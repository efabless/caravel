VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_io_buffer
  CLASS BLOCK ;
  FOREIGN mprj_io_buffer ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 50.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.880 5.200 14.480 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.505 5.200 23.105 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.130 5.200 31.730 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.755 5.200 40.355 43.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.570 5.200 10.170 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.195 5.200 18.795 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.820 5.200 27.420 43.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.445 5.200 36.045 43.760 ;
    END
  END VPWR
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 46.000 39.930 50.000 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 46.000 12.330 50.000 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 46.000 9.570 50.000 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 46.000 6.810 50.000 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 46.000 4.050 50.000 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 46.000 37.170 50.000 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 46.000 34.410 50.000 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 46.000 31.650 50.000 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 46.000 28.890 50.000 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 46.000 26.130 50.000 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 46.000 23.370 50.000 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 46.000 20.610 50.000 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 46.000 17.850 50.000 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 46.000 15.090 50.000 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_in_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 8.880 45.000 9.480 ;
    END
  END mgmt_gpio_in_buf[0]
  PIN mgmt_gpio_in_buf[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 29.280 45.000 29.880 ;
    END
  END mgmt_gpio_in_buf[10]
  PIN mgmt_gpio_in_buf[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 31.320 45.000 31.920 ;
    END
  END mgmt_gpio_in_buf[11]
  PIN mgmt_gpio_in_buf[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 33.360 45.000 33.960 ;
    END
  END mgmt_gpio_in_buf[12]
  PIN mgmt_gpio_in_buf[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 35.400 45.000 36.000 ;
    END
  END mgmt_gpio_in_buf[13]
  PIN mgmt_gpio_in_buf[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 37.440 45.000 38.040 ;
    END
  END mgmt_gpio_in_buf[14]
  PIN mgmt_gpio_in_buf[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 39.480 45.000 40.080 ;
    END
  END mgmt_gpio_in_buf[15]
  PIN mgmt_gpio_in_buf[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 41.520 45.000 42.120 ;
    END
  END mgmt_gpio_in_buf[16]
  PIN mgmt_gpio_in_buf[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 43.560 45.000 44.160 ;
    END
  END mgmt_gpio_in_buf[17]
  PIN mgmt_gpio_in_buf[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 45.600 45.000 46.200 ;
    END
  END mgmt_gpio_in_buf[18]
  PIN mgmt_gpio_in_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 10.920 45.000 11.520 ;
    END
  END mgmt_gpio_in_buf[1]
  PIN mgmt_gpio_in_buf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 12.960 45.000 13.560 ;
    END
  END mgmt_gpio_in_buf[2]
  PIN mgmt_gpio_in_buf[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 15.000 45.000 15.600 ;
    END
  END mgmt_gpio_in_buf[3]
  PIN mgmt_gpio_in_buf[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 17.040 45.000 17.640 ;
    END
  END mgmt_gpio_in_buf[4]
  PIN mgmt_gpio_in_buf[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 19.080 45.000 19.680 ;
    END
  END mgmt_gpio_in_buf[5]
  PIN mgmt_gpio_in_buf[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 21.120 45.000 21.720 ;
    END
  END mgmt_gpio_in_buf[6]
  PIN mgmt_gpio_in_buf[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 23.160 45.000 23.760 ;
    END
  END mgmt_gpio_in_buf[7]
  PIN mgmt_gpio_in_buf[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 25.200 45.000 25.800 ;
    END
  END mgmt_gpio_in_buf[8]
  PIN mgmt_gpio_in_buf[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 27.240 45.000 27.840 ;
    END
  END mgmt_gpio_in_buf[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 2.760 45.000 3.360 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 4.800 45.000 5.400 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 6.840 45.000 7.440 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END mgmt_gpio_oeb_buf[0]
  PIN mgmt_gpio_oeb_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END mgmt_gpio_oeb_buf[1]
  PIN mgmt_gpio_oeb_buf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END mgmt_gpio_oeb_buf[2]
  PIN mgmt_gpio_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END mgmt_gpio_out[9]
  PIN mgmt_gpio_out_buf[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 46.000 41.310 50.000 ;
    END
  END mgmt_gpio_out_buf[0]
  PIN mgmt_gpio_out_buf[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 46.000 13.710 50.000 ;
    END
  END mgmt_gpio_out_buf[10]
  PIN mgmt_gpio_out_buf[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 46.000 10.950 50.000 ;
    END
  END mgmt_gpio_out_buf[11]
  PIN mgmt_gpio_out_buf[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 46.000 8.190 50.000 ;
    END
  END mgmt_gpio_out_buf[12]
  PIN mgmt_gpio_out_buf[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 46.000 5.430 50.000 ;
    END
  END mgmt_gpio_out_buf[13]
  PIN mgmt_gpio_out_buf[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END mgmt_gpio_out_buf[14]
  PIN mgmt_gpio_out_buf[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END mgmt_gpio_out_buf[15]
  PIN mgmt_gpio_out_buf[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END mgmt_gpio_out_buf[16]
  PIN mgmt_gpio_out_buf[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END mgmt_gpio_out_buf[17]
  PIN mgmt_gpio_out_buf[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END mgmt_gpio_out_buf[18]
  PIN mgmt_gpio_out_buf[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 46.000 38.550 50.000 ;
    END
  END mgmt_gpio_out_buf[1]
  PIN mgmt_gpio_out_buf[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 46.000 35.790 50.000 ;
    END
  END mgmt_gpio_out_buf[2]
  PIN mgmt_gpio_out_buf[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 46.000 33.030 50.000 ;
    END
  END mgmt_gpio_out_buf[3]
  PIN mgmt_gpio_out_buf[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 46.000 30.270 50.000 ;
    END
  END mgmt_gpio_out_buf[4]
  PIN mgmt_gpio_out_buf[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 46.000 27.510 50.000 ;
    END
  END mgmt_gpio_out_buf[5]
  PIN mgmt_gpio_out_buf[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 46.000 24.750 50.000 ;
    END
  END mgmt_gpio_out_buf[6]
  PIN mgmt_gpio_out_buf[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 46.000 21.990 50.000 ;
    END
  END mgmt_gpio_out_buf[7]
  PIN mgmt_gpio_out_buf[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 46.000 19.230 50.000 ;
    END
  END mgmt_gpio_out_buf[8]
  PIN mgmt_gpio_out_buf[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 46.000 16.470 50.000 ;
    END
  END mgmt_gpio_out_buf[9]
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 39.560 43.605 ;
      LAYER met1 ;
        RECT 1.450 5.200 43.170 44.500 ;
      LAYER met2 ;
        RECT 1.480 45.720 3.490 46.650 ;
        RECT 4.330 45.720 4.870 46.650 ;
        RECT 5.710 45.720 6.250 46.650 ;
        RECT 7.090 45.720 7.630 46.650 ;
        RECT 8.470 45.720 9.010 46.650 ;
        RECT 9.850 45.720 10.390 46.650 ;
        RECT 11.230 45.720 11.770 46.650 ;
        RECT 12.610 45.720 13.150 46.650 ;
        RECT 13.990 45.720 14.530 46.650 ;
        RECT 15.370 45.720 15.910 46.650 ;
        RECT 16.750 45.720 17.290 46.650 ;
        RECT 18.130 45.720 18.670 46.650 ;
        RECT 19.510 45.720 20.050 46.650 ;
        RECT 20.890 45.720 21.430 46.650 ;
        RECT 22.270 45.720 22.810 46.650 ;
        RECT 23.650 45.720 24.190 46.650 ;
        RECT 25.030 45.720 25.570 46.650 ;
        RECT 26.410 45.720 26.950 46.650 ;
        RECT 27.790 45.720 28.330 46.650 ;
        RECT 29.170 45.720 29.710 46.650 ;
        RECT 30.550 45.720 31.090 46.650 ;
        RECT 31.930 45.720 32.470 46.650 ;
        RECT 33.310 45.720 33.850 46.650 ;
        RECT 34.690 45.720 35.230 46.650 ;
        RECT 36.070 45.720 36.610 46.650 ;
        RECT 37.450 45.720 37.990 46.650 ;
        RECT 38.830 45.720 39.370 46.650 ;
        RECT 40.210 45.720 40.750 46.650 ;
        RECT 41.590 45.720 43.140 46.650 ;
        RECT 1.480 4.280 43.140 45.720 ;
        RECT 2.030 2.875 3.490 4.280 ;
        RECT 4.330 2.875 5.790 4.280 ;
        RECT 6.630 2.875 8.090 4.280 ;
        RECT 8.930 2.875 10.390 4.280 ;
        RECT 11.230 2.875 12.690 4.280 ;
        RECT 13.530 2.875 14.990 4.280 ;
        RECT 15.830 2.875 17.290 4.280 ;
        RECT 18.130 2.875 19.590 4.280 ;
        RECT 20.430 2.875 21.890 4.280 ;
        RECT 22.730 2.875 24.190 4.280 ;
        RECT 25.030 2.875 26.490 4.280 ;
        RECT 27.330 2.875 28.790 4.280 ;
        RECT 29.630 2.875 31.090 4.280 ;
        RECT 31.930 2.875 33.390 4.280 ;
        RECT 34.230 2.875 35.690 4.280 ;
        RECT 36.530 2.875 37.990 4.280 ;
        RECT 38.830 2.875 40.290 4.280 ;
        RECT 41.130 2.875 42.590 4.280 ;
      LAYER met3 ;
        RECT 4.000 45.920 40.600 46.065 ;
        RECT 4.400 45.200 40.600 45.920 ;
        RECT 4.400 44.560 41.090 45.200 ;
        RECT 4.400 44.520 40.600 44.560 ;
        RECT 4.000 43.160 40.600 44.520 ;
        RECT 4.000 42.520 41.090 43.160 ;
        RECT 4.400 41.120 40.600 42.520 ;
        RECT 4.000 40.480 41.090 41.120 ;
        RECT 4.000 39.120 40.600 40.480 ;
        RECT 4.400 39.080 40.600 39.120 ;
        RECT 4.400 38.440 41.090 39.080 ;
        RECT 4.400 37.720 40.600 38.440 ;
        RECT 4.000 37.040 40.600 37.720 ;
        RECT 4.000 36.400 41.090 37.040 ;
        RECT 4.000 35.720 40.600 36.400 ;
        RECT 4.400 35.000 40.600 35.720 ;
        RECT 4.400 34.360 41.090 35.000 ;
        RECT 4.400 34.320 40.600 34.360 ;
        RECT 4.000 32.960 40.600 34.320 ;
        RECT 4.000 32.320 41.090 32.960 ;
        RECT 4.400 30.920 40.600 32.320 ;
        RECT 4.000 30.280 41.090 30.920 ;
        RECT 4.000 28.920 40.600 30.280 ;
        RECT 4.400 28.880 40.600 28.920 ;
        RECT 4.400 28.240 41.090 28.880 ;
        RECT 4.400 27.520 40.600 28.240 ;
        RECT 4.000 26.840 40.600 27.520 ;
        RECT 4.000 26.200 41.090 26.840 ;
        RECT 4.000 25.520 40.600 26.200 ;
        RECT 4.400 24.800 40.600 25.520 ;
        RECT 4.400 24.160 41.090 24.800 ;
        RECT 4.400 24.120 40.600 24.160 ;
        RECT 4.000 22.760 40.600 24.120 ;
        RECT 4.000 22.120 41.090 22.760 ;
        RECT 4.400 20.720 40.600 22.120 ;
        RECT 4.000 20.080 41.090 20.720 ;
        RECT 4.000 18.720 40.600 20.080 ;
        RECT 4.400 18.680 40.600 18.720 ;
        RECT 4.400 18.040 41.090 18.680 ;
        RECT 4.400 17.320 40.600 18.040 ;
        RECT 4.000 16.640 40.600 17.320 ;
        RECT 4.000 16.000 41.090 16.640 ;
        RECT 4.000 15.320 40.600 16.000 ;
        RECT 4.400 14.600 40.600 15.320 ;
        RECT 4.400 13.960 41.090 14.600 ;
        RECT 4.400 13.920 40.600 13.960 ;
        RECT 4.000 12.560 40.600 13.920 ;
        RECT 4.000 11.920 41.090 12.560 ;
        RECT 4.400 10.520 40.600 11.920 ;
        RECT 4.000 9.880 41.090 10.520 ;
        RECT 4.000 8.520 40.600 9.880 ;
        RECT 4.400 8.480 40.600 8.520 ;
        RECT 4.400 7.840 41.090 8.480 ;
        RECT 4.400 7.120 40.600 7.840 ;
        RECT 4.000 6.440 40.600 7.120 ;
        RECT 4.000 5.800 41.090 6.440 ;
        RECT 4.000 5.120 40.600 5.800 ;
        RECT 4.400 4.400 40.600 5.120 ;
        RECT 4.400 3.760 41.090 4.400 ;
        RECT 4.400 3.720 40.600 3.760 ;
        RECT 4.000 2.895 40.600 3.720 ;
  END
END mprj_io_buffer
END LIBRARY

