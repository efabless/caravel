VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_clocking
  CLASS BLOCK ;
  FOREIGN caravel_clocking ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 60.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 1.840 24.060 94.300 25.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.840 40.960 94.300 42.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.110 -0.240 26.710 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.610 -0.240 42.210 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.110 -0.240 57.710 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.610 -0.240 73.210 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.110 -0.240 88.710 54.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 1.840 15.610 94.300 17.210 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.840 32.510 94.300 34.110 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.840 49.410 94.300 51.010 ;
    END
    PORT
      LAYER met4 ;
        RECT 17.360 -0.240 18.960 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.860 -0.240 34.460 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.360 -0.240 49.960 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.860 -0.240 65.460 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.360 -0.240 80.960 54.640 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 56.000 35.790 60.000 ;
    END
  END core_clk
  PIN ext_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 56.000 21.530 60.000 ;
    END
  END ext_clk
  PIN ext_clk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END ext_clk_sel
  PIN ext_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END ext_reset
  PIN pll_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 56.000 78.570 60.000 ;
    END
  END pll_clk
  PIN pll_clk90
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 56.000 92.830 60.000 ;
    END
  END pll_clk90
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 56.000 7.270 60.000 ;
    END
  END resetb
  PIN resetb_sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 56.000 64.310 60.000 ;
    END
  END resetb_sync
  PIN sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 33.360 100.000 33.960 ;
    END
  END sel2[0]
  PIN sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END sel2[1]
  PIN sel2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 48.320 100.000 48.920 ;
    END
  END sel2[2]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 18.400 100.000 19.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.880 100.000 26.480 ;
    END
  END sel[2]
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 56.000 50.050 60.000 ;
    END
  END user_clk
  OBS
      LAYER pwell ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 7.055 -0.050 7.215 0.060 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 20.385 -0.085 20.555 0.085 ;
        RECT 24.060 -0.055 24.180 0.055 ;
        RECT 25.450 -0.085 25.620 0.085 ;
        RECT 26.360 -0.055 26.480 0.055 ;
        RECT 27.285 -0.085 27.455 0.085 ;
        RECT 27.755 -0.050 27.915 0.060 ;
        RECT 30.040 -0.085 30.210 0.085 ;
        RECT 30.505 -0.085 30.675 0.085 ;
        RECT 32.350 -0.085 32.520 0.085 ;
        RECT 34.185 -0.085 34.355 0.085 ;
        RECT 38.335 -0.050 38.495 0.060 ;
        RECT 39.245 -0.085 39.415 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 44.305 -0.085 44.475 0.085 ;
        RECT 47.525 -0.085 47.695 0.085 ;
        RECT 49.360 -0.055 49.480 0.055 ;
        RECT 50.285 -0.085 50.455 0.085 ;
        RECT 56.265 -0.085 56.435 0.085 ;
        RECT 62.245 -0.085 62.415 0.085 ;
        RECT 65.460 -0.055 65.580 0.055 ;
        RECT 66.840 -0.085 67.010 0.085 ;
        RECT 67.300 -0.055 67.420 0.055 ;
        RECT 68.225 -0.085 68.395 0.085 ;
        RECT 74.200 -0.055 74.320 0.055 ;
        RECT 75.125 -0.085 75.295 0.085 ;
        RECT 75.585 -0.085 75.755 0.085 ;
        RECT 79.260 -0.055 79.380 0.055 ;
        RECT 80.185 -0.085 80.355 0.085 ;
        RECT 86.165 -0.085 86.335 0.085 ;
        RECT 89.395 -0.050 89.555 0.060 ;
        RECT 91.225 -0.085 91.395 0.085 ;
        RECT 92.145 -0.085 92.315 0.085 ;
        RECT 93.985 -0.085 94.155 0.085 ;
      LAYER li1 ;
        RECT 1.065 0.085 94.300 54.485 ;
        RECT 1.065 0.000 1.840 0.085 ;
      LAYER li1 ;
        RECT 1.840 -0.085 94.300 0.085 ;
      LAYER met1 ;
        RECT 1.005 0.000 94.300 54.640 ;
        RECT 1.840 -0.240 94.300 0.000 ;
      LAYER met2 ;
        RECT 3.320 55.720 6.710 56.285 ;
        RECT 7.550 55.720 20.970 56.285 ;
        RECT 21.810 55.720 35.230 56.285 ;
        RECT 36.070 55.720 49.490 56.285 ;
        RECT 50.330 55.720 63.750 56.285 ;
        RECT 64.590 55.720 78.010 56.285 ;
        RECT 78.850 55.720 92.270 56.285 ;
        RECT 93.110 55.720 94.210 56.285 ;
        RECT 3.320 0.000 94.210 55.720 ;
        RECT 25.140 -0.240 26.680 0.000 ;
        RECT 40.640 -0.240 42.180 0.000 ;
        RECT 56.140 -0.240 57.680 0.000 ;
        RECT 71.640 -0.240 73.180 0.000 ;
        RECT 87.140 -0.240 88.680 0.000 ;
      LAYER met3 ;
        RECT 12.485 55.400 95.600 56.265 ;
        RECT 12.485 49.320 96.000 55.400 ;
        RECT 12.485 47.920 95.600 49.320 ;
        RECT 12.485 41.840 96.000 47.920 ;
        RECT 12.485 40.440 95.600 41.840 ;
        RECT 12.485 34.360 96.000 40.440 ;
        RECT 12.485 32.960 95.600 34.360 ;
        RECT 12.485 26.880 96.000 32.960 ;
        RECT 12.485 25.480 95.600 26.880 ;
        RECT 12.485 19.400 96.000 25.480 ;
        RECT 12.485 18.000 95.600 19.400 ;
        RECT 12.485 11.920 96.000 18.000 ;
        RECT 12.485 10.520 95.600 11.920 ;
        RECT 12.485 4.440 96.000 10.520 ;
        RECT 12.485 3.040 95.600 4.440 ;
        RECT 12.485 0.000 96.000 3.040 ;
        RECT 25.110 -0.165 26.710 0.000 ;
        RECT 40.610 -0.165 42.210 0.000 ;
        RECT 56.110 -0.165 57.710 0.000 ;
        RECT 71.610 -0.165 73.210 0.000 ;
        RECT 87.110 -0.165 88.710 0.000 ;
  END
END caravel_clocking
END LIBRARY

