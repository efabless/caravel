VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128
  CLASS BLOCK ;
  FOREIGN RAM128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 406.180 BY 437.920 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 51.720 406.180 52.320 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 85.040 406.180 85.640 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 118.360 406.180 118.960 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 151.680 406.180 152.280 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 185.000 406.180 185.600 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 218.320 406.180 218.920 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 251.640 406.180 252.240 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 284.960 406.180 285.560 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 435.920 10.490 437.920 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 435.920 134.690 437.920 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 435.920 147.110 437.920 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 435.920 159.530 437.920 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 435.920 171.950 437.920 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 435.920 184.370 437.920 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 435.920 196.790 437.920 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 435.920 209.210 437.920 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 435.920 221.630 437.920 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 435.920 234.050 437.920 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 435.920 246.470 437.920 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 435.920 22.910 437.920 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 435.920 258.890 437.920 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 435.920 271.310 437.920 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 435.920 283.730 437.920 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 435.920 296.150 437.920 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 435.920 308.570 437.920 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 435.920 320.990 437.920 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 435.920 333.410 437.920 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 435.920 345.830 437.920 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 435.920 358.250 437.920 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 435.920 370.670 437.920 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 435.920 35.330 437.920 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 435.920 383.090 437.920 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 435.920 395.510 437.920 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 435.920 47.750 437.920 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 435.920 60.170 437.920 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 435.920 72.590 437.920 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 435.920 85.010 437.920 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 435.920 97.430 437.920 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 435.920 109.850 437.920 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 435.920 122.270 437.920 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 18.400 406.180 19.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 435.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 435.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 435.440 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 318.280 406.180 318.880 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 351.600 406.180 352.200 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 384.920 406.180 385.520 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 404.180 418.240 406.180 418.840 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 403.420 435.285 ;
      LAYER met1 ;
        RECT 2.460 0.040 406.110 437.880 ;
      LAYER met2 ;
        RECT 2.860 435.640 9.930 437.910 ;
        RECT 10.770 435.640 22.350 437.910 ;
        RECT 23.190 435.640 34.770 437.910 ;
        RECT 35.610 435.640 47.190 437.910 ;
        RECT 48.030 435.640 59.610 437.910 ;
        RECT 60.450 435.640 72.030 437.910 ;
        RECT 72.870 435.640 84.450 437.910 ;
        RECT 85.290 435.640 96.870 437.910 ;
        RECT 97.710 435.640 109.290 437.910 ;
        RECT 110.130 435.640 121.710 437.910 ;
        RECT 122.550 435.640 134.130 437.910 ;
        RECT 134.970 435.640 146.550 437.910 ;
        RECT 147.390 435.640 158.970 437.910 ;
        RECT 159.810 435.640 171.390 437.910 ;
        RECT 172.230 435.640 183.810 437.910 ;
        RECT 184.650 435.640 196.230 437.910 ;
        RECT 197.070 435.640 208.650 437.910 ;
        RECT 209.490 435.640 221.070 437.910 ;
        RECT 221.910 435.640 233.490 437.910 ;
        RECT 234.330 435.640 245.910 437.910 ;
        RECT 246.750 435.640 258.330 437.910 ;
        RECT 259.170 435.640 270.750 437.910 ;
        RECT 271.590 435.640 283.170 437.910 ;
        RECT 284.010 435.640 295.590 437.910 ;
        RECT 296.430 435.640 308.010 437.910 ;
        RECT 308.850 435.640 320.430 437.910 ;
        RECT 321.270 435.640 332.850 437.910 ;
        RECT 333.690 435.640 345.270 437.910 ;
        RECT 346.110 435.640 357.690 437.910 ;
        RECT 358.530 435.640 370.110 437.910 ;
        RECT 370.950 435.640 382.530 437.910 ;
        RECT 383.370 435.640 394.950 437.910 ;
        RECT 395.790 435.640 406.080 437.910 ;
        RECT 2.860 2.280 406.080 435.640 ;
        RECT 2.860 0.010 9.930 2.280 ;
        RECT 10.770 0.010 22.350 2.280 ;
        RECT 23.190 0.010 34.770 2.280 ;
        RECT 35.610 0.010 47.190 2.280 ;
        RECT 48.030 0.010 59.610 2.280 ;
        RECT 60.450 0.010 72.030 2.280 ;
        RECT 72.870 0.010 84.450 2.280 ;
        RECT 85.290 0.010 96.870 2.280 ;
        RECT 97.710 0.010 109.290 2.280 ;
        RECT 110.130 0.010 121.710 2.280 ;
        RECT 122.550 0.010 134.130 2.280 ;
        RECT 134.970 0.010 146.550 2.280 ;
        RECT 147.390 0.010 158.970 2.280 ;
        RECT 159.810 0.010 171.390 2.280 ;
        RECT 172.230 0.010 183.810 2.280 ;
        RECT 184.650 0.010 196.230 2.280 ;
        RECT 197.070 0.010 208.650 2.280 ;
        RECT 209.490 0.010 221.070 2.280 ;
        RECT 221.910 0.010 233.490 2.280 ;
        RECT 234.330 0.010 245.910 2.280 ;
        RECT 246.750 0.010 258.330 2.280 ;
        RECT 259.170 0.010 270.750 2.280 ;
        RECT 271.590 0.010 283.170 2.280 ;
        RECT 284.010 0.010 295.590 2.280 ;
        RECT 296.430 0.010 308.010 2.280 ;
        RECT 308.850 0.010 320.430 2.280 ;
        RECT 321.270 0.010 332.850 2.280 ;
        RECT 333.690 0.010 345.270 2.280 ;
        RECT 346.110 0.010 357.690 2.280 ;
        RECT 358.530 0.010 370.110 2.280 ;
        RECT 370.950 0.010 382.530 2.280 ;
        RECT 383.370 0.010 394.950 2.280 ;
        RECT 395.790 0.010 406.080 2.280 ;
      LAYER met3 ;
        RECT 3.285 419.240 404.490 437.745 ;
        RECT 3.285 417.840 403.780 419.240 ;
        RECT 3.285 385.920 404.490 417.840 ;
        RECT 3.285 384.520 403.780 385.920 ;
        RECT 3.285 352.600 404.490 384.520 ;
        RECT 3.285 351.200 403.780 352.600 ;
        RECT 3.285 319.280 404.490 351.200 ;
        RECT 3.285 317.880 403.780 319.280 ;
        RECT 3.285 285.960 404.490 317.880 ;
        RECT 3.285 284.560 403.780 285.960 ;
        RECT 3.285 252.640 404.490 284.560 ;
        RECT 3.285 251.240 403.780 252.640 ;
        RECT 3.285 219.320 404.490 251.240 ;
        RECT 3.285 217.920 403.780 219.320 ;
        RECT 3.285 186.000 404.490 217.920 ;
        RECT 3.285 184.600 403.780 186.000 ;
        RECT 3.285 152.680 404.490 184.600 ;
        RECT 3.285 151.280 403.780 152.680 ;
        RECT 3.285 119.360 404.490 151.280 ;
        RECT 3.285 117.960 403.780 119.360 ;
        RECT 3.285 86.040 404.490 117.960 ;
        RECT 3.285 84.640 403.780 86.040 ;
        RECT 3.285 52.720 404.490 84.640 ;
        RECT 3.285 51.320 403.780 52.720 ;
        RECT 3.285 19.400 404.490 51.320 ;
        RECT 3.285 18.000 403.780 19.400 ;
        RECT 3.285 0.175 404.490 18.000 ;
      LAYER met4 ;
        RECT 97.815 435.840 384.265 437.065 ;
        RECT 97.815 6.975 171.480 435.840 ;
        RECT 173.880 6.975 248.280 435.840 ;
        RECT 250.680 6.975 325.080 435.840 ;
        RECT 327.480 6.975 384.265 435.840 ;
  END
END RAM128
END LIBRARY

