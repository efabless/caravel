module housekeeping (debug_in,
    debug_mode,
    debug_oeb,
    debug_out,
    pad_flash_clk,
    pad_flash_clk_oeb,
    pad_flash_csb,
    pad_flash_csb_oeb,
    pad_flash_io0_di,
    pad_flash_io0_do,
    pad_flash_io0_ieb,
    pad_flash_io0_oeb,
    pad_flash_io1_di,
    pad_flash_io1_do,
    pad_flash_io1_ieb,
    pad_flash_io1_oeb,
    pll_bypass,
    pll_dco_ena,
    pll_ena,
    porb,
    qspi_enabled,
    reset,
    ser_rx,
    ser_tx,
    serial_clock,
    serial_data_1,
    serial_data_2,
    serial_load,
    serial_resetn,
    spi_csb,
    spi_enabled,
    spi_sck,
    spi_sdi,
    spi_sdo,
    spi_sdoenb,
    spimemio_flash_clk,
    spimemio_flash_csb,
    spimemio_flash_io0_di,
    spimemio_flash_io0_do,
    spimemio_flash_io0_oeb,
    spimemio_flash_io1_di,
    spimemio_flash_io1_do,
    spimemio_flash_io1_oeb,
    spimemio_flash_io2_di,
    spimemio_flash_io2_do,
    spimemio_flash_io2_oeb,
    spimemio_flash_io3_di,
    spimemio_flash_io3_do,
    spimemio_flash_io3_oeb,
    trap,
    uart_enabled,
    user_clock,
    usr1_vcc_pwrgood,
    usr1_vdd_pwrgood,
    usr2_vcc_pwrgood,
    usr2_vdd_pwrgood,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rstn_i,
    wb_stb_i,
    wb_we_i,
    irq,
    mask_rev_in,
    mgmt_gpio_in,
    mgmt_gpio_oeb,
    mgmt_gpio_out,
    pll90_sel,
    pll_div,
    pll_sel,
    pll_trim,
    pwr_ctrl_out,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output debug_in;
 input debug_mode;
 input debug_oeb;
 input debug_out;
 output pad_flash_clk;
 output pad_flash_clk_oeb;
 output pad_flash_csb;
 output pad_flash_csb_oeb;
 input pad_flash_io0_di;
 output pad_flash_io0_do;
 output pad_flash_io0_ieb;
 output pad_flash_io0_oeb;
 input pad_flash_io1_di;
 output pad_flash_io1_do;
 output pad_flash_io1_ieb;
 output pad_flash_io1_oeb;
 output pll_bypass;
 output pll_dco_ena;
 output pll_ena;
 input porb;
 input qspi_enabled;
 output reset;
 output ser_rx;
 input ser_tx;
 output serial_clock;
 output serial_data_1;
 output serial_data_2;
 output serial_load;
 output serial_resetn;
 input spi_csb;
 input spi_enabled;
 input spi_sck;
 output spi_sdi;
 input spi_sdo;
 input spi_sdoenb;
 input spimemio_flash_clk;
 input spimemio_flash_csb;
 output spimemio_flash_io0_di;
 input spimemio_flash_io0_do;
 input spimemio_flash_io0_oeb;
 output spimemio_flash_io1_di;
 input spimemio_flash_io1_do;
 input spimemio_flash_io1_oeb;
 output spimemio_flash_io2_di;
 input spimemio_flash_io2_do;
 input spimemio_flash_io2_oeb;
 output spimemio_flash_io3_di;
 input spimemio_flash_io3_do;
 input spimemio_flash_io3_oeb;
 input trap;
 input uart_enabled;
 input user_clock;
 input usr1_vcc_pwrgood;
 input usr1_vdd_pwrgood;
 input usr2_vcc_pwrgood;
 input usr2_vdd_pwrgood;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rstn_i;
 input wb_stb_i;
 input wb_we_i;
 output [2:0] irq;
 input [31:0] mask_rev_in;
 input [37:0] mgmt_gpio_in;
 output [37:0] mgmt_gpio_oeb;
 output [37:0] mgmt_gpio_out;
 output [2:0] pll90_sel;
 output [4:0] pll_div;
 output [2:0] pll_sel;
 output [25:0] pll_trim;
 output [3:0] pwr_ctrl_out;
 input [31:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire clknet_0_wb_clk_i;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire net461;
 wire clk1_output_dest;
 wire clk2_output_dest;
 wire csclk;
 wire \gpio_configure[0][0] ;
 wire \gpio_configure[0][10] ;
 wire \gpio_configure[0][11] ;
 wire \gpio_configure[0][12] ;
 wire \gpio_configure[0][1] ;
 wire \gpio_configure[0][2] ;
 wire \gpio_configure[0][3] ;
 wire \gpio_configure[0][4] ;
 wire \gpio_configure[0][5] ;
 wire \gpio_configure[0][6] ;
 wire \gpio_configure[0][7] ;
 wire \gpio_configure[0][8] ;
 wire \gpio_configure[0][9] ;
 wire \gpio_configure[10][0] ;
 wire \gpio_configure[10][10] ;
 wire \gpio_configure[10][11] ;
 wire \gpio_configure[10][12] ;
 wire \gpio_configure[10][1] ;
 wire \gpio_configure[10][2] ;
 wire \gpio_configure[10][3] ;
 wire \gpio_configure[10][4] ;
 wire \gpio_configure[10][5] ;
 wire \gpio_configure[10][6] ;
 wire \gpio_configure[10][7] ;
 wire \gpio_configure[10][8] ;
 wire \gpio_configure[10][9] ;
 wire \gpio_configure[11][0] ;
 wire \gpio_configure[11][10] ;
 wire \gpio_configure[11][11] ;
 wire \gpio_configure[11][12] ;
 wire \gpio_configure[11][1] ;
 wire \gpio_configure[11][2] ;
 wire \gpio_configure[11][3] ;
 wire \gpio_configure[11][4] ;
 wire \gpio_configure[11][5] ;
 wire \gpio_configure[11][6] ;
 wire \gpio_configure[11][7] ;
 wire \gpio_configure[11][8] ;
 wire \gpio_configure[11][9] ;
 wire \gpio_configure[12][0] ;
 wire \gpio_configure[12][10] ;
 wire \gpio_configure[12][11] ;
 wire \gpio_configure[12][12] ;
 wire \gpio_configure[12][1] ;
 wire \gpio_configure[12][2] ;
 wire \gpio_configure[12][3] ;
 wire \gpio_configure[12][4] ;
 wire \gpio_configure[12][5] ;
 wire \gpio_configure[12][6] ;
 wire \gpio_configure[12][7] ;
 wire \gpio_configure[12][8] ;
 wire \gpio_configure[12][9] ;
 wire \gpio_configure[13][0] ;
 wire \gpio_configure[13][10] ;
 wire \gpio_configure[13][11] ;
 wire \gpio_configure[13][12] ;
 wire \gpio_configure[13][1] ;
 wire \gpio_configure[13][2] ;
 wire \gpio_configure[13][3] ;
 wire \gpio_configure[13][4] ;
 wire \gpio_configure[13][5] ;
 wire \gpio_configure[13][6] ;
 wire \gpio_configure[13][7] ;
 wire \gpio_configure[13][8] ;
 wire \gpio_configure[13][9] ;
 wire \gpio_configure[14][0] ;
 wire \gpio_configure[14][10] ;
 wire \gpio_configure[14][11] ;
 wire \gpio_configure[14][12] ;
 wire \gpio_configure[14][1] ;
 wire \gpio_configure[14][2] ;
 wire \gpio_configure[14][3] ;
 wire \gpio_configure[14][4] ;
 wire \gpio_configure[14][5] ;
 wire \gpio_configure[14][6] ;
 wire \gpio_configure[14][7] ;
 wire \gpio_configure[14][8] ;
 wire \gpio_configure[14][9] ;
 wire \gpio_configure[15][0] ;
 wire \gpio_configure[15][10] ;
 wire \gpio_configure[15][11] ;
 wire \gpio_configure[15][12] ;
 wire \gpio_configure[15][1] ;
 wire \gpio_configure[15][2] ;
 wire \gpio_configure[15][3] ;
 wire \gpio_configure[15][4] ;
 wire \gpio_configure[15][5] ;
 wire \gpio_configure[15][6] ;
 wire \gpio_configure[15][7] ;
 wire \gpio_configure[15][8] ;
 wire \gpio_configure[15][9] ;
 wire \gpio_configure[16][0] ;
 wire \gpio_configure[16][10] ;
 wire \gpio_configure[16][11] ;
 wire \gpio_configure[16][12] ;
 wire \gpio_configure[16][1] ;
 wire \gpio_configure[16][2] ;
 wire \gpio_configure[16][3] ;
 wire \gpio_configure[16][4] ;
 wire \gpio_configure[16][5] ;
 wire \gpio_configure[16][6] ;
 wire \gpio_configure[16][7] ;
 wire \gpio_configure[16][8] ;
 wire \gpio_configure[16][9] ;
 wire \gpio_configure[17][0] ;
 wire \gpio_configure[17][10] ;
 wire \gpio_configure[17][11] ;
 wire \gpio_configure[17][12] ;
 wire \gpio_configure[17][1] ;
 wire \gpio_configure[17][2] ;
 wire \gpio_configure[17][3] ;
 wire \gpio_configure[17][4] ;
 wire \gpio_configure[17][5] ;
 wire \gpio_configure[17][6] ;
 wire \gpio_configure[17][7] ;
 wire \gpio_configure[17][8] ;
 wire \gpio_configure[17][9] ;
 wire \gpio_configure[18][0] ;
 wire \gpio_configure[18][10] ;
 wire \gpio_configure[18][11] ;
 wire \gpio_configure[18][12] ;
 wire \gpio_configure[18][1] ;
 wire \gpio_configure[18][2] ;
 wire \gpio_configure[18][3] ;
 wire \gpio_configure[18][4] ;
 wire \gpio_configure[18][5] ;
 wire \gpio_configure[18][6] ;
 wire \gpio_configure[18][7] ;
 wire \gpio_configure[18][8] ;
 wire \gpio_configure[18][9] ;
 wire \gpio_configure[19][0] ;
 wire \gpio_configure[19][10] ;
 wire \gpio_configure[19][11] ;
 wire \gpio_configure[19][12] ;
 wire \gpio_configure[19][1] ;
 wire \gpio_configure[19][2] ;
 wire \gpio_configure[19][3] ;
 wire \gpio_configure[19][4] ;
 wire \gpio_configure[19][5] ;
 wire \gpio_configure[19][6] ;
 wire \gpio_configure[19][7] ;
 wire \gpio_configure[19][8] ;
 wire \gpio_configure[19][9] ;
 wire \gpio_configure[1][0] ;
 wire \gpio_configure[1][10] ;
 wire \gpio_configure[1][11] ;
 wire \gpio_configure[1][12] ;
 wire \gpio_configure[1][1] ;
 wire \gpio_configure[1][2] ;
 wire \gpio_configure[1][3] ;
 wire \gpio_configure[1][4] ;
 wire \gpio_configure[1][5] ;
 wire \gpio_configure[1][6] ;
 wire \gpio_configure[1][7] ;
 wire \gpio_configure[1][8] ;
 wire \gpio_configure[1][9] ;
 wire \gpio_configure[20][0] ;
 wire \gpio_configure[20][10] ;
 wire \gpio_configure[20][11] ;
 wire \gpio_configure[20][12] ;
 wire \gpio_configure[20][1] ;
 wire \gpio_configure[20][2] ;
 wire \gpio_configure[20][3] ;
 wire \gpio_configure[20][4] ;
 wire \gpio_configure[20][5] ;
 wire \gpio_configure[20][6] ;
 wire \gpio_configure[20][7] ;
 wire \gpio_configure[20][8] ;
 wire \gpio_configure[20][9] ;
 wire \gpio_configure[21][0] ;
 wire \gpio_configure[21][10] ;
 wire \gpio_configure[21][11] ;
 wire \gpio_configure[21][12] ;
 wire \gpio_configure[21][1] ;
 wire \gpio_configure[21][2] ;
 wire \gpio_configure[21][3] ;
 wire \gpio_configure[21][4] ;
 wire \gpio_configure[21][5] ;
 wire \gpio_configure[21][6] ;
 wire \gpio_configure[21][7] ;
 wire \gpio_configure[21][8] ;
 wire \gpio_configure[21][9] ;
 wire \gpio_configure[22][0] ;
 wire \gpio_configure[22][10] ;
 wire \gpio_configure[22][11] ;
 wire \gpio_configure[22][12] ;
 wire \gpio_configure[22][1] ;
 wire \gpio_configure[22][2] ;
 wire \gpio_configure[22][3] ;
 wire \gpio_configure[22][4] ;
 wire \gpio_configure[22][5] ;
 wire \gpio_configure[22][6] ;
 wire \gpio_configure[22][7] ;
 wire \gpio_configure[22][8] ;
 wire \gpio_configure[22][9] ;
 wire \gpio_configure[23][0] ;
 wire \gpio_configure[23][10] ;
 wire \gpio_configure[23][11] ;
 wire \gpio_configure[23][12] ;
 wire \gpio_configure[23][1] ;
 wire \gpio_configure[23][2] ;
 wire \gpio_configure[23][3] ;
 wire \gpio_configure[23][4] ;
 wire \gpio_configure[23][5] ;
 wire \gpio_configure[23][6] ;
 wire \gpio_configure[23][7] ;
 wire \gpio_configure[23][8] ;
 wire \gpio_configure[23][9] ;
 wire \gpio_configure[24][0] ;
 wire \gpio_configure[24][10] ;
 wire \gpio_configure[24][11] ;
 wire \gpio_configure[24][12] ;
 wire \gpio_configure[24][1] ;
 wire \gpio_configure[24][2] ;
 wire \gpio_configure[24][3] ;
 wire \gpio_configure[24][4] ;
 wire \gpio_configure[24][5] ;
 wire \gpio_configure[24][6] ;
 wire \gpio_configure[24][7] ;
 wire \gpio_configure[24][8] ;
 wire \gpio_configure[24][9] ;
 wire \gpio_configure[25][0] ;
 wire \gpio_configure[25][10] ;
 wire \gpio_configure[25][11] ;
 wire \gpio_configure[25][12] ;
 wire \gpio_configure[25][1] ;
 wire \gpio_configure[25][2] ;
 wire \gpio_configure[25][3] ;
 wire \gpio_configure[25][4] ;
 wire \gpio_configure[25][5] ;
 wire \gpio_configure[25][6] ;
 wire \gpio_configure[25][7] ;
 wire \gpio_configure[25][8] ;
 wire \gpio_configure[25][9] ;
 wire \gpio_configure[26][0] ;
 wire \gpio_configure[26][10] ;
 wire \gpio_configure[26][11] ;
 wire \gpio_configure[26][12] ;
 wire \gpio_configure[26][1] ;
 wire \gpio_configure[26][2] ;
 wire \gpio_configure[26][3] ;
 wire \gpio_configure[26][4] ;
 wire \gpio_configure[26][5] ;
 wire \gpio_configure[26][6] ;
 wire \gpio_configure[26][7] ;
 wire \gpio_configure[26][8] ;
 wire \gpio_configure[26][9] ;
 wire \gpio_configure[27][0] ;
 wire \gpio_configure[27][10] ;
 wire \gpio_configure[27][11] ;
 wire \gpio_configure[27][12] ;
 wire \gpio_configure[27][1] ;
 wire \gpio_configure[27][2] ;
 wire \gpio_configure[27][3] ;
 wire \gpio_configure[27][4] ;
 wire \gpio_configure[27][5] ;
 wire \gpio_configure[27][6] ;
 wire \gpio_configure[27][7] ;
 wire \gpio_configure[27][8] ;
 wire \gpio_configure[27][9] ;
 wire \gpio_configure[28][0] ;
 wire \gpio_configure[28][10] ;
 wire \gpio_configure[28][11] ;
 wire \gpio_configure[28][12] ;
 wire \gpio_configure[28][1] ;
 wire \gpio_configure[28][2] ;
 wire \gpio_configure[28][3] ;
 wire \gpio_configure[28][4] ;
 wire \gpio_configure[28][5] ;
 wire \gpio_configure[28][6] ;
 wire \gpio_configure[28][7] ;
 wire \gpio_configure[28][8] ;
 wire \gpio_configure[28][9] ;
 wire \gpio_configure[29][0] ;
 wire \gpio_configure[29][10] ;
 wire \gpio_configure[29][11] ;
 wire \gpio_configure[29][12] ;
 wire \gpio_configure[29][1] ;
 wire \gpio_configure[29][2] ;
 wire \gpio_configure[29][3] ;
 wire \gpio_configure[29][4] ;
 wire \gpio_configure[29][5] ;
 wire \gpio_configure[29][6] ;
 wire \gpio_configure[29][7] ;
 wire \gpio_configure[29][8] ;
 wire \gpio_configure[29][9] ;
 wire \gpio_configure[2][0] ;
 wire \gpio_configure[2][10] ;
 wire \gpio_configure[2][11] ;
 wire \gpio_configure[2][12] ;
 wire \gpio_configure[2][1] ;
 wire \gpio_configure[2][2] ;
 wire \gpio_configure[2][3] ;
 wire \gpio_configure[2][4] ;
 wire \gpio_configure[2][5] ;
 wire \gpio_configure[2][6] ;
 wire \gpio_configure[2][7] ;
 wire \gpio_configure[2][8] ;
 wire \gpio_configure[2][9] ;
 wire \gpio_configure[30][0] ;
 wire \gpio_configure[30][10] ;
 wire \gpio_configure[30][11] ;
 wire \gpio_configure[30][12] ;
 wire \gpio_configure[30][1] ;
 wire \gpio_configure[30][2] ;
 wire \gpio_configure[30][3] ;
 wire \gpio_configure[30][4] ;
 wire \gpio_configure[30][5] ;
 wire \gpio_configure[30][6] ;
 wire \gpio_configure[30][7] ;
 wire \gpio_configure[30][8] ;
 wire \gpio_configure[30][9] ;
 wire \gpio_configure[31][0] ;
 wire \gpio_configure[31][10] ;
 wire \gpio_configure[31][11] ;
 wire \gpio_configure[31][12] ;
 wire \gpio_configure[31][1] ;
 wire \gpio_configure[31][2] ;
 wire \gpio_configure[31][3] ;
 wire \gpio_configure[31][4] ;
 wire \gpio_configure[31][5] ;
 wire \gpio_configure[31][6] ;
 wire \gpio_configure[31][7] ;
 wire \gpio_configure[31][8] ;
 wire \gpio_configure[31][9] ;
 wire \gpio_configure[32][0] ;
 wire \gpio_configure[32][10] ;
 wire \gpio_configure[32][11] ;
 wire \gpio_configure[32][12] ;
 wire \gpio_configure[32][1] ;
 wire \gpio_configure[32][2] ;
 wire \gpio_configure[32][3] ;
 wire \gpio_configure[32][4] ;
 wire \gpio_configure[32][5] ;
 wire \gpio_configure[32][6] ;
 wire \gpio_configure[32][7] ;
 wire \gpio_configure[32][8] ;
 wire \gpio_configure[32][9] ;
 wire \gpio_configure[33][0] ;
 wire \gpio_configure[33][10] ;
 wire \gpio_configure[33][11] ;
 wire \gpio_configure[33][12] ;
 wire \gpio_configure[33][1] ;
 wire \gpio_configure[33][2] ;
 wire \gpio_configure[33][3] ;
 wire \gpio_configure[33][4] ;
 wire \gpio_configure[33][5] ;
 wire \gpio_configure[33][6] ;
 wire \gpio_configure[33][7] ;
 wire \gpio_configure[33][8] ;
 wire \gpio_configure[33][9] ;
 wire \gpio_configure[34][0] ;
 wire \gpio_configure[34][10] ;
 wire \gpio_configure[34][11] ;
 wire \gpio_configure[34][12] ;
 wire \gpio_configure[34][1] ;
 wire \gpio_configure[34][2] ;
 wire \gpio_configure[34][3] ;
 wire \gpio_configure[34][4] ;
 wire \gpio_configure[34][5] ;
 wire \gpio_configure[34][6] ;
 wire \gpio_configure[34][7] ;
 wire \gpio_configure[34][8] ;
 wire \gpio_configure[34][9] ;
 wire \gpio_configure[35][0] ;
 wire \gpio_configure[35][10] ;
 wire \gpio_configure[35][11] ;
 wire \gpio_configure[35][12] ;
 wire \gpio_configure[35][1] ;
 wire \gpio_configure[35][2] ;
 wire \gpio_configure[35][3] ;
 wire \gpio_configure[35][4] ;
 wire \gpio_configure[35][5] ;
 wire \gpio_configure[35][6] ;
 wire \gpio_configure[35][7] ;
 wire \gpio_configure[35][8] ;
 wire \gpio_configure[35][9] ;
 wire \gpio_configure[36][0] ;
 wire \gpio_configure[36][10] ;
 wire \gpio_configure[36][11] ;
 wire \gpio_configure[36][12] ;
 wire \gpio_configure[36][1] ;
 wire \gpio_configure[36][2] ;
 wire \gpio_configure[36][3] ;
 wire \gpio_configure[36][4] ;
 wire \gpio_configure[36][5] ;
 wire \gpio_configure[36][6] ;
 wire \gpio_configure[36][7] ;
 wire \gpio_configure[36][8] ;
 wire \gpio_configure[36][9] ;
 wire \gpio_configure[37][0] ;
 wire \gpio_configure[37][10] ;
 wire \gpio_configure[37][11] ;
 wire \gpio_configure[37][12] ;
 wire \gpio_configure[37][1] ;
 wire \gpio_configure[37][2] ;
 wire \gpio_configure[37][3] ;
 wire \gpio_configure[37][4] ;
 wire \gpio_configure[37][5] ;
 wire \gpio_configure[37][6] ;
 wire \gpio_configure[37][7] ;
 wire \gpio_configure[37][8] ;
 wire \gpio_configure[37][9] ;
 wire \gpio_configure[3][0] ;
 wire \gpio_configure[3][10] ;
 wire \gpio_configure[3][11] ;
 wire \gpio_configure[3][12] ;
 wire \gpio_configure[3][1] ;
 wire \gpio_configure[3][2] ;
 wire \gpio_configure[3][3] ;
 wire \gpio_configure[3][4] ;
 wire \gpio_configure[3][5] ;
 wire \gpio_configure[3][6] ;
 wire \gpio_configure[3][7] ;
 wire \gpio_configure[3][8] ;
 wire \gpio_configure[3][9] ;
 wire \gpio_configure[4][0] ;
 wire \gpio_configure[4][10] ;
 wire \gpio_configure[4][11] ;
 wire \gpio_configure[4][12] ;
 wire \gpio_configure[4][1] ;
 wire \gpio_configure[4][2] ;
 wire \gpio_configure[4][3] ;
 wire \gpio_configure[4][4] ;
 wire \gpio_configure[4][5] ;
 wire \gpio_configure[4][6] ;
 wire \gpio_configure[4][7] ;
 wire \gpio_configure[4][8] ;
 wire \gpio_configure[4][9] ;
 wire \gpio_configure[5][0] ;
 wire \gpio_configure[5][10] ;
 wire \gpio_configure[5][11] ;
 wire \gpio_configure[5][12] ;
 wire \gpio_configure[5][1] ;
 wire \gpio_configure[5][2] ;
 wire \gpio_configure[5][3] ;
 wire \gpio_configure[5][4] ;
 wire \gpio_configure[5][5] ;
 wire \gpio_configure[5][6] ;
 wire \gpio_configure[5][7] ;
 wire \gpio_configure[5][8] ;
 wire \gpio_configure[5][9] ;
 wire \gpio_configure[6][0] ;
 wire \gpio_configure[6][10] ;
 wire \gpio_configure[6][11] ;
 wire \gpio_configure[6][12] ;
 wire \gpio_configure[6][1] ;
 wire \gpio_configure[6][2] ;
 wire \gpio_configure[6][3] ;
 wire \gpio_configure[6][4] ;
 wire \gpio_configure[6][5] ;
 wire \gpio_configure[6][6] ;
 wire \gpio_configure[6][7] ;
 wire \gpio_configure[6][8] ;
 wire \gpio_configure[6][9] ;
 wire \gpio_configure[7][0] ;
 wire \gpio_configure[7][10] ;
 wire \gpio_configure[7][11] ;
 wire \gpio_configure[7][12] ;
 wire \gpio_configure[7][1] ;
 wire \gpio_configure[7][2] ;
 wire \gpio_configure[7][3] ;
 wire \gpio_configure[7][4] ;
 wire \gpio_configure[7][5] ;
 wire \gpio_configure[7][6] ;
 wire \gpio_configure[7][7] ;
 wire \gpio_configure[7][8] ;
 wire \gpio_configure[7][9] ;
 wire \gpio_configure[8][0] ;
 wire \gpio_configure[8][10] ;
 wire \gpio_configure[8][11] ;
 wire \gpio_configure[8][12] ;
 wire \gpio_configure[8][1] ;
 wire \gpio_configure[8][2] ;
 wire \gpio_configure[8][3] ;
 wire \gpio_configure[8][4] ;
 wire \gpio_configure[8][5] ;
 wire \gpio_configure[8][6] ;
 wire \gpio_configure[8][7] ;
 wire \gpio_configure[8][8] ;
 wire \gpio_configure[8][9] ;
 wire \gpio_configure[9][0] ;
 wire \gpio_configure[9][10] ;
 wire \gpio_configure[9][11] ;
 wire \gpio_configure[9][12] ;
 wire \gpio_configure[9][1] ;
 wire \gpio_configure[9][2] ;
 wire \gpio_configure[9][3] ;
 wire \gpio_configure[9][4] ;
 wire \gpio_configure[9][5] ;
 wire \gpio_configure[9][6] ;
 wire \gpio_configure[9][7] ;
 wire \gpio_configure[9][8] ;
 wire \gpio_configure[9][9] ;
 wire \hkspi.SDO ;
 wire \hkspi.addr[0] ;
 wire \hkspi.addr[1] ;
 wire \hkspi.addr[2] ;
 wire \hkspi.addr[3] ;
 wire \hkspi.addr[4] ;
 wire \hkspi.addr[5] ;
 wire \hkspi.addr[6] ;
 wire \hkspi.addr[7] ;
 wire \hkspi.count[0] ;
 wire \hkspi.count[1] ;
 wire \hkspi.count[2] ;
 wire \hkspi.fixed[0] ;
 wire \hkspi.fixed[1] ;
 wire \hkspi.fixed[2] ;
 wire \hkspi.ldata[0] ;
 wire \hkspi.ldata[1] ;
 wire \hkspi.ldata[2] ;
 wire \hkspi.ldata[3] ;
 wire \hkspi.ldata[4] ;
 wire \hkspi.ldata[5] ;
 wire \hkspi.ldata[6] ;
 wire \hkspi.odata[1] ;
 wire \hkspi.odata[2] ;
 wire \hkspi.odata[3] ;
 wire \hkspi.odata[4] ;
 wire \hkspi.odata[5] ;
 wire \hkspi.odata[6] ;
 wire \hkspi.odata[7] ;
 wire \hkspi.pass_thru_mgmt ;
 wire \hkspi.pass_thru_mgmt_delay ;
 wire \hkspi.pass_thru_user ;
 wire \hkspi.pass_thru_user_delay ;
 wire \hkspi.pre_pass_thru_mgmt ;
 wire \hkspi.pre_pass_thru_user ;
 wire \hkspi.rdstb ;
 wire \hkspi.readmode ;
 wire \hkspi.sdoenb ;
 wire \hkspi.state[0] ;
 wire \hkspi.state[1] ;
 wire \hkspi.state[2] ;
 wire \hkspi.state[3] ;
 wire \hkspi.state[4] ;
 wire \hkspi.writemode ;
 wire \hkspi.wrstb ;
 wire hkspi_disable;
 wire irq_1_inputsrc;
 wire irq_2_inputsrc;
 wire \mgmt_gpio_data[0] ;
 wire \mgmt_gpio_data[10] ;
 wire \mgmt_gpio_data[13] ;
 wire \mgmt_gpio_data[14] ;
 wire \mgmt_gpio_data[15] ;
 wire \mgmt_gpio_data[1] ;
 wire \mgmt_gpio_data[32] ;
 wire \mgmt_gpio_data[33] ;
 wire \mgmt_gpio_data[35] ;
 wire \mgmt_gpio_data[36] ;
 wire \mgmt_gpio_data[37] ;
 wire \mgmt_gpio_data[6] ;
 wire \mgmt_gpio_data[8] ;
 wire \mgmt_gpio_data[9] ;
 wire \mgmt_gpio_data_buf[0] ;
 wire \mgmt_gpio_data_buf[10] ;
 wire \mgmt_gpio_data_buf[11] ;
 wire \mgmt_gpio_data_buf[12] ;
 wire \mgmt_gpio_data_buf[13] ;
 wire \mgmt_gpio_data_buf[14] ;
 wire \mgmt_gpio_data_buf[15] ;
 wire \mgmt_gpio_data_buf[16] ;
 wire \mgmt_gpio_data_buf[17] ;
 wire \mgmt_gpio_data_buf[18] ;
 wire \mgmt_gpio_data_buf[19] ;
 wire \mgmt_gpio_data_buf[1] ;
 wire \mgmt_gpio_data_buf[20] ;
 wire \mgmt_gpio_data_buf[21] ;
 wire \mgmt_gpio_data_buf[22] ;
 wire \mgmt_gpio_data_buf[23] ;
 wire \mgmt_gpio_data_buf[2] ;
 wire \mgmt_gpio_data_buf[3] ;
 wire \mgmt_gpio_data_buf[4] ;
 wire \mgmt_gpio_data_buf[5] ;
 wire \mgmt_gpio_data_buf[6] ;
 wire \mgmt_gpio_data_buf[7] ;
 wire \mgmt_gpio_data_buf[8] ;
 wire \mgmt_gpio_data_buf[9] ;
 wire \pad_count_1[0] ;
 wire \pad_count_1[1] ;
 wire \pad_count_1[2] ;
 wire \pad_count_1[3] ;
 wire \pad_count_1[4] ;
 wire \pad_count_2[0] ;
 wire \pad_count_2[1] ;
 wire \pad_count_2[2] ;
 wire \pad_count_2[3] ;
 wire \pad_count_2[4] ;
 wire \pad_count_2[5] ;
 wire reset_reg;
 wire serial_bb_clock;
 wire serial_bb_data_1;
 wire serial_bb_data_2;
 wire serial_bb_enable;
 wire serial_bb_load;
 wire serial_bb_resetn;
 wire serial_busy;
 wire serial_clock_pre;
 wire \serial_data_staging_1[0] ;
 wire \serial_data_staging_1[10] ;
 wire \serial_data_staging_1[11] ;
 wire \serial_data_staging_1[12] ;
 wire \serial_data_staging_1[1] ;
 wire \serial_data_staging_1[2] ;
 wire \serial_data_staging_1[3] ;
 wire \serial_data_staging_1[4] ;
 wire \serial_data_staging_1[5] ;
 wire \serial_data_staging_1[6] ;
 wire \serial_data_staging_1[7] ;
 wire \serial_data_staging_1[8] ;
 wire \serial_data_staging_1[9] ;
 wire \serial_data_staging_2[0] ;
 wire \serial_data_staging_2[10] ;
 wire \serial_data_staging_2[11] ;
 wire \serial_data_staging_2[12] ;
 wire \serial_data_staging_2[1] ;
 wire \serial_data_staging_2[2] ;
 wire \serial_data_staging_2[3] ;
 wire \serial_data_staging_2[4] ;
 wire \serial_data_staging_2[5] ;
 wire \serial_data_staging_2[6] ;
 wire \serial_data_staging_2[7] ;
 wire \serial_data_staging_2[8] ;
 wire \serial_data_staging_2[9] ;
 wire serial_load_pre;
 wire serial_resetn_pre;
 wire serial_xfer;
 wire trap_output_dest;
 wire \wbbd_addr[0] ;
 wire \wbbd_addr[1] ;
 wire \wbbd_addr[2] ;
 wire \wbbd_addr[3] ;
 wire \wbbd_addr[4] ;
 wire \wbbd_addr[5] ;
 wire \wbbd_addr[6] ;
 wire wbbd_busy;
 wire \wbbd_data[0] ;
 wire \wbbd_data[1] ;
 wire \wbbd_data[2] ;
 wire \wbbd_data[3] ;
 wire \wbbd_data[4] ;
 wire \wbbd_data[5] ;
 wire \wbbd_data[6] ;
 wire \wbbd_data[7] ;
 wire wbbd_sck;
 wire \wbbd_state[0] ;
 wire \wbbd_state[1] ;
 wire \wbbd_state[2] ;
 wire \wbbd_state[3] ;
 wire \wbbd_state[4] ;
 wire \wbbd_state[5] ;
 wire \wbbd_state[6] ;
 wire \wbbd_state[7] ;
 wire \wbbd_state[8] ;
 wire \wbbd_state[9] ;
 wire wbbd_write;
 wire \xfer_count[0] ;
 wire \xfer_count[1] ;
 wire \xfer_count[2] ;
 wire \xfer_count[3] ;
 wire \xfer_state[0] ;
 wire \xfer_state[1] ;
 wire \xfer_state[2] ;
 wire \xfer_state[3] ;
 wire net108;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net462;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_0_1_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_1_1_1_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_leaf_0_csclk;
 wire clknet_leaf_1_csclk;
 wire clknet_leaf_2_csclk;
 wire clknet_leaf_3_csclk;
 wire clknet_leaf_4_csclk;
 wire clknet_leaf_5_csclk;
 wire clknet_leaf_7_csclk;
 wire clknet_leaf_8_csclk;
 wire clknet_leaf_10_csclk;
 wire clknet_leaf_11_csclk;
 wire clknet_leaf_12_csclk;
 wire clknet_leaf_13_csclk;
 wire clknet_leaf_14_csclk;
 wire clknet_leaf_15_csclk;
 wire clknet_leaf_16_csclk;
 wire clknet_leaf_17_csclk;
 wire clknet_leaf_18_csclk;
 wire clknet_leaf_19_csclk;
 wire clknet_leaf_20_csclk;
 wire clknet_leaf_21_csclk;
 wire clknet_leaf_22_csclk;
 wire clknet_leaf_23_csclk;
 wire clknet_leaf_24_csclk;
 wire clknet_leaf_25_csclk;
 wire clknet_leaf_26_csclk;
 wire clknet_leaf_27_csclk;
 wire clknet_leaf_28_csclk;
 wire clknet_leaf_29_csclk;
 wire clknet_leaf_30_csclk;
 wire clknet_leaf_31_csclk;
 wire clknet_leaf_32_csclk;
 wire clknet_leaf_33_csclk;
 wire clknet_leaf_34_csclk;
 wire clknet_leaf_35_csclk;
 wire clknet_leaf_36_csclk;
 wire clknet_leaf_37_csclk;
 wire clknet_leaf_38_csclk;
 wire clknet_leaf_39_csclk;
 wire clknet_leaf_40_csclk;
 wire clknet_leaf_42_csclk;
 wire clknet_leaf_43_csclk;
 wire clknet_leaf_44_csclk;
 wire clknet_leaf_45_csclk;
 wire clknet_leaf_46_csclk;
 wire clknet_leaf_47_csclk;
 wire clknet_leaf_48_csclk;
 wire clknet_leaf_49_csclk;
 wire clknet_leaf_50_csclk;
 wire clknet_leaf_51_csclk;
 wire clknet_leaf_52_csclk;
 wire clknet_leaf_53_csclk;
 wire clknet_leaf_54_csclk;
 wire clknet_leaf_55_csclk;
 wire clknet_leaf_56_csclk;
 wire clknet_leaf_57_csclk;
 wire clknet_leaf_58_csclk;
 wire clknet_leaf_59_csclk;
 wire clknet_leaf_60_csclk;
 wire clknet_leaf_61_csclk;
 wire clknet_leaf_62_csclk;
 wire clknet_leaf_63_csclk;
 wire clknet_leaf_64_csclk;
 wire clknet_leaf_65_csclk;
 wire clknet_leaf_67_csclk;
 wire clknet_leaf_68_csclk;
 wire clknet_leaf_69_csclk;
 wire clknet_leaf_70_csclk;
 wire clknet_leaf_71_csclk;
 wire clknet_leaf_72_csclk;
 wire clknet_leaf_73_csclk;
 wire clknet_leaf_74_csclk;
 wire clknet_leaf_75_csclk;
 wire clknet_leaf_76_csclk;
 wire clknet_leaf_77_csclk;
 wire clknet_leaf_78_csclk;
 wire clknet_0_csclk;
 wire clknet_1_0_0_csclk;
 wire clknet_1_0_1_csclk;
 wire clknet_1_1_0_csclk;
 wire clknet_1_1_1_csclk;
 wire clknet_2_0_0_csclk;
 wire clknet_2_1_0_csclk;
 wire clknet_2_2_0_csclk;
 wire clknet_2_3_0_csclk;
 wire clknet_3_0_0_csclk;
 wire clknet_3_1_0_csclk;
 wire clknet_3_2_0_csclk;
 wire clknet_3_3_0_csclk;
 wire clknet_3_4_0_csclk;
 wire clknet_3_5_0_csclk;
 wire clknet_3_6_0_csclk;
 wire clknet_3_7_0_csclk;
 wire clknet_opt_1_0_csclk;
 wire clknet_opt_2_0_csclk;
 wire clknet_opt_3_0_csclk;
 wire clknet_opt_4_0_csclk;
 wire clknet_0__1132_;
 wire clknet_1_0__leaf__1132_;
 wire clknet_1_1__leaf__1132_;
 wire clknet_0_wbbd_sck;
 wire clknet_1_0__leaf_wbbd_sck;
 wire clknet_1_1__leaf_wbbd_sck;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire [4:0] clknet_0_mgmt_gpio_in;
 wire [4:0] clknet_1_0_0_mgmt_gpio_in;
 wire [4:0] clknet_1_1_0_mgmt_gpio_in;
 wire [4:0] clknet_2_0_0_mgmt_gpio_in;
 wire [4:0] clknet_2_1_0_mgmt_gpio_in;
 wire [4:0] clknet_2_2_0_mgmt_gpio_in;
 wire [4:0] clknet_2_3_0_mgmt_gpio_in;

 sky130_fd_sc_hd__inv_2 _3191_ (.A(\hkspi.addr[0] ),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _3192_ (.A(\hkspi.pre_pass_thru_mgmt ),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _3193_ (.A(\wbbd_state[0] ),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _3194_ (.A(\gpio_configure[3][3] ),
    .Y(net206));
 sky130_fd_sc_hd__clkinv_8 _3195_ (.A(\wbbd_state[6] ),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _3196_ (.A(\hkspi.state[2] ),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_8 _3197_ (.A(net407),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _3198_ (.A(\xfer_state[0] ),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _3199_ (.A(\xfer_state[3] ),
    .Y(_0821_));
 sky130_fd_sc_hd__clkinv_8 _3200_ (.A(\xfer_state[2] ),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _3201_ (.A(\hkspi.state[4] ),
    .Y(_0823_));
 sky130_fd_sc_hd__clkinv_2 _3202_ (.A(net38),
    .Y(_0824_));
 sky130_fd_sc_hd__clkinv_2 _3203_ (.A(\gpio_configure[37][3] ),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _3204_ (.A(\gpio_configure[36][3] ),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _3205_ (.A(\gpio_configure[35][3] ),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_2 _3206_ (.A(\gpio_configure[34][3] ),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _3207_ (.A(\gpio_configure[33][3] ),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(\gpio_configure[32][3] ),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _3209_ (.A(\gpio_configure[31][3] ),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _3210_ (.A(\gpio_configure[30][3] ),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _3211_ (.A(\gpio_configure[29][3] ),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _3212_ (.A(\gpio_configure[28][3] ),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _3213_ (.A(\gpio_configure[27][3] ),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _3214_ (.A(\gpio_configure[26][3] ),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _3215_ (.A(\gpio_configure[25][3] ),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(\gpio_configure[24][3] ),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(\gpio_configure[23][3] ),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _3218_ (.A(\gpio_configure[22][3] ),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _3219_ (.A(\gpio_configure[21][3] ),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _3220_ (.A(\gpio_configure[20][3] ),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _3221_ (.A(\gpio_configure[19][3] ),
    .Y(net185));
 sky130_fd_sc_hd__clkinv_2 _3222_ (.A(\gpio_configure[18][3] ),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _3223_ (.A(\gpio_configure[17][3] ),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _3224_ (.A(\gpio_configure[16][3] ),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _3225_ (.A(\gpio_configure[15][3] ),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _3226_ (.A(\gpio_configure[14][3] ),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _3227_ (.A(\gpio_configure[13][3] ),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _3228_ (.A(\gpio_configure[12][3] ),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _3229_ (.A(\gpio_configure[11][3] ),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _3230_ (.A(\gpio_configure[10][3] ),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _3231_ (.A(\gpio_configure[9][3] ),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _3232_ (.A(\gpio_configure[8][3] ),
    .Y(net211));
 sky130_fd_sc_hd__clkinv_2 _3233_ (.A(\gpio_configure[7][3] ),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _3234_ (.A(\gpio_configure[6][3] ),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _3235_ (.A(\gpio_configure[5][3] ),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _3236_ (.A(\gpio_configure[4][3] ),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _3237_ (.A(\gpio_configure[2][3] ),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _3238_ (.A(\gpio_configure[1][3] ),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_2 _3239_ (.A(\gpio_configure[0][3] ),
    .Y(_0829_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__inv_8 _3241_ (.A(\pad_count_1[4] ),
    .Y(_0830_));
 sky130_fd_sc_hd__clkinv_4 _3242_ (.A(net110),
    .Y(_0831_));
 sky130_fd_sc_hd__clkinv_4 _3243_ (.A(net99),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_8 _3244_ (.A(net124),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_6 _3245_ (.A(net121),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_6 _3246_ (.A(net128),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_4 _3247_ (.A(net459),
    .Y(_0836_));
 sky130_fd_sc_hd__or3_4 _3248_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_0837_));
 sky130_fd_sc_hd__nand2b_1 _3249_ (.A_N(net409),
    .B(net565),
    .Y(_0838_));
 sky130_fd_sc_hd__a21bo_2 _3250_ (.A1(net573),
    .A2(net409),
    .B1_N(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_8 _3251_ (.A0(net520),
    .A1(net635),
    .S(net406),
    .X(_0840_));
 sky130_fd_sc_hd__inv_2 _3252_ (.A(net521),
    .Y(_0841_));
 sky130_fd_sc_hd__mux2_2 _3253_ (.A0(\hkspi.addr[5] ),
    .A1(net565),
    .S(net409),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_8 _3254_ (.A0(net566),
    .A1(net606),
    .S(net406),
    .X(_0843_));
 sky130_fd_sc_hd__and2b_2 _3255_ (.A_N(net409),
    .B(net684),
    .X(_0844_));
 sky130_fd_sc_hd__a21oi_4 _3256_ (.A1(net512),
    .A2(net409),
    .B1(net685),
    .Y(_0845_));
 sky130_fd_sc_hd__a21o_1 _3257_ (.A1(net653),
    .A2(net409),
    .B1(net512),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_4 _3258_ (.A0(net654),
    .A1(\wbbd_addr[6] ),
    .S(net406),
    .X(_0847_));
 sky130_fd_sc_hd__o21ai_4 _3259_ (.A1(net406),
    .A2(net513),
    .B1(net655),
    .Y(_0848_));
 sky130_fd_sc_hd__or3_4 _3260_ (.A(net637),
    .B(net608),
    .C(net657),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(net486),
    .A1(net478),
    .S(net409),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_8 _3262_ (.A0(net487),
    .A1(net583),
    .S(net406),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(net573),
    .A1(net486),
    .S(net409),
    .X(_0852_));
 sky130_fd_sc_hd__and2b_4 _3264_ (.A_N(net406),
    .B(net574),
    .X(_0853_));
 sky130_fd_sc_hd__a21o_4 _3265_ (.A1(net406),
    .A2(net748),
    .B1(net575),
    .X(_0854_));
 sky130_fd_sc_hd__a21oi_4 _3266_ (.A1(net406),
    .A2(net550),
    .B1(net575),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_2 _3267_ (.A(net488),
    .B(net551),
    .Y(_0856_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(net478),
    .A1(net542),
    .S(net409),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_8 _3269_ (.A0(net479),
    .A1(net787),
    .S(net406),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(net542),
    .A1(net58),
    .S(net409),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_8 _3271_ (.A0(net543),
    .A1(net819),
    .S(net406),
    .X(_0860_));
 sky130_fd_sc_hd__or2_4 _3272_ (.A(net480),
    .B(net544),
    .X(_0861_));
 sky130_fd_sc_hd__or2_4 _3273_ (.A(net552),
    .B(net481),
    .X(_0862_));
 sky130_fd_sc_hd__nor2_8 _3274_ (.A(net360),
    .B(net553),
    .Y(_0863_));
 sky130_fd_sc_hd__or3_4 _3275_ (.A(_0841_),
    .B(net608),
    .C(net657),
    .X(_0864_));
 sky130_fd_sc_hd__nor2_8 _3276_ (.A(net553),
    .B(net357),
    .Y(_0865_));
 sky130_fd_sc_hd__o21bai_4 _3277_ (.A1(net406),
    .A2(net513),
    .B1_N(net655),
    .Y(_0866_));
 sky130_fd_sc_hd__or2_1 _3278_ (.A(net567),
    .B(net687),
    .X(_0867_));
 sky130_fd_sc_hd__or2_4 _3279_ (.A(net637),
    .B(net568),
    .X(_0868_));
 sky130_fd_sc_hd__inv_2 _3280_ (.A(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_2 _3281_ (.A(net480),
    .B(net544),
    .Y(_0870_));
 sky130_fd_sc_hd__or2_4 _3282_ (.A(net552),
    .B(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_8 _3283_ (.A(net356),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__or2_4 _3284_ (.A(net585),
    .B(net551),
    .X(_0873_));
 sky130_fd_sc_hd__or2_4 _3285_ (.A(net481),
    .B(net586),
    .X(_0874_));
 sky130_fd_sc_hd__nor2_8 _3286_ (.A(net515),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__a22o_1 _3287_ (.A1(net33),
    .A2(_0872_),
    .B1(_0875_),
    .B2(\gpio_configure[29][7] ),
    .X(_0876_));
 sky130_fd_sc_hd__nand2b_4 _3288_ (.A_N(net544),
    .B(net480),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_2 _3289_ (.A(net488),
    .B(net576),
    .Y(_0878_));
 sky130_fd_sc_hd__or2_4 _3290_ (.A(net545),
    .B(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_8 _3291_ (.A(net360),
    .B(net546),
    .Y(_0880_));
 sky130_fd_sc_hd__or3_4 _3292_ (.A(net488),
    .B(net576),
    .C(net481),
    .X(_0881_));
 sky130_fd_sc_hd__nand2b_1 _3293_ (.A_N(net687),
    .B(net567),
    .Y(_0882_));
 sky130_fd_sc_hd__or2_4 _3294_ (.A(net521),
    .B(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_8 _3295_ (.A(net489),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__a221o_1 _3296_ (.A1(\gpio_configure[24][7] ),
    .A2(_0880_),
    .B1(_0884_),
    .B2(\gpio_configure[1][7] ),
    .C1(_0876_),
    .X(_0885_));
 sky130_fd_sc_hd__a221o_1 _3297_ (.A1(\gpio_configure[19][7] ),
    .A2(_0863_),
    .B1(_0865_),
    .B2(\gpio_configure[27][7] ),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_8 _3298_ (.A(net357),
    .B(net578),
    .Y(_0887_));
 sky130_fd_sc_hd__nor2_8 _3299_ (.A(net360),
    .B(net578),
    .Y(_0888_));
 sky130_fd_sc_hd__a22o_1 _3300_ (.A1(\gpio_configure[25][7] ),
    .A2(_0887_),
    .B1(_0888_),
    .B2(\gpio_configure[17][7] ),
    .X(_0889_));
 sky130_fd_sc_hd__nor2_8 _3301_ (.A(net609),
    .B(_0874_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_8 _3302_ (.A(_0862_),
    .B(net356),
    .Y(_0891_));
 sky130_fd_sc_hd__a221o_2 _3303_ (.A1(\gpio_configure[21][7] ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(net28),
    .C1(_0889_),
    .X(_0892_));
 sky130_fd_sc_hd__or2_4 _3304_ (.A(_0841_),
    .B(_0882_),
    .X(_0893_));
 sky130_fd_sc_hd__nor2_8 _3305_ (.A(_0874_),
    .B(net354),
    .Y(_0894_));
 sky130_fd_sc_hd__nor2_8 _3306_ (.A(net578),
    .B(_0893_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_4 _3307_ (.A(net481),
    .B(_0878_),
    .X(_0896_));
 sky130_fd_sc_hd__inv_2 _3308_ (.A(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__or3b_4 _3309_ (.A(net637),
    .B(net514),
    .C_N(net567),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_8 _3310_ (.A(net482),
    .B(net358),
    .Y(_0899_));
 sky130_fd_sc_hd__nor2_8 _3311_ (.A(net357),
    .B(net546),
    .Y(_0900_));
 sky130_fd_sc_hd__a22o_1 _3312_ (.A1(net42),
    .A2(_0899_),
    .B1(_0900_),
    .B2(\gpio_configure[32][7] ),
    .X(_0901_));
 sky130_fd_sc_hd__a221o_4 _3313_ (.A1(\gpio_configure[13][7] ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\gpio_configure[9][7] ),
    .C1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__or2_4 _3314_ (.A(_0841_),
    .B(net568),
    .X(_0903_));
 sky130_fd_sc_hd__nor2_8 _3315_ (.A(net546),
    .B(net569),
    .Y(_0904_));
 sky130_fd_sc_hd__or3_4 _3316_ (.A(net585),
    .B(net576),
    .C(net545),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_8 _3317_ (.A(net357),
    .B(net749),
    .Y(_0906_));
 sky130_fd_sc_hd__a22o_1 _3318_ (.A1(\gpio_configure[0][7] ),
    .A2(_0904_),
    .B1(_0906_),
    .B2(\gpio_configure[26][7] ),
    .X(_0907_));
 sky130_fd_sc_hd__or2_4 _3319_ (.A(net552),
    .B(net545),
    .X(_0908_));
 sky130_fd_sc_hd__nor2_8 _3320_ (.A(net356),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__or2_4 _3321_ (.A(net586),
    .B(net545),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_8 _3322_ (.A(net359),
    .B(net587),
    .Y(_0911_));
 sky130_fd_sc_hd__a221o_1 _3323_ (.A1(net10),
    .A2(_0909_),
    .B1(_0911_),
    .B2(net60),
    .C1(_0907_),
    .X(_0912_));
 sky130_fd_sc_hd__nor2_8 _3324_ (.A(net546),
    .B(_0883_),
    .Y(_0913_));
 sky130_fd_sc_hd__nor2_8 _3325_ (.A(_0883_),
    .B(net482),
    .Y(_0914_));
 sky130_fd_sc_hd__a22o_1 _3326_ (.A1(\gpio_configure[8][7] ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\gpio_configure[7][7] ),
    .X(_0915_));
 sky130_fd_sc_hd__nor2_8 _3327_ (.A(_0893_),
    .B(net587),
    .Y(_0916_));
 sky130_fd_sc_hd__or2_4 _3328_ (.A(_0870_),
    .B(net586),
    .X(_0917_));
 sky130_fd_sc_hd__nor2_8 _3329_ (.A(net358),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__a221o_4 _3330_ (.A1(\gpio_configure[14][7] ),
    .A2(_0916_),
    .B1(_0918_),
    .B2(net51),
    .C1(_0915_),
    .X(_0919_));
 sky130_fd_sc_hd__or4_1 _3331_ (.A(_0892_),
    .B(_0902_),
    .C(_0912_),
    .D(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__or2_4 _3332_ (.A(_0870_),
    .B(_0878_),
    .X(_0921_));
 sky130_fd_sc_hd__nor2_8 _3333_ (.A(_0868_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__nor2_8 _3334_ (.A(net609),
    .B(net482),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_8 _3335_ (.A(net356),
    .B(net546),
    .Y(_0924_));
 sky130_fd_sc_hd__a22o_1 _3336_ (.A1(\gpio_configure[23][7] ),
    .A2(_0923_),
    .B1(_0924_),
    .B2(net281),
    .X(_0925_));
 sky130_fd_sc_hd__a21o_2 _3337_ (.A1(net290),
    .A2(_0922_),
    .B1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__nor2_8 _3338_ (.A(_0883_),
    .B(net587),
    .Y(_0927_));
 sky130_fd_sc_hd__nor2_8 _3339_ (.A(net360),
    .B(net587),
    .Y(_0928_));
 sky130_fd_sc_hd__a22o_1 _3340_ (.A1(\gpio_configure[6][7] ),
    .A2(_0927_),
    .B1(_0928_),
    .B2(\gpio_configure[22][7] ),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_8 _3341_ (.A(net357),
    .B(net587),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2b_4 _3342_ (.A_N(net789),
    .B(net544),
    .Y(_0931_));
 sky130_fd_sc_hd__or2_4 _3343_ (.A(_0878_),
    .B(net790),
    .X(_0932_));
 sky130_fd_sc_hd__nor2_8 _3344_ (.A(_0868_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__a221o_1 _3345_ (.A1(\gpio_configure[30][7] ),
    .A2(_0930_),
    .B1(_0933_),
    .B2(net298),
    .C1(_0929_),
    .X(_0934_));
 sky130_fd_sc_hd__nor2_8 _3346_ (.A(net359),
    .B(_0908_),
    .Y(_0935_));
 sky130_fd_sc_hd__nor2_8 _3347_ (.A(net355),
    .B(_0908_),
    .Y(_0936_));
 sky130_fd_sc_hd__a22o_1 _3348_ (.A1(\gpio_configure[36][7] ),
    .A2(_0935_),
    .B1(_0936_),
    .B2(\gpio_configure[4][7] ),
    .X(_0937_));
 sky130_fd_sc_hd__nor2_8 _3349_ (.A(net609),
    .B(_0905_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_8 _3350_ (.A(_0874_),
    .B(net358),
    .Y(_0939_));
 sky130_fd_sc_hd__a221o_4 _3351_ (.A1(\gpio_configure[18][7] ),
    .A2(_0938_),
    .B1(_0939_),
    .B2(\gpio_configure[37][7] ),
    .C1(_0937_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_8 _3352_ (.A(_0874_),
    .B(net355),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_8 _3353_ (.A(net553),
    .B(_0883_),
    .Y(_0942_));
 sky130_fd_sc_hd__a22o_1 _3354_ (.A1(\gpio_configure[5][7] ),
    .A2(_0941_),
    .B1(_0942_),
    .B2(\gpio_configure[3][7] ),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_8 _3355_ (.A(net357),
    .B(net482),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_8 _3356_ (.A(_0893_),
    .B(net749),
    .Y(_0945_));
 sky130_fd_sc_hd__a221o_2 _3357_ (.A1(\gpio_configure[31][7] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(\gpio_configure[10][7] ),
    .C1(_0943_),
    .X(_0946_));
 sky130_fd_sc_hd__nor2_8 _3358_ (.A(net359),
    .B(net749),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_8 _3359_ (.A(net609),
    .B(_0908_),
    .Y(_0948_));
 sky130_fd_sc_hd__a22o_1 _3360_ (.A1(\gpio_configure[34][7] ),
    .A2(_0947_),
    .B1(_0948_),
    .B2(\gpio_configure[20][7] ),
    .X(_0949_));
 sky130_fd_sc_hd__nor2_8 _3361_ (.A(net359),
    .B(_0932_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_8 _3362_ (.A(net553),
    .B(_0893_),
    .Y(_0951_));
 sky130_fd_sc_hd__a221o_1 _3363_ (.A1(net70),
    .A2(_0950_),
    .B1(_0951_),
    .B2(\gpio_configure[11][7] ),
    .C1(_0949_),
    .X(_0952_));
 sky130_fd_sc_hd__nor2_8 _3364_ (.A(net357),
    .B(_0908_),
    .Y(_0953_));
 sky130_fd_sc_hd__nor2_8 _3365_ (.A(_0862_),
    .B(net522),
    .Y(_0954_));
 sky130_fd_sc_hd__a22o_1 _3366_ (.A1(\gpio_configure[28][7] ),
    .A2(_0953_),
    .B1(_0954_),
    .B2(\gpio_configure[35][7] ),
    .X(_0955_));
 sky130_fd_sc_hd__or2_4 _3367_ (.A(net552),
    .B(net790),
    .X(_0956_));
 sky130_fd_sc_hd__nor2_8 _3368_ (.A(net356),
    .B(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_8 _3369_ (.A(_0893_),
    .B(net482),
    .Y(_0958_));
 sky130_fd_sc_hd__a221o_1 _3370_ (.A1(net19),
    .A2(_0957_),
    .B1(_0958_),
    .B2(\gpio_configure[15][7] ),
    .C1(_0955_),
    .X(_0959_));
 sky130_fd_sc_hd__nor2_8 _3371_ (.A(net578),
    .B(net359),
    .Y(_0960_));
 sky130_fd_sc_hd__nor2_8 _3372_ (.A(net546),
    .B(_0893_),
    .Y(_0961_));
 sky130_fd_sc_hd__a22o_1 _3373_ (.A1(\gpio_configure[33][7] ),
    .A2(_0960_),
    .B1(_0961_),
    .B2(\gpio_configure[16][7] ),
    .X(_0962_));
 sky130_fd_sc_hd__nor2_8 _3374_ (.A(_0883_),
    .B(net749),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2_8 _3375_ (.A(net354),
    .B(_0908_),
    .Y(_0964_));
 sky130_fd_sc_hd__a221o_4 _3376_ (.A1(\gpio_configure[2][7] ),
    .A2(_0963_),
    .B1(_0964_),
    .B2(\gpio_configure[12][7] ),
    .C1(_0962_),
    .X(_0965_));
 sky130_fd_sc_hd__or4_1 _3377_ (.A(_0946_),
    .B(_0952_),
    .C(_0959_),
    .D(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__or4_2 _3378_ (.A(_0926_),
    .B(_0934_),
    .C(_0940_),
    .D(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__or3_4 _3379_ (.A(_0886_),
    .B(_0920_),
    .C(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__nand2_8 _3380_ (.A(\hkspi.readmode ),
    .B(\hkspi.state[2] ),
    .Y(_0969_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(_0968_),
    .A1(\hkspi.ldata[6] ),
    .S(_0837_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(_0970_),
    .A1(\hkspi.SDO ),
    .S(_0969_),
    .X(_0386_));
 sky130_fd_sc_hd__or3_4 _3383_ (.A(net585),
    .B(net576),
    .C(_0870_),
    .X(_0971_));
 sky130_fd_sc_hd__nor2_8 _3384_ (.A(net569),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux2_8 _3385_ (.A0(\serial_data_staging_2[12] ),
    .A1(serial_bb_data_2),
    .S(serial_bb_enable),
    .X(net309));
 sky130_fd_sc_hd__nor2_8 _3386_ (.A(_0868_),
    .B(_0905_),
    .Y(_0973_));
 sky130_fd_sc_hd__a22o_1 _3387_ (.A1(net41),
    .A2(_0899_),
    .B1(_0914_),
    .B2(\gpio_configure[7][6] ),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _3388_ (.A1(\gpio_configure[36][6] ),
    .A2(_0935_),
    .B1(_0950_),
    .B2(net69),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _3389_ (.A1(net32),
    .A2(_0872_),
    .B1(_0880_),
    .B2(\gpio_configure[24][6] ),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _3390_ (.A1(\gpio_configure[4][6] ),
    .A2(_0936_),
    .B1(_0961_),
    .B2(\gpio_configure[16][6] ),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _3391_ (.A1(\gpio_configure[21][6] ),
    .A2(_0890_),
    .B1(_0944_),
    .B2(\gpio_configure[31][6] ),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _3392_ (.A1(\gpio_configure[29][6] ),
    .A2(_0875_),
    .B1(_0948_),
    .B2(\gpio_configure[20][6] ),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _3393_ (.A1(\gpio_configure[13][6] ),
    .A2(_0894_),
    .B1(_0954_),
    .B2(\gpio_configure[35][6] ),
    .C1(_0977_),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _3394_ (.A1(\gpio_configure[25][6] ),
    .A2(_0887_),
    .B1(_0938_),
    .B2(\gpio_configure[18][6] ),
    .X(_0981_));
 sky130_fd_sc_hd__a221o_1 _3395_ (.A1(\gpio_configure[1][6] ),
    .A2(_0884_),
    .B1(_0923_),
    .B2(\gpio_configure[23][6] ),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a221o_4 _3396_ (.A1(\gpio_configure[10][6] ),
    .A2(_0945_),
    .B1(_0964_),
    .B2(\gpio_configure[12][6] ),
    .C1(_0974_),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_4 _3397_ (.A1(net9),
    .A2(_0909_),
    .B1(_0928_),
    .B2(\gpio_configure[22][6] ),
    .C1(_0979_),
    .X(_0984_));
 sky130_fd_sc_hd__or4_2 _3398_ (.A(_0980_),
    .B(_0982_),
    .C(_0983_),
    .D(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__a221o_1 _3399_ (.A1(\gpio_configure[30][6] ),
    .A2(_0930_),
    .B1(_0953_),
    .B2(\gpio_configure[28][6] ),
    .C1(_0978_),
    .X(_0986_));
 sky130_fd_sc_hd__a221o_2 _3400_ (.A1(\gpio_configure[26][6] ),
    .A2(_0906_),
    .B1(_0922_),
    .B2(net289),
    .C1(_0976_),
    .X(_0987_));
 sky130_fd_sc_hd__a211o_1 _3401_ (.A1(\gpio_configure[15][6] ),
    .A2(_0958_),
    .B1(_0986_),
    .C1(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__a221o_4 _3402_ (.A1(\gpio_configure[3][6] ),
    .A2(_0942_),
    .B1(_0951_),
    .B2(\gpio_configure[11][6] ),
    .C1(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _3403_ (.A1(\gpio_configure[34][6] ),
    .A2(_0947_),
    .B1(_0963_),
    .B2(\gpio_configure[2][6] ),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_4 _3404_ (.A1(\gpio_configure[32][6] ),
    .A2(_0900_),
    .B1(_0939_),
    .B2(\gpio_configure[37][6] ),
    .X(_0991_));
 sky130_fd_sc_hd__a221o_1 _3405_ (.A1(\gpio_configure[19][6] ),
    .A2(_0863_),
    .B1(_0933_),
    .B2(net297),
    .C1(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__a2111o_1 _3406_ (.A1(\gpio_configure[6][6] ),
    .A2(_0927_),
    .B1(_0973_),
    .C1(_0990_),
    .D1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a22o_1 _3407_ (.A1(\gpio_configure[27][6] ),
    .A2(_0865_),
    .B1(_0913_),
    .B2(\gpio_configure[8][6] ),
    .X(_0994_));
 sky130_fd_sc_hd__a221o_1 _3408_ (.A1(\gpio_configure[0][6] ),
    .A2(_0904_),
    .B1(_0918_),
    .B2(net50),
    .C1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _3409_ (.A1(\gpio_configure[5][6] ),
    .A2(_0941_),
    .B1(_0972_),
    .B2(net309),
    .X(_0996_));
 sky130_fd_sc_hd__a221o_2 _3410_ (.A1(\gpio_configure[9][6] ),
    .A2(_0895_),
    .B1(_0916_),
    .B2(\gpio_configure[14][6] ),
    .C1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__a221o_1 _3411_ (.A1(\gpio_configure[17][6] ),
    .A2(_0888_),
    .B1(_0924_),
    .B2(net280),
    .C1(_0975_),
    .X(_0998_));
 sky130_fd_sc_hd__a22o_1 _3412_ (.A1(net27),
    .A2(_0891_),
    .B1(_0960_),
    .B2(\gpio_configure[33][6] ),
    .X(_0999_));
 sky130_fd_sc_hd__a221o_1 _3413_ (.A1(net59),
    .A2(_0911_),
    .B1(_0957_),
    .B2(net18),
    .C1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__or4_1 _3414_ (.A(_0995_),
    .B(_0997_),
    .C(_0998_),
    .D(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__or4_4 _3415_ (.A(_0985_),
    .B(_0989_),
    .C(_0993_),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(_1002_),
    .A1(\hkspi.ldata[5] ),
    .S(_0837_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(_1003_),
    .A1(\hkspi.ldata[6] ),
    .S(_0969_),
    .X(_0385_));
 sky130_fd_sc_hd__a22o_1 _3418_ (.A1(\gpio_configure[34][5] ),
    .A2(_0947_),
    .B1(_0960_),
    .B2(\gpio_configure[33][5] ),
    .X(_1004_));
 sky130_fd_sc_hd__or2_4 _3419_ (.A(net586),
    .B(net790),
    .X(_1005_));
 sky130_fd_sc_hd__nor2_8 _3420_ (.A(net358),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__or3_4 _3421_ (.A(net585),
    .B(net576),
    .C(net790),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_8 _3422_ (.A(net569),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__mux2_8 _3423_ (.A0(\serial_data_staging_1[12] ),
    .A1(serial_bb_data_1),
    .S(serial_bb_enable),
    .X(net308));
 sky130_fd_sc_hd__a22o_1 _3424_ (.A1(\gpio_configure[13][5] ),
    .A2(_0894_),
    .B1(_0941_),
    .B2(\gpio_configure[5][5] ),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _3425_ (.A1(\gpio_configure[10][5] ),
    .A2(_0945_),
    .B1(_0963_),
    .B2(\gpio_configure[2][5] ),
    .X(_1010_));
 sky130_fd_sc_hd__a22o_4 _3426_ (.A1(\gpio_configure[25][5] ),
    .A2(_0887_),
    .B1(_0900_),
    .B2(\gpio_configure[32][5] ),
    .X(_1011_));
 sky130_fd_sc_hd__a221o_1 _3427_ (.A1(net288),
    .A2(_0922_),
    .B1(_0928_),
    .B2(\gpio_configure[22][5] ),
    .C1(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_2 _3428_ (.A1(net31),
    .A2(_0872_),
    .B1(_0924_),
    .B2(net279),
    .X(_1013_));
 sky130_fd_sc_hd__a221o_1 _3429_ (.A1(\gpio_configure[23][5] ),
    .A2(_0923_),
    .B1(_0938_),
    .B2(\gpio_configure[18][5] ),
    .C1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_2 _3430_ (.A1(net296),
    .A2(_0933_),
    .B1(_0957_),
    .B2(net17),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_2 _3431_ (.A1(\gpio_configure[1][5] ),
    .A2(_0884_),
    .B1(_1006_),
    .B2(net66),
    .X(_1016_));
 sky130_fd_sc_hd__a221o_1 _3432_ (.A1(\gpio_configure[0][5] ),
    .A2(_0904_),
    .B1(_0906_),
    .B2(\gpio_configure[26][5] ),
    .C1(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__a221o_2 _3433_ (.A1(\gpio_configure[29][5] ),
    .A2(_0875_),
    .B1(_0890_),
    .B2(\gpio_configure[21][5] ),
    .C1(_1010_),
    .X(_1018_));
 sky130_fd_sc_hd__a221o_1 _3434_ (.A1(net40),
    .A2(_0899_),
    .B1(_0913_),
    .B2(\gpio_configure[8][5] ),
    .C1(_1004_),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_4 _3435_ (.A1(net57),
    .A2(_0911_),
    .B1(_0939_),
    .B2(\gpio_configure[37][5] ),
    .C1(_1009_),
    .X(_1020_));
 sky130_fd_sc_hd__or4_4 _3436_ (.A(_1017_),
    .B(_1018_),
    .C(_1019_),
    .D(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__a22o_1 _3437_ (.A1(\gpio_configure[27][5] ),
    .A2(_0865_),
    .B1(_0972_),
    .B2(net308),
    .X(_1022_));
 sky130_fd_sc_hd__a221o_1 _3438_ (.A1(\gpio_configure[17][5] ),
    .A2(_0888_),
    .B1(_0944_),
    .B2(\gpio_configure[31][5] ),
    .C1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_4 _3439_ (.A1(\gpio_configure[3][5] ),
    .A2(_0942_),
    .B1(_0961_),
    .B2(\gpio_configure[16][5] ),
    .X(_1024_));
 sky130_fd_sc_hd__a221o_1 _3440_ (.A1(\gpio_configure[30][5] ),
    .A2(_0930_),
    .B1(_0951_),
    .B2(\gpio_configure[11][5] ),
    .C1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a22o_4 _3441_ (.A1(\gpio_configure[14][5] ),
    .A2(_0916_),
    .B1(_0950_),
    .B2(net68),
    .X(_1026_));
 sky130_fd_sc_hd__a221o_4 _3442_ (.A1(\gpio_configure[36][5] ),
    .A2(_0935_),
    .B1(_0964_),
    .B2(\gpio_configure[12][5] ),
    .C1(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a221o_1 _3443_ (.A1(\gpio_configure[6][5] ),
    .A2(_0927_),
    .B1(_0953_),
    .B2(\gpio_configure[28][5] ),
    .C1(_1015_),
    .X(_1028_));
 sky130_fd_sc_hd__a22o_4 _3444_ (.A1(net25),
    .A2(_0891_),
    .B1(_0909_),
    .B2(net8),
    .X(_1029_));
 sky130_fd_sc_hd__a221o_1 _3445_ (.A1(\gpio_configure[19][5] ),
    .A2(_0863_),
    .B1(_0914_),
    .B2(\gpio_configure[7][5] ),
    .C1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_1 _3446_ (.A1(\gpio_configure[9][5] ),
    .A2(_0895_),
    .B1(_1008_),
    .B2(net263),
    .X(_1031_));
 sky130_fd_sc_hd__a221o_1 _3447_ (.A1(\gpio_configure[20][5] ),
    .A2(_0948_),
    .B1(_0958_),
    .B2(\gpio_configure[15][5] ),
    .C1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__a22o_1 _3448_ (.A1(\gpio_configure[24][5] ),
    .A2(_0880_),
    .B1(_0936_),
    .B2(\gpio_configure[4][5] ),
    .X(_1033_));
 sky130_fd_sc_hd__a221o_4 _3449_ (.A1(net49),
    .A2(_0918_),
    .B1(_0954_),
    .B2(\gpio_configure[35][5] ),
    .C1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__or4_2 _3450_ (.A(_1012_),
    .B(_1014_),
    .C(_1032_),
    .D(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__or4_1 _3451_ (.A(_1027_),
    .B(_1028_),
    .C(_1030_),
    .D(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or4_4 _3452_ (.A(_1021_),
    .B(_1023_),
    .C(_1025_),
    .D(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(_1037_),
    .A1(\hkspi.ldata[4] ),
    .S(_0837_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(_1038_),
    .A1(\hkspi.ldata[5] ),
    .S(_0969_),
    .X(_0384_));
 sky130_fd_sc_hd__nor2_8 _3455_ (.A(_0893_),
    .B(_1007_),
    .Y(_1039_));
 sky130_fd_sc_hd__a22o_1 _3456_ (.A1(net16),
    .A2(_0957_),
    .B1(_1039_),
    .B2(\gpio_configure[10][12] ),
    .X(_1040_));
 sky130_fd_sc_hd__nor2_8 _3457_ (.A(_0893_),
    .B(_0932_),
    .Y(_1041_));
 sky130_fd_sc_hd__a221o_1 _3458_ (.A1(\gpio_configure[18][4] ),
    .A2(_0938_),
    .B1(_1041_),
    .B2(\gpio_configure[16][12] ),
    .C1(_1040_),
    .X(_1042_));
 sky130_fd_sc_hd__nor2_8 _3459_ (.A(net357),
    .B(_0932_),
    .Y(_1043_));
 sky130_fd_sc_hd__nor2_8 _3460_ (.A(net360),
    .B(_0917_),
    .Y(_1044_));
 sky130_fd_sc_hd__a22o_2 _3461_ (.A1(\gpio_configure[32][12] ),
    .A2(_1043_),
    .B1(_1044_),
    .B2(\gpio_configure[23][12] ),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_8 _3462_ (.A(net354),
    .B(_0917_),
    .Y(_1046_));
 sky130_fd_sc_hd__a221o_1 _3463_ (.A1(\gpio_configure[6][4] ),
    .A2(_0927_),
    .B1(_1046_),
    .B2(\gpio_configure[15][12] ),
    .C1(_1045_),
    .X(_1047_));
 sky130_fd_sc_hd__nor2_8 _3464_ (.A(net515),
    .B(net791),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _3465_ (.A1(\gpio_configure[5][4] ),
    .A2(_0941_),
    .B1(_1048_),
    .B2(\gpio_configure[28][12] ),
    .X(_1049_));
 sky130_fd_sc_hd__a221o_4 _3466_ (.A1(\gpio_configure[13][4] ),
    .A2(_0894_),
    .B1(_0954_),
    .B2(\gpio_configure[35][4] ),
    .C1(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__nor2_8 _3467_ (.A(net609),
    .B(net791),
    .Y(_1051_));
 sky130_fd_sc_hd__nor2_8 _3468_ (.A(net360),
    .B(_0921_),
    .Y(_1052_));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(\gpio_configure[20][12] ),
    .A2(_1051_),
    .B1(_1052_),
    .B2(\gpio_configure[25][12] ),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_8 _3470_ (.A(net609),
    .B(_0871_),
    .Y(_1054_));
 sky130_fd_sc_hd__a221o_2 _3471_ (.A1(\gpio_configure[31][4] ),
    .A2(_0944_),
    .B1(_1054_),
    .B2(\gpio_configure[21][12] ),
    .C1(_1053_),
    .X(_1055_));
 sky130_fd_sc_hd__or4_1 _3472_ (.A(_1042_),
    .B(_1047_),
    .C(_1050_),
    .D(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__nor2_8 _3473_ (.A(_0883_),
    .B(_0956_),
    .Y(_1057_));
 sky130_fd_sc_hd__a22o_1 _3474_ (.A1(\gpio_configure[8][4] ),
    .A2(_0913_),
    .B1(_1057_),
    .B2(\gpio_configure[4][12] ),
    .X(_1058_));
 sky130_fd_sc_hd__a221o_4 _3475_ (.A1(\gpio_configure[3][4] ),
    .A2(_0942_),
    .B1(_0961_),
    .B2(\gpio_configure[16][4] ),
    .C1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__nor2_4 _3476_ (.A(_0868_),
    .B(_0971_),
    .Y(_1060_));
 sky130_fd_sc_hd__a211o_4 _3477_ (.A1(net39),
    .A2(_0899_),
    .B1(_0973_),
    .C1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__nor2_8 _3478_ (.A(_0871_),
    .B(net354),
    .Y(_1062_));
 sky130_fd_sc_hd__a221o_1 _3479_ (.A1(\gpio_configure[2][4] ),
    .A2(_0963_),
    .B1(_1062_),
    .B2(\gpio_configure[13][12] ),
    .C1(_1061_),
    .X(_1063_));
 sky130_fd_sc_hd__nor2_8 _3480_ (.A(net355),
    .B(_0932_),
    .Y(_1064_));
 sky130_fd_sc_hd__nor2_8 _3481_ (.A(_0871_),
    .B(net355),
    .Y(_1065_));
 sky130_fd_sc_hd__a22o_1 _3482_ (.A1(\gpio_configure[25][4] ),
    .A2(_0887_),
    .B1(_1065_),
    .B2(\gpio_configure[5][12] ),
    .X(_1066_));
 sky130_fd_sc_hd__a221o_1 _3483_ (.A1(\gpio_configure[29][4] ),
    .A2(_0875_),
    .B1(_1064_),
    .B2(\gpio_configure[8][12] ),
    .C1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__nor2_8 _3484_ (.A(net355),
    .B(_0971_),
    .Y(_1068_));
 sky130_fd_sc_hd__nor2_8 _3485_ (.A(net569),
    .B(_0932_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22o_4 _3486_ (.A1(\gpio_configure[3][12] ),
    .A2(_1068_),
    .B1(_1069_),
    .B2(\gpio_configure[0][12] ),
    .X(_1070_));
 sky130_fd_sc_hd__a221o_4 _3487_ (.A1(\gpio_configure[32][4] ),
    .A2(_0900_),
    .B1(_0964_),
    .B2(\gpio_configure[12][4] ),
    .C1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__or4_2 _3488_ (.A(_1059_),
    .B(_1063_),
    .C(_1067_),
    .D(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_8 _3489_ (.A(net354),
    .B(_0971_),
    .Y(_1073_));
 sky130_fd_sc_hd__a22o_2 _3490_ (.A1(net65),
    .A2(_1006_),
    .B1(_1073_),
    .B2(\gpio_configure[11][12] ),
    .X(_1074_));
 sky130_fd_sc_hd__nor2_8 _3491_ (.A(net515),
    .B(_1005_),
    .Y(_1075_));
 sky130_fd_sc_hd__a221o_4 _3492_ (.A1(\gpio_configure[4][4] ),
    .A2(_0936_),
    .B1(_1075_),
    .B2(\gpio_configure[30][12] ),
    .C1(_1074_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_8 _3493_ (.A(net609),
    .B(_1007_),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_8 _3494_ (.A(net515),
    .B(_1007_),
    .Y(_1078_));
 sky130_fd_sc_hd__a22o_1 _3495_ (.A1(\gpio_configure[18][12] ),
    .A2(_1077_),
    .B1(_1078_),
    .B2(\gpio_configure[26][12] ),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_2 _3496_ (.A1(net24),
    .A2(_0891_),
    .B1(_0951_),
    .B2(\gpio_configure[11][4] ),
    .C1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__nor2_8 _3497_ (.A(net515),
    .B(_0971_),
    .Y(_1081_));
 sky130_fd_sc_hd__a22o_1 _3498_ (.A1(\gpio_configure[17][4] ),
    .A2(_0888_),
    .B1(_1081_),
    .B2(\gpio_configure[27][12] ),
    .X(_1082_));
 sky130_fd_sc_hd__a221o_2 _3499_ (.A1(net7),
    .A2(_0909_),
    .B1(_1008_),
    .B2(net262),
    .C1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__nor2_8 _3500_ (.A(net515),
    .B(_0917_),
    .Y(_1084_));
 sky130_fd_sc_hd__nor2_8 _3501_ (.A(net357),
    .B(_0871_),
    .Y(_1085_));
 sky130_fd_sc_hd__a22o_2 _3502_ (.A1(\gpio_configure[27][4] ),
    .A2(_0865_),
    .B1(_1085_),
    .B2(\gpio_configure[29][12] ),
    .X(_1086_));
 sky130_fd_sc_hd__a221o_1 _3503_ (.A1(\gpio_configure[20][4] ),
    .A2(_0948_),
    .B1(_1084_),
    .B2(\gpio_configure[31][12] ),
    .C1(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__or4_4 _3504_ (.A(_1076_),
    .B(_1080_),
    .C(_1083_),
    .D(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nor2_8 _3505_ (.A(net360),
    .B(_0932_),
    .Y(_1089_));
 sky130_fd_sc_hd__nor2_8 _3506_ (.A(net609),
    .B(_0971_),
    .Y(_1090_));
 sky130_fd_sc_hd__a22o_1 _3507_ (.A1(\gpio_configure[24][12] ),
    .A2(_1089_),
    .B1(_1090_),
    .B2(\gpio_configure[19][12] ),
    .X(_1091_));
 sky130_fd_sc_hd__nor2_8 _3508_ (.A(net515),
    .B(_0921_),
    .Y(_1092_));
 sky130_fd_sc_hd__a221o_4 _3509_ (.A1(serial_bb_clock),
    .A2(_0972_),
    .B1(_1092_),
    .B2(\gpio_configure[33][12] ),
    .C1(_1091_),
    .X(_1093_));
 sky130_fd_sc_hd__nor2_8 _3510_ (.A(net569),
    .B(_0921_),
    .Y(_1094_));
 sky130_fd_sc_hd__nor2_8 _3511_ (.A(net354),
    .B(net791),
    .Y(_1095_));
 sky130_fd_sc_hd__a22o_1 _3512_ (.A1(\gpio_configure[28][4] ),
    .A2(_0953_),
    .B1(_1095_),
    .B2(\gpio_configure[12][12] ),
    .X(_1096_));
 sky130_fd_sc_hd__a221o_1 _3513_ (.A1(net56),
    .A2(_0911_),
    .B1(_1094_),
    .B2(\gpio_configure[1][12] ),
    .C1(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_8 _3514_ (.A(net360),
    .B(_1005_),
    .Y(_1098_));
 sky130_fd_sc_hd__nor2_8 _3515_ (.A(net569),
    .B(net749),
    .Y(_1099_));
 sky130_fd_sc_hd__a22o_2 _3516_ (.A1(\gpio_configure[22][12] ),
    .A2(_1098_),
    .B1(_1099_),
    .B2(net270),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _3517_ (.A1(\gpio_configure[19][4] ),
    .A2(_0863_),
    .B1(_0906_),
    .B2(\gpio_configure[26][4] ),
    .C1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__nor2_8 _3518_ (.A(net355),
    .B(_0921_),
    .Y(_1102_));
 sky130_fd_sc_hd__a22o_2 _3519_ (.A1(\gpio_configure[33][4] ),
    .A2(_0960_),
    .B1(_1102_),
    .B2(\gpio_configure[9][12] ),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_8 _3520_ (.A(net358),
    .B(_0971_),
    .Y(_1104_));
 sky130_fd_sc_hd__a221o_4 _3521_ (.A1(\gpio_configure[10][4] ),
    .A2(_0945_),
    .B1(_1104_),
    .B2(\gpio_configure[35][12] ),
    .C1(_1103_),
    .X(_1105_));
 sky130_fd_sc_hd__or4_1 _3522_ (.A(_1093_),
    .B(_1097_),
    .C(_1101_),
    .D(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _3523_ (.A1(\gpio_configure[0][4] ),
    .A2(_0904_),
    .B1(_0923_),
    .B2(\gpio_configure[23][4] ),
    .X(_1107_));
 sky130_fd_sc_hd__nor2_8 _3524_ (.A(net358),
    .B(_1007_),
    .Y(_1108_));
 sky130_fd_sc_hd__a221o_1 _3525_ (.A1(\gpio_configure[22][4] ),
    .A2(_0928_),
    .B1(_1108_),
    .B2(\gpio_configure[34][12] ),
    .C1(_1107_),
    .X(_1109_));
 sky130_fd_sc_hd__a22o_4 _3526_ (.A1(net287),
    .A2(_0922_),
    .B1(_0933_),
    .B2(net295),
    .X(_1110_));
 sky130_fd_sc_hd__a221o_4 _3527_ (.A1(net48),
    .A2(_0918_),
    .B1(_0935_),
    .B2(\gpio_configure[36][4] ),
    .C1(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__nor2_8 _3528_ (.A(net359),
    .B(net791),
    .Y(_1112_));
 sky130_fd_sc_hd__nor2_8 _3529_ (.A(net355),
    .B(_0917_),
    .Y(_1113_));
 sky130_fd_sc_hd__a22o_1 _3530_ (.A1(\gpio_configure[36][12] ),
    .A2(_1112_),
    .B1(_1113_),
    .B2(\gpio_configure[7][12] ),
    .X(_1114_));
 sky130_fd_sc_hd__nor2_8 _3531_ (.A(net355),
    .B(_1005_),
    .Y(_1115_));
 sky130_fd_sc_hd__a221o_1 _3532_ (.A1(\gpio_configure[30][4] ),
    .A2(_0930_),
    .B1(_1115_),
    .B2(\gpio_configure[6][12] ),
    .C1(_1114_),
    .X(_1116_));
 sky130_fd_sc_hd__or3_1 _3533_ (.A(_1109_),
    .B(_1111_),
    .C(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__nor2_8 _3534_ (.A(_0871_),
    .B(net359),
    .Y(_1118_));
 sky130_fd_sc_hd__a22o_4 _3535_ (.A1(net30),
    .A2(_0872_),
    .B1(_0947_),
    .B2(\gpio_configure[34][4] ),
    .X(_1119_));
 sky130_fd_sc_hd__a221o_1 _3536_ (.A1(\gpio_configure[24][4] ),
    .A2(_0880_),
    .B1(_1118_),
    .B2(\gpio_configure[37][12] ),
    .C1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a22o_1 _3537_ (.A1(\gpio_configure[9][4] ),
    .A2(_0895_),
    .B1(_0958_),
    .B2(\gpio_configure[15][4] ),
    .X(_1121_));
 sky130_fd_sc_hd__a221o_2 _3538_ (.A1(\gpio_configure[1][4] ),
    .A2(_0884_),
    .B1(_0916_),
    .B2(\gpio_configure[14][4] ),
    .C1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_8 _3539_ (.A(net354),
    .B(_1005_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor2_8 _3540_ (.A(net354),
    .B(_0921_),
    .Y(_1124_));
 sky130_fd_sc_hd__a22o_1 _3541_ (.A1(\gpio_configure[14][12] ),
    .A2(_1123_),
    .B1(_1124_),
    .B2(\gpio_configure[17][12] ),
    .X(_1125_));
 sky130_fd_sc_hd__a221o_1 _3542_ (.A1(\gpio_configure[21][4] ),
    .A2(_0890_),
    .B1(_0914_),
    .B2(\gpio_configure[7][4] ),
    .C1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_8 _3543_ (.A(net355),
    .B(_1007_),
    .Y(_1127_));
 sky130_fd_sc_hd__a22o_1 _3544_ (.A1(net278),
    .A2(_0924_),
    .B1(_0939_),
    .B2(\gpio_configure[37][4] ),
    .X(_1128_));
 sky130_fd_sc_hd__a221o_2 _3545_ (.A1(clknet_2_2_0_mgmt_gpio_in[4]),
    .A2(_0950_),
    .B1(_1127_),
    .B2(\gpio_configure[2][12] ),
    .C1(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__or4_2 _3546_ (.A(_1120_),
    .B(_1122_),
    .C(_1126_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__or4_2 _3547_ (.A(_1088_),
    .B(_1106_),
    .C(_1117_),
    .D(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__or3_2 _3548_ (.A(_1056_),
    .B(_1072_),
    .C(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(clknet_1_0__leaf__1132_),
    .A1(\hkspi.ldata[3] ),
    .S(_0837_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(_1133_),
    .A1(\hkspi.ldata[4] ),
    .S(_0969_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_4 _3551_ (.A(_0903_),
    .B(_0910_),
    .Y(_1134_));
 sky130_fd_sc_hd__nor2_8 _3552_ (.A(net546),
    .B(net639),
    .Y(_1135_));
 sky130_fd_sc_hd__a22o_1 _3553_ (.A1(\gpio_configure[31][3] ),
    .A2(_0944_),
    .B1(_1043_),
    .B2(\gpio_configure[32][11] ),
    .X(_1136_));
 sky130_fd_sc_hd__a22o_1 _3554_ (.A1(\gpio_configure[11][3] ),
    .A2(_0951_),
    .B1(_0964_),
    .B2(\gpio_configure[12][3] ),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _3555_ (.A1(net38),
    .A2(_0899_),
    .B1(_1108_),
    .B2(\gpio_configure[34][11] ),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_4 _3556_ (.A1(\gpio_configure[25][3] ),
    .A2(_0887_),
    .B1(_0953_),
    .B2(\gpio_configure[28][3] ),
    .X(_1139_));
 sky130_fd_sc_hd__a22o_1 _3557_ (.A1(\gpio_configure[24][3] ),
    .A2(_0880_),
    .B1(_1089_),
    .B2(\gpio_configure[24][11] ),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _3558_ (.A1(\gpio_configure[29][3] ),
    .A2(_0875_),
    .B1(_1069_),
    .B2(\gpio_configure[0][11] ),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_2 _3559_ (.A1(\gpio_configure[32][3] ),
    .A2(_0900_),
    .B1(_0972_),
    .B2(serial_bb_load),
    .X(_1142_));
 sky130_fd_sc_hd__a22o_2 _3560_ (.A1(\gpio_configure[19][3] ),
    .A2(_0863_),
    .B1(_0957_),
    .B2(net14),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _3561_ (.A1(\gpio_configure[17][3] ),
    .A2(_0888_),
    .B1(_0923_),
    .B2(\gpio_configure[23][3] ),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_4 _3562_ (.A1(\gpio_configure[25][11] ),
    .A2(_1052_),
    .B1(_1090_),
    .B2(\gpio_configure[19][11] ),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _3563_ (.A1(\gpio_configure[0][3] ),
    .A2(_0904_),
    .B1(_1078_),
    .B2(\gpio_configure[26][11] ),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _3564_ (.A1(\gpio_configure[18][3] ),
    .A2(_0938_),
    .B1(_1054_),
    .B2(\gpio_configure[21][11] ),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _3565_ (.A1(\gpio_configure[20][3] ),
    .A2(_0948_),
    .B1(_1077_),
    .B2(\gpio_configure[18][11] ),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _3566_ (.A1(\gpio_configure[10][3] ),
    .A2(_0945_),
    .B1(_1046_),
    .B2(\gpio_configure[15][11] ),
    .X(_1149_));
 sky130_fd_sc_hd__a221o_2 _3567_ (.A1(\gpio_configure[7][3] ),
    .A2(_0914_),
    .B1(_0916_),
    .B2(\gpio_configure[14][3] ),
    .C1(_1137_),
    .X(_1150_));
 sky130_fd_sc_hd__a221o_4 _3568_ (.A1(\gpio_configure[9][11] ),
    .A2(_1102_),
    .B1(_1113_),
    .B2(\gpio_configure[7][11] ),
    .C1(_1138_),
    .X(_1151_));
 sky130_fd_sc_hd__a211o_1 _3569_ (.A1(\gpio_configure[9][3] ),
    .A2(_0895_),
    .B1(_1150_),
    .C1(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a22o_4 _3570_ (.A1(\gpio_configure[35][11] ),
    .A2(_1104_),
    .B1(_1124_),
    .B2(\gpio_configure[17][11] ),
    .X(_1153_));
 sky130_fd_sc_hd__a221o_1 _3571_ (.A1(net46),
    .A2(_0918_),
    .B1(_0954_),
    .B2(\gpio_configure[35][3] ),
    .C1(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__a22o_4 _3572_ (.A1(\gpio_configure[10][11] ),
    .A2(_1039_),
    .B1(_1062_),
    .B2(\gpio_configure[13][11] ),
    .X(_1155_));
 sky130_fd_sc_hd__a221o_1 _3573_ (.A1(\gpio_configure[13][3] ),
    .A2(_0894_),
    .B1(_1135_),
    .B2(net304),
    .C1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _3574_ (.A1(\gpio_configure[37][3] ),
    .A2(_0939_),
    .B1(_0960_),
    .B2(\gpio_configure[33][3] ),
    .X(_1157_));
 sky130_fd_sc_hd__a221o_4 _3575_ (.A1(\gpio_configure[4][3] ),
    .A2(_0936_),
    .B1(_0961_),
    .B2(\gpio_configure[16][3] ),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__a22o_1 _3576_ (.A1(\gpio_configure[3][3] ),
    .A2(_0942_),
    .B1(_1065_),
    .B2(\gpio_configure[5][11] ),
    .X(_1159_));
 sky130_fd_sc_hd__a221o_2 _3577_ (.A1(\gpio_configure[2][3] ),
    .A2(_0963_),
    .B1(_1068_),
    .B2(\gpio_configure[3][11] ),
    .C1(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__or4_1 _3578_ (.A(_1154_),
    .B(_1156_),
    .C(_1158_),
    .D(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__a22o_2 _3579_ (.A1(\gpio_configure[12][11] ),
    .A2(_1095_),
    .B1(_1123_),
    .B2(\gpio_configure[14][11] ),
    .X(_1162_));
 sky130_fd_sc_hd__a221o_2 _3580_ (.A1(\gpio_configure[1][3] ),
    .A2(_0884_),
    .B1(_1127_),
    .B2(\gpio_configure[2][11] ),
    .C1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__a22o_1 _3581_ (.A1(\gpio_configure[6][3] ),
    .A2(_0927_),
    .B1(_1115_),
    .B2(\gpio_configure[6][11] ),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _3582_ (.A1(\gpio_configure[8][3] ),
    .A2(_0913_),
    .B1(_0941_),
    .B2(\gpio_configure[5][3] ),
    .C1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__a22o_1 _3583_ (.A1(\gpio_configure[34][3] ),
    .A2(_0947_),
    .B1(_1112_),
    .B2(\gpio_configure[36][11] ),
    .X(_1166_));
 sky130_fd_sc_hd__a221o_4 _3584_ (.A1(net55),
    .A2(_0911_),
    .B1(_1041_),
    .B2(\gpio_configure[16][11] ),
    .C1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a22o_4 _3585_ (.A1(\gpio_configure[4][11] ),
    .A2(_1057_),
    .B1(_1073_),
    .B2(\gpio_configure[11][11] ),
    .X(_1168_));
 sky130_fd_sc_hd__a221o_4 _3586_ (.A1(\gpio_configure[15][3] ),
    .A2(_0958_),
    .B1(_1006_),
    .B2(net64),
    .C1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__or4_1 _3587_ (.A(_1163_),
    .B(_1165_),
    .C(_1167_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__or4_4 _3588_ (.A(_1149_),
    .B(_1152_),
    .C(_1161_),
    .D(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__a221o_1 _3589_ (.A1(net23),
    .A2(_0891_),
    .B1(_0928_),
    .B2(\gpio_configure[22][3] ),
    .C1(_1136_),
    .X(_1172_));
 sky130_fd_sc_hd__a221o_1 _3590_ (.A1(net261),
    .A2(_1008_),
    .B1(_1134_),
    .B2(net95),
    .C1(_1142_),
    .X(_1173_));
 sky130_fd_sc_hd__a221o_2 _3591_ (.A1(\gpio_configure[28][11] ),
    .A2(_1048_),
    .B1(_1081_),
    .B2(\gpio_configure[27][11] ),
    .C1(_1148_),
    .X(_1174_));
 sky130_fd_sc_hd__a221o_2 _3592_ (.A1(\gpio_configure[30][11] ),
    .A2(_1075_),
    .B1(_1099_),
    .B2(net269),
    .C1(_1139_),
    .X(_1175_));
 sky130_fd_sc_hd__or4_1 _3593_ (.A(_1172_),
    .B(_1173_),
    .C(_1174_),
    .D(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__a221o_1 _3594_ (.A1(net277),
    .A2(_0924_),
    .B1(_1051_),
    .B2(\gpio_configure[20][11] ),
    .C1(_1140_),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_4 _3595_ (.A1(\gpio_configure[26][3] ),
    .A2(_0906_),
    .B1(_1085_),
    .B2(\gpio_configure[29][11] ),
    .C1(_1141_),
    .X(_1178_));
 sky130_fd_sc_hd__a221o_1 _3596_ (.A1(net285),
    .A2(_0922_),
    .B1(_0933_),
    .B2(net294),
    .C1(_1147_),
    .X(_1179_));
 sky130_fd_sc_hd__a221o_2 _3597_ (.A1(net29),
    .A2(_0872_),
    .B1(_0909_),
    .B2(net6),
    .C1(_1145_),
    .X(_1180_));
 sky130_fd_sc_hd__or4_4 _3598_ (.A(_1177_),
    .B(_1178_),
    .C(_1179_),
    .D(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_1 _3599_ (.A1(\gpio_configure[27][3] ),
    .A2(_0865_),
    .B1(_1084_),
    .B2(\gpio_configure[31][11] ),
    .C1(_1146_),
    .X(_1182_));
 sky130_fd_sc_hd__a221o_1 _3600_ (.A1(\gpio_configure[33][11] ),
    .A2(_1092_),
    .B1(_1094_),
    .B2(\gpio_configure[1][11] ),
    .C1(_1143_),
    .X(_1183_));
 sky130_fd_sc_hd__a221o_1 _3601_ (.A1(\gpio_configure[21][3] ),
    .A2(_0890_),
    .B1(_1044_),
    .B2(\gpio_configure[23][11] ),
    .C1(_1144_),
    .X(_1184_));
 sky130_fd_sc_hd__a22o_1 _3602_ (.A1(\gpio_configure[36][3] ),
    .A2(_0935_),
    .B1(_1064_),
    .B2(\gpio_configure[8][11] ),
    .X(_1185_));
 sky130_fd_sc_hd__a221o_4 _3603_ (.A1(net67),
    .A2(_0950_),
    .B1(_1118_),
    .B2(\gpio_configure[37][11] ),
    .C1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__a221o_1 _3604_ (.A1(\gpio_configure[30][3] ),
    .A2(_0930_),
    .B1(_1098_),
    .B2(\gpio_configure[22][11] ),
    .C1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__or4_1 _3605_ (.A(_1182_),
    .B(_1183_),
    .C(_1184_),
    .D(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__or4_4 _3606_ (.A(_1171_),
    .B(_1176_),
    .C(_1181_),
    .D(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _3607_ (.A0(_1189_),
    .A1(\hkspi.ldata[2] ),
    .S(_0837_),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(_1190_),
    .A1(\hkspi.ldata[3] ),
    .S(_0969_),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_8 _3609_ (.A(net569),
    .B(_0917_),
    .Y(_1191_));
 sky130_fd_sc_hd__a22o_1 _3610_ (.A1(net63),
    .A2(_1006_),
    .B1(_1102_),
    .B2(\gpio_configure[9][10] ),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _3611_ (.A1(net37),
    .A2(_0899_),
    .B1(_1064_),
    .B2(\gpio_configure[8][10] ),
    .X(_1193_));
 sky130_fd_sc_hd__a22o_1 _3612_ (.A1(\gpio_configure[4][10] ),
    .A2(_1057_),
    .B1(_1127_),
    .B2(\gpio_configure[2][10] ),
    .X(_1194_));
 sky130_fd_sc_hd__a22o_4 _3613_ (.A1(net58),
    .A2(_0950_),
    .B1(_0960_),
    .B2(\gpio_configure[33][2] ),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_2 _3614_ (.A1(\gpio_configure[37][2] ),
    .A2(_0939_),
    .B1(_1135_),
    .B2(net303),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _3615_ (.A1(\gpio_configure[10][2] ),
    .A2(_0945_),
    .B1(_1095_),
    .B2(\gpio_configure[12][10] ),
    .X(_1197_));
 sky130_fd_sc_hd__a22o_1 _3616_ (.A1(\gpio_configure[13][2] ),
    .A2(_0894_),
    .B1(_0958_),
    .B2(\gpio_configure[15][2] ),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _3617_ (.A1(\gpio_configure[4][2] ),
    .A2(_0936_),
    .B1(_0942_),
    .B2(\gpio_configure[3][2] ),
    .X(_1199_));
 sky130_fd_sc_hd__a22o_1 _3618_ (.A1(\gpio_configure[10][10] ),
    .A2(_1039_),
    .B1(_1065_),
    .B2(\gpio_configure[5][10] ),
    .X(_1200_));
 sky130_fd_sc_hd__a22o_2 _3619_ (.A1(\gpio_configure[14][2] ),
    .A2(_0916_),
    .B1(_0951_),
    .B2(\gpio_configure[11][2] ),
    .X(_1201_));
 sky130_fd_sc_hd__a22o_1 _3620_ (.A1(\gpio_configure[36][2] ),
    .A2(_0935_),
    .B1(_1104_),
    .B2(\gpio_configure[35][10] ),
    .X(_1202_));
 sky130_fd_sc_hd__a221o_4 _3621_ (.A1(\gpio_configure[7][2] ),
    .A2(_0914_),
    .B1(_0918_),
    .B2(net45),
    .C1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__a221o_1 _3622_ (.A1(\gpio_configure[7][10] ),
    .A2(_1113_),
    .B1(_1123_),
    .B2(\gpio_configure[14][10] ),
    .C1(_1196_),
    .X(_1204_));
 sky130_fd_sc_hd__a221o_1 _3623_ (.A1(\gpio_configure[13][10] ),
    .A2(_1062_),
    .B1(_1124_),
    .B2(\gpio_configure[17][10] ),
    .C1(_1201_),
    .X(_1205_));
 sky130_fd_sc_hd__a2111o_2 _3624_ (.A1(\gpio_configure[36][10] ),
    .A2(_1112_),
    .B1(_1195_),
    .C1(_1204_),
    .D1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a221o_1 _3625_ (.A1(\gpio_configure[12][2] ),
    .A2(_0964_),
    .B1(_1118_),
    .B2(\gpio_configure[37][10] ),
    .C1(_1192_),
    .X(_1207_));
 sky130_fd_sc_hd__a221o_1 _3626_ (.A1(\gpio_configure[8][2] ),
    .A2(_0913_),
    .B1(_1068_),
    .B2(\gpio_configure[3][10] ),
    .C1(_1197_),
    .X(_1208_));
 sky130_fd_sc_hd__a221o_1 _3627_ (.A1(\gpio_configure[16][2] ),
    .A2(_0961_),
    .B1(_1046_),
    .B2(\gpio_configure[15][10] ),
    .C1(_1198_),
    .X(_1209_));
 sky130_fd_sc_hd__a221o_1 _3628_ (.A1(net54),
    .A2(_0911_),
    .B1(_1108_),
    .B2(\gpio_configure[34][10] ),
    .C1(_1199_),
    .X(_1210_));
 sky130_fd_sc_hd__or4_1 _3629_ (.A(_1207_),
    .B(_1208_),
    .C(_1209_),
    .D(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _3630_ (.A1(\gpio_configure[9][2] ),
    .A2(_0895_),
    .B1(_1073_),
    .B2(\gpio_configure[11][10] ),
    .C1(_1200_),
    .X(_1212_));
 sky130_fd_sc_hd__a221o_1 _3631_ (.A1(\gpio_configure[6][2] ),
    .A2(_0927_),
    .B1(_0963_),
    .B2(\gpio_configure[2][2] ),
    .C1(_1193_),
    .X(_1213_));
 sky130_fd_sc_hd__a221o_1 _3632_ (.A1(\gpio_configure[16][10] ),
    .A2(_1041_),
    .B1(_1115_),
    .B2(\gpio_configure[6][10] ),
    .C1(_1194_),
    .X(_1214_));
 sky130_fd_sc_hd__a22o_1 _3633_ (.A1(\gpio_configure[34][2] ),
    .A2(_0947_),
    .B1(_0954_),
    .B2(\gpio_configure[35][2] ),
    .X(_1215_));
 sky130_fd_sc_hd__a221o_1 _3634_ (.A1(\gpio_configure[1][2] ),
    .A2(_0884_),
    .B1(_0941_),
    .B2(\gpio_configure[5][2] ),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__or4_1 _3635_ (.A(_1212_),
    .B(_1213_),
    .C(_1214_),
    .D(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__or4_4 _3636_ (.A(_1203_),
    .B(_1206_),
    .C(_1211_),
    .D(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__a22o_1 _3637_ (.A1(\gpio_configure[27][2] ),
    .A2(_0865_),
    .B1(_1085_),
    .B2(\gpio_configure[29][10] ),
    .X(_1219_));
 sky130_fd_sc_hd__a221o_2 _3638_ (.A1(\gpio_configure[22][2] ),
    .A2(_0928_),
    .B1(_0953_),
    .B2(\gpio_configure[28][2] ),
    .C1(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__a22o_1 _3639_ (.A1(net22),
    .A2(_0891_),
    .B1(_1090_),
    .B2(\gpio_configure[19][10] ),
    .X(_1221_));
 sky130_fd_sc_hd__a221o_4 _3640_ (.A1(net5),
    .A2(_0909_),
    .B1(_0933_),
    .B2(net293),
    .C1(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__a22o_1 _3641_ (.A1(\gpio_configure[32][10] ),
    .A2(_1043_),
    .B1(_1092_),
    .B2(\gpio_configure[33][10] ),
    .X(_1223_));
 sky130_fd_sc_hd__a221o_1 _3642_ (.A1(\gpio_configure[25][2] ),
    .A2(_0887_),
    .B1(_0972_),
    .B2(serial_bb_resetn),
    .C1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a22o_1 _3643_ (.A1(net26),
    .A2(_0872_),
    .B1(_1048_),
    .B2(\gpio_configure[28][10] ),
    .X(_1225_));
 sky130_fd_sc_hd__a221o_1 _3644_ (.A1(\gpio_configure[21][2] ),
    .A2(_0890_),
    .B1(_1077_),
    .B2(\gpio_configure[18][10] ),
    .C1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__or4_1 _3645_ (.A(_1220_),
    .B(_1222_),
    .C(_1224_),
    .D(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_1 _3646_ (.A1(\gpio_configure[27][10] ),
    .A2(_1081_),
    .B1(_1099_),
    .B2(net268),
    .X(_1228_));
 sky130_fd_sc_hd__a221o_2 _3647_ (.A1(net274),
    .A2(_1008_),
    .B1(_1075_),
    .B2(\gpio_configure[30][10] ),
    .C1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__a22o_1 _3648_ (.A1(\gpio_configure[23][2] ),
    .A2(_0923_),
    .B1(_1078_),
    .B2(\gpio_configure[26][10] ),
    .X(_1230_));
 sky130_fd_sc_hd__a221o_1 _3649_ (.A1(\gpio_configure[24][2] ),
    .A2(_0880_),
    .B1(_0922_),
    .B2(net284),
    .C1(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__a22o_4 _3650_ (.A1(net13),
    .A2(_0957_),
    .B1(_1191_),
    .B2(clk1_output_dest),
    .X(_1232_));
 sky130_fd_sc_hd__a221o_4 _3651_ (.A1(\gpio_configure[0][10] ),
    .A2(_1069_),
    .B1(_1084_),
    .B2(\gpio_configure[31][10] ),
    .C1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__a22o_2 _3652_ (.A1(\gpio_configure[31][2] ),
    .A2(_0944_),
    .B1(_1134_),
    .B2(net97),
    .X(_1234_));
 sky130_fd_sc_hd__a221o_1 _3653_ (.A1(\gpio_configure[29][2] ),
    .A2(_0875_),
    .B1(_0924_),
    .B2(net276),
    .C1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__or4_1 _3654_ (.A(_1229_),
    .B(_1231_),
    .C(_1233_),
    .D(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__a22o_1 _3655_ (.A1(\gpio_configure[17][2] ),
    .A2(_0888_),
    .B1(_1054_),
    .B2(\gpio_configure[21][10] ),
    .X(_1237_));
 sky130_fd_sc_hd__a221o_1 _3656_ (.A1(\gpio_configure[19][2] ),
    .A2(_0863_),
    .B1(_0948_),
    .B2(\gpio_configure[20][2] ),
    .C1(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__a22o_1 _3657_ (.A1(\gpio_configure[26][2] ),
    .A2(_0906_),
    .B1(_0930_),
    .B2(\gpio_configure[30][2] ),
    .X(_1239_));
 sky130_fd_sc_hd__a221o_4 _3658_ (.A1(\gpio_configure[32][2] ),
    .A2(_0900_),
    .B1(_0904_),
    .B2(\gpio_configure[0][2] ),
    .C1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_1 _3659_ (.A1(\gpio_configure[23][10] ),
    .A2(_1044_),
    .B1(_1089_),
    .B2(\gpio_configure[24][10] ),
    .X(_1241_));
 sky130_fd_sc_hd__a221o_1 _3660_ (.A1(\gpio_configure[20][10] ),
    .A2(_1051_),
    .B1(_1052_),
    .B2(\gpio_configure[25][10] ),
    .C1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__a2bb2o_1 _3661_ (.A1_N(_0868_),
    .A2_N(_1007_),
    .B1(_1094_),
    .B2(\gpio_configure[1][10] ),
    .X(_1243_));
 sky130_fd_sc_hd__a22o_1 _3662_ (.A1(\gpio_configure[18][2] ),
    .A2(_0938_),
    .B1(_1098_),
    .B2(\gpio_configure[22][10] ),
    .X(_1244_));
 sky130_fd_sc_hd__or4_1 _3663_ (.A(_0973_),
    .B(_1242_),
    .C(_1243_),
    .D(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__or4_1 _3664_ (.A(_1236_),
    .B(_1238_),
    .C(_1240_),
    .D(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__or3_4 _3665_ (.A(_1218_),
    .B(_1227_),
    .C(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(_1247_),
    .A1(\hkspi.ldata[1] ),
    .S(_0837_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(_1248_),
    .A1(\hkspi.ldata[2] ),
    .S(_0969_),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_2 _3668_ (.A(net578),
    .B(net569),
    .Y(_1249_));
 sky130_fd_sc_hd__a22o_2 _3669_ (.A1(\gpio_configure[18][9] ),
    .A2(_1077_),
    .B1(_1249_),
    .B2(net292),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_1 _3670_ (.A1(\gpio_configure[1][1] ),
    .A2(_0884_),
    .B1(_0916_),
    .B2(\gpio_configure[14][1] ),
    .X(_1251_));
 sky130_fd_sc_hd__a22o_4 _3671_ (.A1(\gpio_configure[19][9] ),
    .A2(_1090_),
    .B1(_1099_),
    .B2(net267),
    .X(_1252_));
 sky130_fd_sc_hd__nor2_8 _3672_ (.A(net482),
    .B(net569),
    .Y(_1253_));
 sky130_fd_sc_hd__nor2_4 _3673_ (.A(net356),
    .B(_0874_),
    .Y(_1254_));
 sky130_fd_sc_hd__a22o_4 _3674_ (.A1(\gpio_configure[37][1] ),
    .A2(_0939_),
    .B1(_1006_),
    .B2(net62),
    .X(_1255_));
 sky130_fd_sc_hd__a22o_1 _3675_ (.A1(\gpio_configure[34][1] ),
    .A2(_0947_),
    .B1(_0950_),
    .B2(net47),
    .X(_1256_));
 sky130_fd_sc_hd__a22o_1 _3676_ (.A1(net35),
    .A2(_0909_),
    .B1(_1094_),
    .B2(\gpio_configure[1][9] ),
    .X(_1257_));
 sky130_fd_sc_hd__a221o_1 _3677_ (.A1(net300),
    .A2(_0924_),
    .B1(_1098_),
    .B2(\gpio_configure[22][9] ),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__a22o_1 _3678_ (.A1(serial_bb_enable),
    .A2(_0972_),
    .B1(_1051_),
    .B2(\gpio_configure[20][9] ),
    .X(_1259_));
 sky130_fd_sc_hd__a22o_1 _3679_ (.A1(\gpio_configure[33][1] ),
    .A2(_0960_),
    .B1(_1112_),
    .B2(\gpio_configure[36][9] ),
    .X(_1260_));
 sky130_fd_sc_hd__a22o_4 _3680_ (.A1(\gpio_configure[13][1] ),
    .A2(_0894_),
    .B1(_0961_),
    .B2(\gpio_configure[16][1] ),
    .X(_1261_));
 sky130_fd_sc_hd__a22o_1 _3681_ (.A1(\gpio_configure[23][1] ),
    .A2(_0923_),
    .B1(_1191_),
    .B2(clk2_output_dest),
    .X(_1262_));
 sky130_fd_sc_hd__a221o_1 _3682_ (.A1(net15),
    .A2(_0872_),
    .B1(_1104_),
    .B2(\gpio_configure[35][9] ),
    .C1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__a22o_1 _3683_ (.A1(\gpio_configure[0][1] ),
    .A2(_0904_),
    .B1(_0945_),
    .B2(\gpio_configure[10][1] ),
    .X(_1264_));
 sky130_fd_sc_hd__a221o_1 _3684_ (.A1(\gpio_configure[29][1] ),
    .A2(_0875_),
    .B1(_0953_),
    .B2(\gpio_configure[28][1] ),
    .C1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__a22o_1 _3685_ (.A1(\gpio_configure[8][1] ),
    .A2(_0913_),
    .B1(_1113_),
    .B2(\gpio_configure[7][9] ),
    .X(_1266_));
 sky130_fd_sc_hd__a221o_4 _3686_ (.A1(\gpio_configure[5][9] ),
    .A2(_1065_),
    .B1(_1095_),
    .B2(\gpio_configure[12][9] ),
    .C1(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__or3_1 _3687_ (.A(_1263_),
    .B(_1265_),
    .C(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _3688_ (.A1(\gpio_configure[11][1] ),
    .A2(_0951_),
    .B1(_1124_),
    .B2(\gpio_configure[17][9] ),
    .C1(_1251_),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_4 _3689_ (.A1(\gpio_configure[16][9] ),
    .A2(_1041_),
    .B1(_1123_),
    .B2(\gpio_configure[14][9] ),
    .X(_1270_));
 sky130_fd_sc_hd__a221o_4 _3690_ (.A1(\gpio_configure[7][1] ),
    .A2(_0914_),
    .B1(_0936_),
    .B2(\gpio_configure[4][1] ),
    .C1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a221o_1 _3691_ (.A1(\gpio_configure[26][1] ),
    .A2(_0906_),
    .B1(_1039_),
    .B2(\gpio_configure[10][9] ),
    .C1(_1252_),
    .X(_1272_));
 sky130_fd_sc_hd__a221o_1 _3692_ (.A1(\gpio_configure[24][9] ),
    .A2(_1089_),
    .B1(_1134_),
    .B2(net96),
    .C1(_1250_),
    .X(_1273_));
 sky130_fd_sc_hd__or4_2 _3693_ (.A(_1269_),
    .B(_1271_),
    .C(_1272_),
    .D(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _3694_ (.A1(net283),
    .A2(_0922_),
    .B1(_0954_),
    .B2(\gpio_configure[35][1] ),
    .C1(_1259_),
    .X(_1275_));
 sky130_fd_sc_hd__a22o_2 _3695_ (.A1(\gpio_configure[27][1] ),
    .A2(_0865_),
    .B1(_1108_),
    .B2(\gpio_configure[34][9] ),
    .X(_1276_));
 sky130_fd_sc_hd__a221o_1 _3696_ (.A1(net21),
    .A2(_0891_),
    .B1(_0948_),
    .B2(\gpio_configure[20][1] ),
    .C1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__a221o_2 _3697_ (.A1(\gpio_configure[28][9] ),
    .A2(_1048_),
    .B1(_1081_),
    .B2(\gpio_configure[27][9] ),
    .C1(_1255_),
    .X(_1278_));
 sky130_fd_sc_hd__a221o_1 _3698_ (.A1(\gpio_configure[30][1] ),
    .A2(_0930_),
    .B1(_1092_),
    .B2(\gpio_configure[33][9] ),
    .C1(_1256_),
    .X(_1279_));
 sky130_fd_sc_hd__or4_2 _3699_ (.A(_1275_),
    .B(_1277_),
    .C(_1278_),
    .D(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__a22o_1 _3700_ (.A1(\gpio_configure[4][9] ),
    .A2(_1057_),
    .B1(_1078_),
    .B2(\gpio_configure[26][9] ),
    .X(_1281_));
 sky130_fd_sc_hd__a221o_1 _3701_ (.A1(\gpio_configure[24][1] ),
    .A2(_0880_),
    .B1(_1069_),
    .B2(\gpio_configure[0][9] ),
    .C1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__a22o_1 _3702_ (.A1(\gpio_configure[6][1] ),
    .A2(_0927_),
    .B1(_1068_),
    .B2(\gpio_configure[3][9] ),
    .X(_1283_));
 sky130_fd_sc_hd__a221o_2 _3703_ (.A1(\gpio_configure[9][1] ),
    .A2(_0895_),
    .B1(_0958_),
    .B2(\gpio_configure[15][1] ),
    .C1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a22o_1 _3704_ (.A1(\gpio_configure[3][1] ),
    .A2(_0942_),
    .B1(_1062_),
    .B2(\gpio_configure[13][9] ),
    .X(_1285_));
 sky130_fd_sc_hd__a221o_1 _3705_ (.A1(\gpio_configure[5][1] ),
    .A2(_0941_),
    .B1(_1073_),
    .B2(\gpio_configure[11][9] ),
    .C1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a22o_1 _3706_ (.A1(\gpio_configure[2][1] ),
    .A2(_0963_),
    .B1(_1102_),
    .B2(\gpio_configure[9][9] ),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _3707_ (.A1(\gpio_configure[12][1] ),
    .A2(_0964_),
    .B1(_1075_),
    .B2(\gpio_configure[30][9] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a221o_2 _3708_ (.A1(\gpio_configure[25][9] ),
    .A2(_1052_),
    .B1(_1127_),
    .B2(\gpio_configure[2][9] ),
    .C1(_1261_),
    .X(_1289_));
 sky130_fd_sc_hd__or4_4 _3709_ (.A(_1284_),
    .B(_1286_),
    .C(_1288_),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a211o_1 _3710_ (.A1(\gpio_configure[31][9] ),
    .A2(_1084_),
    .B1(_1282_),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a22o_4 _3711_ (.A1(net53),
    .A2(_0911_),
    .B1(_0918_),
    .B2(net44),
    .X(_1292_));
 sky130_fd_sc_hd__a221o_1 _3712_ (.A1(\gpio_configure[32][1] ),
    .A2(_0900_),
    .B1(_1008_),
    .B2(net273),
    .C1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_4 _3713_ (.A1(\gpio_configure[21][9] ),
    .A2(_1054_),
    .B1(_1254_),
    .B2(net265),
    .X(_1294_));
 sky130_fd_sc_hd__a221o_1 _3714_ (.A1(\gpio_configure[36][1] ),
    .A2(_0935_),
    .B1(_1043_),
    .B2(\gpio_configure[32][9] ),
    .C1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__a22o_1 _3715_ (.A1(\gpio_configure[25][1] ),
    .A2(_0887_),
    .B1(_1135_),
    .B2(net302),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _3716_ (.A1(\gpio_configure[19][1] ),
    .A2(_0863_),
    .B1(_0890_),
    .B2(\gpio_configure[21][1] ),
    .C1(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__or4_1 _3717_ (.A(_1258_),
    .B(_1293_),
    .C(_1295_),
    .D(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__a22o_1 _3718_ (.A1(\gpio_configure[31][1] ),
    .A2(_0944_),
    .B1(_1044_),
    .B2(\gpio_configure[23][9] ),
    .X(_1299_));
 sky130_fd_sc_hd__a221o_1 _3719_ (.A1(net72),
    .A2(_0899_),
    .B1(_1085_),
    .B2(\gpio_configure[29][9] ),
    .C1(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__a221o_1 _3720_ (.A1(\gpio_configure[17][1] ),
    .A2(_0888_),
    .B1(_0957_),
    .B2(net12),
    .C1(_1260_),
    .X(_1301_));
 sky130_fd_sc_hd__a22o_1 _3721_ (.A1(net286),
    .A2(_0933_),
    .B1(_1118_),
    .B2(\gpio_configure[37][9] ),
    .X(_1302_));
 sky130_fd_sc_hd__a221o_1 _3722_ (.A1(\gpio_configure[22][1] ),
    .A2(_0928_),
    .B1(_0938_),
    .B2(\gpio_configure[18][1] ),
    .C1(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__a22o_1 _3723_ (.A1(\gpio_configure[6][9] ),
    .A2(_1115_),
    .B1(_1253_),
    .B2(irq_2_inputsrc),
    .X(_1304_));
 sky130_fd_sc_hd__a221o_4 _3724_ (.A1(\gpio_configure[15][9] ),
    .A2(_1046_),
    .B1(_1064_),
    .B2(\gpio_configure[8][9] ),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__or4_1 _3725_ (.A(_1300_),
    .B(_1301_),
    .C(_1303_),
    .D(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__or4_1 _3726_ (.A(_0973_),
    .B(_1291_),
    .C(_1298_),
    .D(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__or4_4 _3727_ (.A(_1268_),
    .B(_1274_),
    .C(_1280_),
    .D(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(_1308_),
    .A1(\hkspi.ldata[0] ),
    .S(_0837_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _3729_ (.A0(_1309_),
    .A1(\hkspi.ldata[1] ),
    .S(_0969_),
    .X(_0380_));
 sky130_fd_sc_hd__or3_4 _3730_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .C(reset_reg),
    .X(net305));
 sky130_fd_sc_hd__nor2_4 _3731_ (.A(net356),
    .B(_0917_),
    .Y(_1310_));
 sky130_fd_sc_hd__nor2_2 _3732_ (.A(net356),
    .B(_1005_),
    .Y(_1311_));
 sky130_fd_sc_hd__nor2_1 _3733_ (.A(net358),
    .B(_0921_),
    .Y(_1312_));
 sky130_fd_sc_hd__a22o_4 _3734_ (.A1(net71),
    .A2(_0899_),
    .B1(_0950_),
    .B2(net36),
    .X(_1313_));
 sky130_fd_sc_hd__nor2_1 _3735_ (.A(net356),
    .B(net587),
    .Y(_1314_));
 sky130_fd_sc_hd__a22o_2 _3736_ (.A1(net43),
    .A2(_0918_),
    .B1(_1135_),
    .B2(net301),
    .X(_1315_));
 sky130_fd_sc_hd__a22o_1 _3737_ (.A1(\gpio_configure[3][0] ),
    .A2(_0942_),
    .B1(_1127_),
    .B2(\gpio_configure[2][8] ),
    .X(_1316_));
 sky130_fd_sc_hd__a22o_2 _3738_ (.A1(\gpio_configure[5][8] ),
    .A2(_1065_),
    .B1(_1102_),
    .B2(\gpio_configure[9][8] ),
    .X(_1317_));
 sky130_fd_sc_hd__a22o_2 _3739_ (.A1(\gpio_configure[9][0] ),
    .A2(_0895_),
    .B1(_0961_),
    .B2(\gpio_configure[16][0] ),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _3740_ (.A1(\gpio_configure[10][0] ),
    .A2(_0945_),
    .B1(_0963_),
    .B2(\gpio_configure[2][0] ),
    .X(_1319_));
 sky130_fd_sc_hd__a22o_1 _3741_ (.A1(\gpio_configure[6][0] ),
    .A2(_0927_),
    .B1(_0935_),
    .B2(\gpio_configure[36][0] ),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_4 _3742_ (.A1(net52),
    .A2(_0911_),
    .B1(_0939_),
    .B2(\gpio_configure[37][0] ),
    .X(_1321_));
 sky130_fd_sc_hd__a22o_1 _3743_ (.A1(\gpio_configure[23][0] ),
    .A2(_0923_),
    .B1(_1311_),
    .B2(net264),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_1 _3744_ (.A1(net299),
    .A2(_0924_),
    .B1(net305),
    .B2(_1310_),
    .X(_1323_));
 sky130_fd_sc_hd__a22o_2 _3745_ (.A1(\gpio_configure[29][0] ),
    .A2(_0875_),
    .B1(_0928_),
    .B2(\gpio_configure[22][0] ),
    .X(_1324_));
 sky130_fd_sc_hd__a22o_1 _3746_ (.A1(\gpio_configure[11][0] ),
    .A2(_0951_),
    .B1(_1124_),
    .B2(\gpio_configure[17][8] ),
    .X(_1325_));
 sky130_fd_sc_hd__a221o_2 _3747_ (.A1(\gpio_configure[1][0] ),
    .A2(_0884_),
    .B1(_0941_),
    .B2(\gpio_configure[5][0] ),
    .C1(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__a22o_1 _3748_ (.A1(\gpio_configure[11][8] ),
    .A2(_1073_),
    .B1(_1095_),
    .B2(\gpio_configure[12][8] ),
    .X(_1327_));
 sky130_fd_sc_hd__a221o_1 _3749_ (.A1(\gpio_configure[14][0] ),
    .A2(_0916_),
    .B1(_1041_),
    .B2(\gpio_configure[16][8] ),
    .C1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a22o_1 _3750_ (.A1(\gpio_configure[13][8] ),
    .A2(_1062_),
    .B1(_1123_),
    .B2(\gpio_configure[14][8] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _3751_ (.A1(\gpio_configure[12][0] ),
    .A2(_0964_),
    .B1(_1057_),
    .B2(\gpio_configure[4][8] ),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a22o_1 _3752_ (.A1(\gpio_configure[34][0] ),
    .A2(_0947_),
    .B1(_1115_),
    .B2(\gpio_configure[6][8] ),
    .X(_1331_));
 sky130_fd_sc_hd__a221o_1 _3753_ (.A1(\gpio_configure[15][0] ),
    .A2(_0958_),
    .B1(_1039_),
    .B2(\gpio_configure[10][8] ),
    .C1(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__or4_2 _3754_ (.A(_1326_),
    .B(_1328_),
    .C(_1330_),
    .D(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a221o_1 _3755_ (.A1(\gpio_configure[8][8] ),
    .A2(_1064_),
    .B1(_1118_),
    .B2(\gpio_configure[37][8] ),
    .C1(_1313_),
    .X(_1334_));
 sky130_fd_sc_hd__a21o_1 _3756_ (.A1(\gpio_configure[7][8] ),
    .A2(_1113_),
    .B1(_1318_),
    .X(_1335_));
 sky130_fd_sc_hd__a221o_1 _3757_ (.A1(\gpio_configure[35][8] ),
    .A2(_1104_),
    .B1(_1312_),
    .B2(hkspi_disable),
    .C1(_1321_),
    .X(_1336_));
 sky130_fd_sc_hd__a221o_2 _3758_ (.A1(\gpio_configure[13][0] ),
    .A2(_0894_),
    .B1(_1046_),
    .B2(\gpio_configure[15][8] ),
    .C1(_1319_),
    .X(_1337_));
 sky130_fd_sc_hd__or4_1 _3759_ (.A(_1334_),
    .B(_1335_),
    .C(_1336_),
    .D(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__a221o_4 _3760_ (.A1(\gpio_configure[33][0] ),
    .A2(_0960_),
    .B1(_1006_),
    .B2(net61),
    .C1(_1320_),
    .X(_1339_));
 sky130_fd_sc_hd__a221o_1 _3761_ (.A1(\gpio_configure[7][0] ),
    .A2(_0914_),
    .B1(_1112_),
    .B2(\gpio_configure[36][8] ),
    .C1(_1315_),
    .X(_1340_));
 sky130_fd_sc_hd__a221o_1 _3762_ (.A1(\gpio_configure[8][0] ),
    .A2(_0913_),
    .B1(_1108_),
    .B2(\gpio_configure[34][8] ),
    .C1(_1316_),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_1 _3763_ (.A1(\gpio_configure[4][0] ),
    .A2(_0936_),
    .B1(_0954_),
    .B2(\gpio_configure[35][0] ),
    .C1(_1317_),
    .X(_1342_));
 sky130_fd_sc_hd__or4_4 _3764_ (.A(_1339_),
    .B(_1340_),
    .C(_1341_),
    .D(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__a22o_1 _3765_ (.A1(net4),
    .A2(_0872_),
    .B1(_0948_),
    .B2(\gpio_configure[20][0] ),
    .X(_1344_));
 sky130_fd_sc_hd__a22o_1 _3766_ (.A1(\gpio_configure[19][0] ),
    .A2(_0863_),
    .B1(_1098_),
    .B2(\gpio_configure[22][8] ),
    .X(_1345_));
 sky130_fd_sc_hd__a211o_2 _3767_ (.A1(net291),
    .A2(_1249_),
    .B1(_1344_),
    .C1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a221o_4 _3768_ (.A1(\gpio_configure[20][8] ),
    .A2(_1051_),
    .B1(_1253_),
    .B2(irq_1_inputsrc),
    .C1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a2111o_1 _3769_ (.A1(\gpio_configure[3][8] ),
    .A2(_1068_),
    .B1(_1343_),
    .C1(_1347_),
    .D1(_1060_),
    .X(_1348_));
 sky130_fd_sc_hd__a221o_4 _3770_ (.A1(\gpio_configure[32][0] ),
    .A2(_0900_),
    .B1(_1075_),
    .B2(\gpio_configure[30][8] ),
    .C1(_1324_),
    .X(_1349_));
 sky130_fd_sc_hd__a22o_1 _3771_ (.A1(\gpio_configure[32][8] ),
    .A2(_1043_),
    .B1(_1078_),
    .B2(\gpio_configure[26][8] ),
    .X(_1350_));
 sky130_fd_sc_hd__a22o_1 _3772_ (.A1(\gpio_configure[23][8] ),
    .A2(_1044_),
    .B1(_1089_),
    .B2(\gpio_configure[24][8] ),
    .X(_1351_));
 sky130_fd_sc_hd__a221o_1 _3773_ (.A1(\gpio_configure[24][0] ),
    .A2(_0880_),
    .B1(_0933_),
    .B2(net275),
    .C1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__a22o_1 _3774_ (.A1(\gpio_configure[1][8] ),
    .A2(_1094_),
    .B1(_1134_),
    .B2(net98),
    .X(_1353_));
 sky130_fd_sc_hd__a221o_4 _3775_ (.A1(\gpio_configure[27][0] ),
    .A2(_0865_),
    .B1(_1048_),
    .B2(\gpio_configure[28][8] ),
    .C1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a2111o_1 _3776_ (.A1(net266),
    .A2(_1099_),
    .B1(_1350_),
    .C1(_1352_),
    .D1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__a22o_2 _3777_ (.A1(\gpio_configure[28][0] ),
    .A2(_0953_),
    .B1(_1085_),
    .B2(\gpio_configure[29][8] ),
    .X(_1356_));
 sky130_fd_sc_hd__a221o_1 _3778_ (.A1(\gpio_configure[0][8] ),
    .A2(_1069_),
    .B1(_1092_),
    .B2(\gpio_configure[33][8] ),
    .C1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__a22o_1 _3779_ (.A1(serial_busy),
    .A2(_0972_),
    .B1(_1081_),
    .B2(\gpio_configure[27][8] ),
    .X(_1358_));
 sky130_fd_sc_hd__a221o_1 _3780_ (.A1(net272),
    .A2(_1008_),
    .B1(_1084_),
    .B2(\gpio_configure[31][8] ),
    .C1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__a22o_2 _3781_ (.A1(net20),
    .A2(_0891_),
    .B1(_0909_),
    .B2(net34),
    .X(_1360_));
 sky130_fd_sc_hd__a221o_2 _3782_ (.A1(\gpio_configure[26][0] ),
    .A2(_0906_),
    .B1(_0944_),
    .B2(\gpio_configure[31][0] ),
    .C1(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__a22o_2 _3783_ (.A1(\gpio_configure[17][0] ),
    .A2(_0888_),
    .B1(_0930_),
    .B2(\gpio_configure[30][0] ),
    .X(_1362_));
 sky130_fd_sc_hd__a221o_1 _3784_ (.A1(net11),
    .A2(_0957_),
    .B1(_1090_),
    .B2(\gpio_configure[19][8] ),
    .C1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__or4_1 _3785_ (.A(_1357_),
    .B(_1359_),
    .C(_1361_),
    .D(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_2 _3786_ (.A1(net282),
    .A2(_0922_),
    .B1(_1254_),
    .B2(net271),
    .C1(_1323_),
    .X(_1365_));
 sky130_fd_sc_hd__a22o_2 _3787_ (.A1(\gpio_configure[0][0] ),
    .A2(_0904_),
    .B1(_1191_),
    .B2(trap_output_dest),
    .X(_1366_));
 sky130_fd_sc_hd__a221o_4 _3788_ (.A1(\gpio_configure[25][0] ),
    .A2(_0887_),
    .B1(_1052_),
    .B2(\gpio_configure[25][8] ),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a32o_1 _3789_ (.A1(net93),
    .A2(_0869_),
    .A3(_0897_),
    .B1(_1077_),
    .B2(\gpio_configure[18][8] ),
    .X(_1368_));
 sky130_fd_sc_hd__a221o_1 _3790_ (.A1(\gpio_configure[18][0] ),
    .A2(_0938_),
    .B1(_1054_),
    .B2(\gpio_configure[21][8] ),
    .C1(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a221o_2 _3791_ (.A1(\gpio_configure[21][0] ),
    .A2(_0890_),
    .B1(_1314_),
    .B2(net172),
    .C1(_1322_),
    .X(_1370_));
 sky130_fd_sc_hd__or4_1 _3792_ (.A(_1365_),
    .B(_1367_),
    .C(_1369_),
    .D(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__or4_4 _3793_ (.A(_1349_),
    .B(_1355_),
    .C(_1364_),
    .D(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__or4_4 _3794_ (.A(_1333_),
    .B(_1338_),
    .C(_1348_),
    .D(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_1 _3795_ (.A(_0837_),
    .B(_0969_),
    .Y(_1374_));
 sky130_fd_sc_hd__a22o_1 _3796_ (.A1(\hkspi.ldata[0] ),
    .A2(_0969_),
    .B1(_1373_),
    .B2(_1374_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_4 _3797_ (.A(\hkspi.state[3] ),
    .B(\hkspi.state[2] ),
    .X(_1375_));
 sky130_fd_sc_hd__o21a_1 _3798_ (.A1(\hkspi.state[0] ),
    .A2(_1375_),
    .B1(\hkspi.count[0] ),
    .X(_1376_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(\hkspi.count[1] ),
    .B(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__xnor2_1 _3800_ (.A(\hkspi.count[2] ),
    .B(_1377_),
    .Y(_0095_));
 sky130_fd_sc_hd__or2_1 _3801_ (.A(\hkspi.count[1] ),
    .B(_1376_),
    .X(_1378_));
 sky130_fd_sc_hd__and2_1 _3802_ (.A(_1377_),
    .B(_1378_),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _3803_ (.A(\hkspi.count[0] ),
    .B(\hkspi.state[0] ),
    .X(_1379_));
 sky130_fd_sc_hd__o21ba_1 _3804_ (.A1(_1375_),
    .A2(_1379_),
    .B1_N(_1376_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2b_2 _3805_ (.A_N(\hkspi.state[0] ),
    .B(net409),
    .Y(_1380_));
 sky130_fd_sc_hd__and2_2 _3806_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .X(_1381_));
 sky130_fd_sc_hd__and3_4 _3807_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_1382_));
 sky130_fd_sc_hd__nand2_4 _3808_ (.A(\hkspi.count[0] ),
    .B(_1381_),
    .Y(_1383_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(\hkspi.fixed[2] ),
    .B(\hkspi.fixed[1] ),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_2 _3810_ (.A(\hkspi.fixed[0] ),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__a31o_4 _3811_ (.A1(\hkspi.state[2] ),
    .A2(_1382_),
    .A3(_1385_),
    .B1(net409),
    .X(_1386_));
 sky130_fd_sc_hd__nand2b_4 _3812_ (.A_N(\hkspi.state[0] ),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__and3_1 _3813_ (.A(\hkspi.addr[2] ),
    .B(\hkspi.addr[1] ),
    .C(\hkspi.addr[0] ),
    .X(_1388_));
 sky130_fd_sc_hd__and2_2 _3814_ (.A(\hkspi.addr[3] ),
    .B(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__nand4_2 _3815_ (.A(\hkspi.addr[6] ),
    .B(\hkspi.addr[5] ),
    .C(\hkspi.addr[4] ),
    .D(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__mux2_1 _3816_ (.A0(_0844_),
    .A1(_0845_),
    .S(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__nor2_1 _3817_ (.A(_1387_),
    .B(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__a21o_1 _3818_ (.A1(\hkspi.addr[7] ),
    .A2(_1387_),
    .B1(_1392_),
    .X(_0092_));
 sky130_fd_sc_hd__a31o_1 _3819_ (.A1(\hkspi.addr[5] ),
    .A2(\hkspi.addr[4] ),
    .A3(_1389_),
    .B1(\hkspi.addr[6] ),
    .X(_1393_));
 sky130_fd_sc_hd__and3b_1 _3820_ (.A_N(net409),
    .B(_1390_),
    .C(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__a21o_1 _3821_ (.A1(\hkspi.addr[5] ),
    .A2(net409),
    .B1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(_1395_),
    .A1(\hkspi.addr[6] ),
    .S(_1387_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _3823_ (.A(net409),
    .B(_1389_),
    .Y(_1396_));
 sky130_fd_sc_hd__or3b_2 _3824_ (.A(_1387_),
    .B(_1396_),
    .C_N(\hkspi.addr[4] ),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(\hkspi.addr[5] ),
    .B(_1380_),
    .Y(_1398_));
 sky130_fd_sc_hd__xor2_1 _3826_ (.A(_1397_),
    .B(_1398_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _3827_ (.A(net409),
    .B(_1388_),
    .Y(_1399_));
 sky130_fd_sc_hd__mux2_1 _3828_ (.A0(_0839_),
    .A1(_0838_),
    .S(_1389_),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _3829_ (.A0(_1400_),
    .A1(\hkspi.addr[4] ),
    .S(_1387_),
    .X(_0089_));
 sky130_fd_sc_hd__or2_1 _3830_ (.A(\hkspi.addr[3] ),
    .B(_1388_),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_1 _3831_ (.A1(\hkspi.addr[2] ),
    .A2(net409),
    .B1(_1396_),
    .B2(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(_1402_),
    .A1(\hkspi.addr[3] ),
    .S(_1387_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _3833_ (.A1(\hkspi.addr[1] ),
    .A2(\hkspi.addr[0] ),
    .B1(\hkspi.addr[2] ),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _3834_ (.A1(\hkspi.addr[1] ),
    .A2(net409),
    .B1(_1399_),
    .B2(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(_1404_),
    .A1(\hkspi.addr[2] ),
    .S(_1387_),
    .X(_0087_));
 sky130_fd_sc_hd__o211a_1 _3836_ (.A1(_0814_),
    .A2(_1387_),
    .B1(_1380_),
    .C1(\hkspi.addr[1] ),
    .X(_1405_));
 sky130_fd_sc_hd__a21oi_1 _3837_ (.A1(\hkspi.addr[1] ),
    .A2(_1380_),
    .B1(_1387_),
    .Y(_1406_));
 sky130_fd_sc_hd__a21o_1 _3838_ (.A1(\hkspi.addr[0] ),
    .A2(_1406_),
    .B1(_1405_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _3839_ (.A0(_0814_),
    .A1(net58),
    .S(net409),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3840_ (.A0(_1407_),
    .A1(\hkspi.addr[0] ),
    .S(_1387_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(\hkspi.state[0] ),
    .B(_1381_),
    .Y(_1408_));
 sky130_fd_sc_hd__and3_1 _3842_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[0] ),
    .C(\hkspi.state[0] ),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(\hkspi.state[0] ),
    .B(_1382_),
    .Y(_1410_));
 sky130_fd_sc_hd__mux2_1 _3844_ (.A0(\hkspi.pre_pass_thru_user ),
    .A1(\hkspi.pass_thru_user_delay ),
    .S(_1410_),
    .X(_0084_));
 sky130_fd_sc_hd__nor2_8 _3845_ (.A(net409),
    .B(\hkspi.state[0] ),
    .Y(_1411_));
 sky130_fd_sc_hd__a41o_1 _3846_ (.A1(_0818_),
    .A2(\hkspi.state[1] ),
    .A3(_0823_),
    .A4(_1411_),
    .B1(\hkspi.pass_thru_user ),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_2 _3847_ (.A(\hkspi.count[0] ),
    .B(_1408_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2_1 _3848_ (.A0(\hkspi.pass_thru_mgmt_delay ),
    .A1(\hkspi.pre_pass_thru_mgmt ),
    .S(_1412_),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _3849_ (.A1(_0818_),
    .A2(\hkspi.state[4] ),
    .A3(_1411_),
    .B1(\hkspi.pass_thru_mgmt ),
    .X(_0081_));
 sky130_fd_sc_hd__a21oi_1 _3850_ (.A1(\hkspi.readmode ),
    .A2(_1375_),
    .B1(\hkspi.rdstb ),
    .Y(_1413_));
 sky130_fd_sc_hd__a211oi_1 _3851_ (.A1(_1375_),
    .A2(_1383_),
    .B1(_1413_),
    .C1(\hkspi.state[0] ),
    .Y(_0080_));
 sky130_fd_sc_hd__or4b_1 _3852_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .D_N(\hkspi.state[0] ),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(net58),
    .A1(\hkspi.writemode ),
    .S(_1414_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2b_1 _3854_ (.A_N(\hkspi.count[1] ),
    .B(\hkspi.count[0] ),
    .Y(_1415_));
 sky130_fd_sc_hd__or3b_1 _3855_ (.A(_1415_),
    .B(\hkspi.count[2] ),
    .C_N(\hkspi.state[0] ),
    .X(_1416_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(net58),
    .A1(\hkspi.readmode ),
    .S(_1416_),
    .X(_0078_));
 sky130_fd_sc_hd__and4b_4 _3857_ (.A_N(_1381_),
    .B(\hkspi.state[0] ),
    .C(_0837_),
    .D(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__inv_2 _3858_ (.A(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_8 _3859_ (.A(\hkspi.state[2] ),
    .B(_1411_),
    .Y(_1419_));
 sky130_fd_sc_hd__o31a_2 _3860_ (.A1(_1383_),
    .A2(_1384_),
    .A3(_1419_),
    .B1(_1418_),
    .X(_1420_));
 sky130_fd_sc_hd__nor2_2 _3861_ (.A(\hkspi.fixed[0] ),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__a21oi_1 _3862_ (.A1(\hkspi.fixed[2] ),
    .A2(_1421_),
    .B1(_1417_),
    .Y(_1422_));
 sky130_fd_sc_hd__o22a_1 _3863_ (.A1(\hkspi.fixed[2] ),
    .A2(_1417_),
    .B1(_1422_),
    .B2(\hkspi.fixed[1] ),
    .X(_0077_));
 sky130_fd_sc_hd__nor2_1 _3864_ (.A(\hkspi.fixed[1] ),
    .B(_1417_),
    .Y(_1423_));
 sky130_fd_sc_hd__xnor2_1 _3865_ (.A(_1421_),
    .B(_1423_),
    .Y(_0076_));
 sky130_fd_sc_hd__and2b_1 _3866_ (.A_N(\hkspi.state[0] ),
    .B(_1421_),
    .X(_1424_));
 sky130_fd_sc_hd__a221o_1 _3867_ (.A1(net58),
    .A2(_1417_),
    .B1(_1420_),
    .B2(\hkspi.fixed[0] ),
    .C1(_1424_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _3868_ (.A0(\hkspi.odata[6] ),
    .A1(\hkspi.odata[7] ),
    .S(_1419_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(\hkspi.odata[5] ),
    .A1(\hkspi.odata[6] ),
    .S(_1419_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3870_ (.A0(\hkspi.odata[4] ),
    .A1(\hkspi.odata[5] ),
    .S(_1419_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3871_ (.A0(\hkspi.odata[3] ),
    .A1(\hkspi.odata[4] ),
    .S(_1419_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _3872_ (.A0(\hkspi.odata[2] ),
    .A1(\hkspi.odata[3] ),
    .S(_1419_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _3873_ (.A0(\hkspi.odata[1] ),
    .A1(\hkspi.odata[2] ),
    .S(_1419_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(net58),
    .A1(\hkspi.odata[1] ),
    .S(_1419_),
    .X(_0068_));
 sky130_fd_sc_hd__and2b_1 _3875_ (.A_N(\hkspi.count[1] ),
    .B(net58),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\hkspi.pre_pass_thru_mgmt ),
    .A1(_1425_),
    .S(_1409_),
    .X(_0067_));
 sky130_fd_sc_hd__nor3_4 _3877_ (.A(hkspi_disable),
    .B(\gpio_configure[3][3] ),
    .C(net67),
    .Y(_1426_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(net416),
    .B(net411),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _3879_ (.A1(\hkspi.count[0] ),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .B1(_1408_),
    .X(_1427_));
 sky130_fd_sc_hd__a22o_1 _3880_ (.A1(net58),
    .A2(_1412_),
    .B1(_1427_),
    .B2(\hkspi.pre_pass_thru_user ),
    .X(_0066_));
 sky130_fd_sc_hd__o211a_1 _3881_ (.A1(\hkspi.writemode ),
    .A2(\hkspi.wrstb ),
    .B1(\hkspi.state[2] ),
    .C1(_1382_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_8 _3882_ (.A0(serial_clock_pre),
    .A1(serial_bb_clock),
    .S(serial_bb_enable),
    .X(net307));
 sky130_fd_sc_hd__o21a_4 _3883_ (.A1(\hkspi.rdstb ),
    .A2(\hkspi.wrstb ),
    .B1(net412),
    .X(_1428_));
 sky130_fd_sc_hd__o21ai_4 _3884_ (.A1(\hkspi.rdstb ),
    .A2(\hkspi.wrstb ),
    .B1(net412),
    .Y(_1429_));
 sky130_fd_sc_hd__or4_1 _3885_ (.A(net101),
    .B(net100),
    .C(net103),
    .D(net102),
    .X(_1430_));
 sky130_fd_sc_hd__or3_4 _3886_ (.A(net130),
    .B(net129),
    .C(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__or4b_4 _3887_ (.A(net109),
    .B(net108),
    .C(net115),
    .D_N(net116),
    .X(_1432_));
 sky130_fd_sc_hd__or4_2 _3888_ (.A(net105),
    .B(net104),
    .C(net107),
    .D(net106),
    .X(_1433_));
 sky130_fd_sc_hd__and2_2 _3889_ (.A(net112),
    .B(net111),
    .X(_1434_));
 sky130_fd_sc_hd__nand2_4 _3890_ (.A(net112),
    .B(net111),
    .Y(_1435_));
 sky130_fd_sc_hd__or2_4 _3891_ (.A(net114),
    .B(net113),
    .X(_1436_));
 sky130_fd_sc_hd__or4bb_1 _3892_ (.A(net123),
    .B(net122),
    .C_N(net131),
    .D_N(net169),
    .X(_1437_));
 sky130_fd_sc_hd__or4bb_1 _3893_ (.A(net118),
    .B(net119),
    .C_N(net120),
    .D_N(net117),
    .X(_1438_));
 sky130_fd_sc_hd__or4_4 _3894_ (.A(_1434_),
    .B(_1436_),
    .C(_1437_),
    .D(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__nor4_4 _3895_ (.A(_1431_),
    .B(_1432_),
    .C(_1433_),
    .D(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__nand2_1 _3896_ (.A(\wbbd_state[0] ),
    .B(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__a22o_1 _3897_ (.A1(\wbbd_state[5] ),
    .A2(_1428_),
    .B1(_1440_),
    .B2(\wbbd_state[0] ),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _3898_ (.A(_1383_),
    .B(_1385_),
    .Y(_1442_));
 sky130_fd_sc_hd__a22o_1 _3899_ (.A1(\hkspi.state[0] ),
    .A2(_1383_),
    .B1(_1442_),
    .B2(\hkspi.state[2] ),
    .X(_0004_));
 sky130_fd_sc_hd__a21o_1 _3900_ (.A1(\wbbd_state[9] ),
    .A2(_1428_),
    .B1(\wbbd_state[4] ),
    .X(_0013_));
 sky130_fd_sc_hd__nand2b_4 _3901_ (.A_N(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_1443_));
 sky130_fd_sc_hd__and2b_4 _3902_ (.A_N(\pad_count_2[0] ),
    .B(\pad_count_2[1] ),
    .X(_1444_));
 sky130_fd_sc_hd__and2b_4 _3903_ (.A_N(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .X(_1445_));
 sky130_fd_sc_hd__nand2_8 _3904_ (.A(_1444_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__or2_4 _3905_ (.A(_1443_),
    .B(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__nor2_1 _3906_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .Y(_1448_));
 sky130_fd_sc_hd__and4b_4 _3907_ (.A_N(net307),
    .B(_1448_),
    .C(\xfer_count[2] ),
    .D(\xfer_count[3] ),
    .X(_1449_));
 sky130_fd_sc_hd__nor2_4 _3908_ (.A(net405),
    .B(net307),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(net407),
    .B(_1449_),
    .Y(_1451_));
 sky130_fd_sc_hd__a32o_1 _3910_ (.A1(net407),
    .A2(_1447_),
    .A3(_1449_),
    .B1(serial_xfer),
    .B2(\xfer_state[0] ),
    .X(_0016_));
 sky130_fd_sc_hd__or4b_2 _3911_ (.A(\xfer_count[0] ),
    .B(\xfer_count[2] ),
    .C(\xfer_count[3] ),
    .D_N(\xfer_count[1] ),
    .X(_1452_));
 sky130_fd_sc_hd__a2bb2o_1 _3912_ (.A1_N(_1447_),
    .A2_N(_1451_),
    .B1(_1452_),
    .B2(\xfer_state[3] ),
    .X(_0017_));
 sky130_fd_sc_hd__a21o_1 _3913_ (.A1(\wbbd_state[7] ),
    .A2(_1428_),
    .B1(\wbbd_state[2] ),
    .X(_0011_));
 sky130_fd_sc_hd__a21o_1 _3914_ (.A1(\wbbd_state[8] ),
    .A2(_1428_),
    .B1(\wbbd_state[3] ),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _3915_ (.A(_0816_),
    .B(_1440_),
    .X(_1453_));
 sky130_fd_sc_hd__nand2_1 _3916_ (.A(_0817_),
    .B(_1453_),
    .Y(_0009_));
 sky130_fd_sc_hd__a41o_1 _3917_ (.A1(\hkspi.pre_pass_thru_user ),
    .A2(_0815_),
    .A3(\hkspi.state[0] ),
    .A4(_1382_),
    .B1(\hkspi.state[1] ),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _3918_ (.A(_0821_),
    .B(_1452_),
    .X(_1454_));
 sky130_fd_sc_hd__o21ai_1 _3919_ (.A1(serial_xfer),
    .A2(_0820_),
    .B1(_1454_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(net407),
    .B(net307),
    .Y(_1455_));
 sky130_fd_sc_hd__nor2_1 _3921_ (.A(net405),
    .B(_1449_),
    .Y(_1456_));
 sky130_fd_sc_hd__or2_1 _3922_ (.A(\xfer_state[2] ),
    .B(_1456_),
    .X(_0015_));
 sky130_fd_sc_hd__a31o_1 _3923_ (.A1(\hkspi.pre_pass_thru_mgmt ),
    .A2(\hkspi.state[0] ),
    .A3(_1382_),
    .B1(\hkspi.state[4] ),
    .X(_0008_));
 sky130_fd_sc_hd__or3_1 _3924_ (.A(\hkspi.pre_pass_thru_user ),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .C(_1410_),
    .X(_1457_));
 sky130_fd_sc_hd__a21bo_1 _3925_ (.A1(\hkspi.state[3] ),
    .A2(_1383_),
    .B1_N(_1457_),
    .X(_0007_));
 sky130_fd_sc_hd__a2bb2o_1 _3926_ (.A1_N(_0818_),
    .A2_N(_1442_),
    .B1(_1382_),
    .B2(\hkspi.state[3] ),
    .X(_0006_));
 sky130_fd_sc_hd__o21ai_1 _3927_ (.A1(\hkspi.state[1] ),
    .A2(\hkspi.state[4] ),
    .B1(_0818_),
    .Y(_1458_));
 sky130_fd_sc_hd__and2_1 _3928_ (.A(_0969_),
    .B(_1458_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_8 _3929_ (.A0(\mgmt_gpio_data[37] ),
    .A1(net91),
    .S(net76),
    .X(net243));
 sky130_fd_sc_hd__mux2_8 _3930_ (.A0(\mgmt_gpio_data[36] ),
    .A1(net89),
    .S(net76),
    .X(net242));
 sky130_fd_sc_hd__mux2_8 _3931_ (.A0(_0825_),
    .A1(net92),
    .S(net76),
    .X(net205));
 sky130_fd_sc_hd__mux2_8 _3932_ (.A0(_0826_),
    .A1(net90),
    .S(net76),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _3933_ (.A0(_0827_),
    .A1(net82),
    .S(net79),
    .X(net203));
 sky130_fd_sc_hd__mux2_8 _3934_ (.A0(\mgmt_gpio_data[32] ),
    .A1(net80),
    .S(net79),
    .X(net238));
 sky130_fd_sc_hd__mux2_8 _3935_ (.A0(\mgmt_gpio_data[33] ),
    .A1(net78),
    .S(net79),
    .X(net239));
 sky130_fd_sc_hd__mux2_8 _3936_ (.A0(\mgmt_gpio_data[35] ),
    .A1(net81),
    .S(net79),
    .X(net241));
 sky130_fd_sc_hd__mux2_2 _3937_ (.A0(\mgmt_gpio_data[10] ),
    .A1(net58),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net214));
 sky130_fd_sc_hd__mux2_1 _3938_ (.A0(\mgmt_gpio_data[9] ),
    .A1(clknet_2_3_0_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_user ),
    .X(net250));
 sky130_fd_sc_hd__mux2_2 _3939_ (.A0(\mgmt_gpio_data[8] ),
    .A1(net67),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net249));
 sky130_fd_sc_hd__mux2_8 _3940_ (.A0(\mgmt_gpio_data[6] ),
    .A1(net77),
    .S(net94),
    .X(net247));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(\mgmt_gpio_data[1] ),
    .A1(\hkspi.SDO ),
    .S(net411),
    .X(_1459_));
 sky130_fd_sc_hd__or2_1 _3942_ (.A(\hkspi.pass_thru_user ),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a21oi_2 _3943_ (.A1(\hkspi.pass_thru_user ),
    .A2(_0824_),
    .B1(\hkspi.pass_thru_mgmt ),
    .Y(_1461_));
 sky130_fd_sc_hd__a22o_4 _3944_ (.A1(\hkspi.pass_thru_mgmt ),
    .A2(net74),
    .B1(_1460_),
    .B2(_1461_),
    .X(net224));
 sky130_fd_sc_hd__mux2_8 _3945_ (.A0(\mgmt_gpio_data[0] ),
    .A1(net3),
    .S(net1),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _3946_ (.A0(_0828_),
    .A1(\hkspi.sdoenb ),
    .S(net412),
    .X(net186));
 sky130_fd_sc_hd__mux2_8 _3947_ (.A0(_0829_),
    .A1(net2),
    .S(net1),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _3948_ (.A0(\mgmt_gpio_data[15] ),
    .A1(user_clock),
    .S(clk2_output_dest),
    .X(net219));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\mgmt_gpio_data[14] ),
    .A1(clknet_3_7_0_wb_clk_i),
    .S(clk1_output_dest),
    .X(net218));
 sky130_fd_sc_hd__mux2_8 _3950_ (.A0(\mgmt_gpio_data[13] ),
    .A1(net93),
    .S(trap_output_dest),
    .X(net217));
 sky130_fd_sc_hd__mux2_4 _3951_ (.A0(serial_resetn_pre),
    .A1(serial_bb_resetn),
    .S(serial_bb_enable),
    .X(net311));
 sky130_fd_sc_hd__mux2_2 _3952_ (.A0(serial_load_pre),
    .A1(serial_bb_load),
    .S(serial_bb_enable),
    .X(net310));
 sky130_fd_sc_hd__nor2_2 _3953_ (.A(net406),
    .B(net462),
    .Y(_1462_));
 sky130_fd_sc_hd__a22o_2 _3954_ (.A1(net406),
    .A2(clknet_1_0__leaf_wbbd_sck),
    .B1(net411),
    .B2(_1462_),
    .X(csclk));
 sky130_fd_sc_hd__mux2_8 _3955_ (.A0(net84),
    .A1(net67),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net253));
 sky130_fd_sc_hd__nor2_1 _3956_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(net415),
    .Y(net254));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(net83),
    .A1(clknet_2_0_0_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_mgmt ),
    .X(net251));
 sky130_fd_sc_hd__nor2_1 _3958_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net415),
    .Y(net252));
 sky130_fd_sc_hd__nand2b_4 _3959_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net86),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(net256),
    .Y(net257));
 sky130_fd_sc_hd__or2_4 _3961_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net88),
    .X(net260));
 sky130_fd_sc_hd__inv_2 _3962_ (.A(net260),
    .Y(net259));
 sky130_fd_sc_hd__mux2_8 _3963_ (.A0(net85),
    .A1(net58),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net255));
 sky130_fd_sc_hd__and2b_4 _3964_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net73),
    .X(net313));
 sky130_fd_sc_hd__and2b_4 _3965_ (.A_N(\hkspi.pass_thru_mgmt ),
    .B(net74),
    .X(net314));
 sky130_fd_sc_hd__and2_1 _3966_ (.A(\wbbd_state[7] ),
    .B(_1429_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(\wbbd_state[5] ),
    .B(_1429_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _3968_ (.A(\wbbd_state[8] ),
    .B(_1429_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_2 _3969_ (.A(net68),
    .B(net94),
    .X(net306));
 sky130_fd_sc_hd__and2_2 _3970_ (.A(net63),
    .B(net79),
    .X(net312));
 sky130_fd_sc_hd__and2_2 _3971_ (.A(net36),
    .B(net1),
    .X(net171));
 sky130_fd_sc_hd__and2_2 _3972_ (.A(irq_1_inputsrc),
    .B(net70),
    .X(net173));
 sky130_fd_sc_hd__and2_4 _3973_ (.A(irq_2_inputsrc),
    .B(net39),
    .X(net174));
 sky130_fd_sc_hd__and2_1 _3974_ (.A(\wbbd_state[9] ),
    .B(_1429_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2b_4 _3975_ (.A_N(net616),
    .B(net676),
    .Y(_1463_));
 sky130_fd_sc_hd__o21a_4 _3976_ (.A1(net560),
    .A2(net406),
    .B1(net617),
    .X(_1464_));
 sky130_fd_sc_hd__o21ai_4 _3977_ (.A1(net560),
    .A2(net676),
    .B1(net617),
    .Y(_1465_));
 sky130_fd_sc_hd__and2_4 _3978_ (.A(_0924_),
    .B(net509),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_8 _3979_ (.A0(net58),
    .A1(net1345),
    .S(net675),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(net1665),
    .A1(net400),
    .S(_1466_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_8 _3981_ (.A0(net527),
    .A1(net621),
    .S(net406),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(net1382),
    .A1(net394),
    .S(_1466_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_4 _3983_ (.A0(net501),
    .A1(\wbbd_data[2] ),
    .S(wbbd_busy),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(net1459),
    .A1(net388),
    .S(_1466_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_8 _3985_ (.A0(net595),
    .A1(net613),
    .S(wbbd_busy),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(net1467),
    .A1(net383),
    .S(_1466_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_8 _3987_ (.A0(net643),
    .A1(net662),
    .S(wbbd_busy),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(net932),
    .A1(net379),
    .S(_1466_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_4 _3989_ (.A0(net536),
    .A1(\wbbd_data[5] ),
    .S(net406),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_1 _3990_ (.A0(net1075),
    .A1(net375),
    .S(_1466_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_8 _3991_ (.A0(net667),
    .A1(\wbbd_data[6] ),
    .S(net406),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(net1088),
    .A1(net372),
    .S(_1466_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_8 _3993_ (.A0(net472),
    .A1(\wbbd_data[7] ),
    .S(wbbd_busy),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _3994_ (.A0(net870),
    .A1(net369),
    .S(_1466_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_4 _3995_ (.A(net688),
    .B(net362),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(net1681),
    .A1(net399),
    .S(_1475_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3997_ (.A0(net1371),
    .A1(net394),
    .S(_1475_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(net1500),
    .A1(net388),
    .S(_1475_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(net1478),
    .A1(net383),
    .S(_1475_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(net1231),
    .A1(net379),
    .S(_1475_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4001_ (.A0(net1081),
    .A1(net375),
    .S(_1475_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4002_ (.A0(net297),
    .A1(net671),
    .S(_1475_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(net950),
    .A1(net369),
    .S(_1475_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(_1249_),
    .B(net363),
    .Y(_1476_));
 sky130_fd_sc_hd__mux2_1 _4005_ (.A0(net400),
    .A1(net1523),
    .S(_1476_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4006_ (.A0(net396),
    .A1(net292),
    .S(_1476_),
    .X(_0113_));
 sky130_fd_sc_hd__and2b_4 _4007_ (.A_N(net413),
    .B(_0911_),
    .X(_1477_));
 sky130_fd_sc_hd__o221a_4 _4008_ (.A1(net482),
    .A2(net413),
    .B1(_1477_),
    .B2(_0899_),
    .C1(net562),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(net1699),
    .A1(net1347),
    .S(_0899_),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _4010_ (.A0(net1410),
    .A1(_1479_),
    .S(_1478_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(net783),
    .A1(net398),
    .S(_0899_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _4012_ (.A0(net1181),
    .A1(_1480_),
    .S(_1478_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(net987),
    .A1(net392),
    .S(_0899_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(net1338),
    .A1(_1481_),
    .S(_1478_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(net1177),
    .A1(net386),
    .S(_0899_),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(net1405),
    .A1(_1482_),
    .S(_1478_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(net729),
    .A1(net382),
    .S(_0899_),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(net1232),
    .A1(_1483_),
    .S(_1478_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(net873),
    .A1(net376),
    .S(_0899_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _4020_ (.A0(net1264),
    .A1(_1484_),
    .S(_1478_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(net1696),
    .A1(net373),
    .S(_0899_),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(net1351),
    .A1(_1485_),
    .S(_1478_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(net817),
    .A1(net476),
    .S(_0899_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(net743),
    .A1(_1486_),
    .S(_1478_),
    .X(_0121_));
 sky130_fd_sc_hd__nand2_8 _4025_ (.A(_0911_),
    .B(net366),
    .Y(_1487_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(net402),
    .A1(net1444),
    .S(_1487_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(net398),
    .A1(net771),
    .S(_1487_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(net392),
    .A1(net971),
    .S(_1487_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(net533),
    .A1(net627),
    .S(_1487_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(net382),
    .A1(net714),
    .S(_1487_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(net376),
    .A1(net846),
    .S(_1487_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(net373),
    .A1(net999),
    .S(_1487_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(net370),
    .A1(net781),
    .S(_1487_),
    .X(_0129_));
 sky130_fd_sc_hd__or4_4 _4034_ (.A(net482),
    .B(net358),
    .C(net413),
    .D(net677),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(net1347),
    .A1(net1699),
    .S(_1488_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(net398),
    .A1(net783),
    .S(_1488_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(net392),
    .A1(net987),
    .S(_1488_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(net386),
    .A1(net1177),
    .S(_1488_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(net382),
    .A1(net729),
    .S(_1488_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(net376),
    .A1(net873),
    .S(_1488_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(net592),
    .A1(net1696),
    .S(_1488_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(net370),
    .A1(net817),
    .S(_1488_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_4 _4043_ (.A(_1069_),
    .B(net362),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(net1692),
    .A1(net399),
    .S(_1489_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4045_ (.A0(net1361),
    .A1(net394),
    .S(_1489_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(net1460),
    .A1(net388),
    .S(_1489_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(net1254),
    .A1(net384),
    .S(_1489_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(net1519),
    .A1(net378),
    .S(_1489_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_4 _4049_ (.A(_1094_),
    .B(net362),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(net1675),
    .A1(net400),
    .S(_1490_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(net1353),
    .A1(net394),
    .S(_1490_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(net1136),
    .A1(net389),
    .S(_1490_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4053_ (.A0(net1451),
    .A1(net383),
    .S(_1490_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(net1518),
    .A1(net378),
    .S(_1490_),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_8 _4055_ (.A(_1127_),
    .B(net365),
    .Y(_1491_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(net403),
    .A1(net1561),
    .S(_1491_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(net394),
    .A1(net1355),
    .S(_1491_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(net390),
    .A1(net1653),
    .S(_1491_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(net383),
    .A1(net1468),
    .S(_1491_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(net378),
    .A1(net1510),
    .S(_1491_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_8 _4061_ (.A(_1068_),
    .B(net365),
    .Y(_1492_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(net403),
    .A1(net1589),
    .S(_1492_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(net397),
    .A1(net785),
    .S(_1492_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(net391),
    .A1(net1420),
    .S(_1492_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(net384),
    .A1(net1248),
    .S(_1492_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(net378),
    .A1(net1505),
    .S(_1492_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_4 _4067_ (.A(_1057_),
    .B(net365),
    .Y(_1493_));
 sky130_fd_sc_hd__mux2_1 _4068_ (.A0(net403),
    .A1(net1583),
    .S(_1493_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(net397),
    .A1(net1119),
    .S(_1493_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4070_ (.A0(net390),
    .A1(net1580),
    .S(_1493_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(net533),
    .A1(net767),
    .S(_1493_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(net381),
    .A1(net1340),
    .S(_1493_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_4 _4073_ (.A(\wbbd_state[4] ),
    .B(net457),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(net325),
    .A1(_1373_),
    .S(_1494_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(net326),
    .A1(_1308_),
    .S(_1494_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(net327),
    .A1(_1247_),
    .S(_1494_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(net328),
    .A1(_1189_),
    .S(_1494_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(net330),
    .A1(clknet_1_1__leaf__1132_),
    .S(_1494_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(net331),
    .A1(_1037_),
    .S(_1494_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(net332),
    .A1(_1002_),
    .S(_1494_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net333),
    .A1(_0968_),
    .S(_1494_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_4 _4082_ (.A(_1065_),
    .B(net365),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(net1641),
    .A1(net403),
    .S(_1495_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(net806),
    .A1(net397),
    .S(_1495_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(net1448),
    .A1(net391),
    .S(_1495_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _4086_ (.A0(net1710),
    .A1(net533),
    .S(_1495_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4087_ (.A0(net673),
    .A1(net382),
    .S(_1495_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_4 _4088_ (.A(\wbbd_state[2] ),
    .B(net457),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(net348),
    .A1(_1373_),
    .S(_1496_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(net349),
    .A1(_1308_),
    .S(_1496_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(net319),
    .A1(_1247_),
    .S(_1496_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(net320),
    .A1(_1189_),
    .S(_1496_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(net321),
    .A1(clknet_1_1__leaf__1132_),
    .S(_1496_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _4094_ (.A0(net322),
    .A1(_1037_),
    .S(_1496_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _4095_ (.A0(net323),
    .A1(_1002_),
    .S(_1496_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(net324),
    .A1(_0968_),
    .S(_1496_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_4 _4097_ (.A(_1115_),
    .B(net509),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(net400),
    .A1(net1587),
    .S(_1497_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(net395),
    .A1(net957),
    .S(_1497_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(net389),
    .A1(net1140),
    .S(_1497_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _4101_ (.A0(net384),
    .A1(net1242),
    .S(_1497_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(net378),
    .A1(net1501),
    .S(_1497_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_4 _4103_ (.A(\wbbd_state[3] ),
    .B(net457),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _4104_ (.A0(net318),
    .A1(_1373_),
    .S(_1498_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(net329),
    .A1(_1308_),
    .S(_1498_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(net340),
    .A1(_1247_),
    .S(_1498_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(net343),
    .A1(_1189_),
    .S(_1498_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(net344),
    .A1(clknet_1_0__leaf__1132_),
    .S(_1498_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(net345),
    .A1(_1037_),
    .S(_1498_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(net346),
    .A1(_1002_),
    .S(_1498_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(net347),
    .A1(_0968_),
    .S(_1498_),
    .X(_0196_));
 sky130_fd_sc_hd__nand2_8 _4112_ (.A(_1113_),
    .B(net365),
    .Y(_1499_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(net403),
    .A1(net1600),
    .S(_1499_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(net395),
    .A1(net1019),
    .S(_1499_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4115_ (.A0(net391),
    .A1(net1414),
    .S(_1499_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(net384),
    .A1(net1291),
    .S(_1499_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(net378),
    .A1(net1527),
    .S(_1499_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_4 _4118_ (.A(_1064_),
    .B(net509),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(net1667),
    .A1(net400),
    .S(_1500_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4120_ (.A0(net975),
    .A1(net395),
    .S(_1500_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(net1174),
    .A1(net389),
    .S(_1500_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(net1223),
    .A1(net384),
    .S(_1500_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(net1492),
    .A1(net378),
    .S(_1500_),
    .X(_0206_));
 sky130_fd_sc_hd__and2_4 _4124_ (.A(_1102_),
    .B(net365),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _4125_ (.A0(net1591),
    .A1(net403),
    .S(_1501_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(net993),
    .A1(net397),
    .S(_1501_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(net1597),
    .A1(net390),
    .S(_1501_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(net694),
    .A1(net533),
    .S(_1501_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(net1268),
    .A1(net381),
    .S(_1501_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_8 _4130_ (.A(_1039_),
    .B(net509),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _4131_ (.A0(net403),
    .A1(net1602),
    .S(_1502_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4132_ (.A0(net395),
    .A1(net965),
    .S(_1502_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _4133_ (.A0(net391),
    .A1(net1417),
    .S(_1502_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4134_ (.A0(net384),
    .A1(net1512),
    .S(_1502_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(net378),
    .A1(net1514),
    .S(_1502_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_4 _4136_ (.A(_1073_),
    .B(net365),
    .Y(_1503_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(net403),
    .A1(net1571),
    .S(_1503_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(net397),
    .A1(net1143),
    .S(_1503_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(net390),
    .A1(net1578),
    .S(_1503_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(net533),
    .A1(net704),
    .S(_1503_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4141_ (.A0(net381),
    .A1(net1256),
    .S(_1503_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_8 _4142_ (.A(net792),
    .B(net365),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_1 _4143_ (.A0(net403),
    .A1(net1629),
    .S(_1504_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(net397),
    .A1(net1706),
    .S(_1504_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _4145_ (.A0(net391),
    .A1(net1441),
    .S(_1504_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(net384),
    .A1(net1270),
    .S(_1504_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(net378),
    .A1(net1525),
    .S(_1504_),
    .X(_0226_));
 sky130_fd_sc_hd__and2_4 _4148_ (.A(_1062_),
    .B(net365),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(net1606),
    .A1(net403),
    .S(_1505_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(net1099),
    .A1(net397),
    .S(_1505_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(net1412),
    .A1(net391),
    .S(_1505_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(net1279),
    .A1(net384),
    .S(_1505_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _4153_ (.A0(net1711),
    .A1(net382),
    .S(_1505_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_4 _4154_ (.A(_1041_),
    .B(net365),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _4155_ (.A0(net1555),
    .A1(net403),
    .S(_1506_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(net997),
    .A1(net397),
    .S(_1506_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _4157_ (.A0(net1579),
    .A1(net390),
    .S(_1506_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(net774),
    .A1(net533),
    .S(_1506_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _4159_ (.A0(net1277),
    .A1(net381),
    .S(_1506_),
    .X(_0236_));
 sky130_fd_sc_hd__nand2_8 _4160_ (.A(_1112_),
    .B(net365),
    .Y(_1507_));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(net403),
    .A1(net1635),
    .S(_1507_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(net395),
    .A1(net1057),
    .S(_1507_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(net391),
    .A1(net1430),
    .S(_1507_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(net533),
    .A1(net838),
    .S(_1507_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _4165_ (.A0(net378),
    .A1(net1559),
    .S(_1507_),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_4 _4166_ (.A(_1084_),
    .B(net362),
    .Y(_1508_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(net399),
    .A1(net1616),
    .S(_1508_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _4168_ (.A0(net394),
    .A1(net1357),
    .S(_1508_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(net388),
    .A1(net1471),
    .S(_1508_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(net383),
    .A1(net1428),
    .S(_1508_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(net379),
    .A1(net1216),
    .S(_1508_),
    .X(_0246_));
 sky130_fd_sc_hd__and2_4 _4172_ (.A(_1089_),
    .B(net362),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(net1690),
    .A1(net399),
    .S(_1509_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(net1372),
    .A1(net394),
    .S(_1509_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(net1454),
    .A1(net388),
    .S(_1509_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(net1481),
    .A1(net383),
    .S(_1509_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(net1206),
    .A1(net379),
    .S(_1509_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_4 _4178_ (.A(_1085_),
    .B(net509),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(net1684),
    .A1(net400),
    .S(_1510_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(net1069),
    .A1(net395),
    .S(_1510_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(net1565),
    .A1(net388),
    .S(_1510_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(net1323),
    .A1(net384),
    .S(_1510_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(net1563),
    .A1(net378),
    .S(_1510_),
    .X(_0256_));
 sky130_fd_sc_hd__and2_4 _4184_ (.A(_1052_),
    .B(net365),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(net1604),
    .A1(net403),
    .S(_1511_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(net804),
    .A1(net397),
    .S(_1511_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(net1151),
    .A1(net389),
    .S(_1511_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(net1266),
    .A1(net384),
    .S(_1511_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(net1520),
    .A1(net378),
    .S(_1511_),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_4 _4190_ (.A(_1048_),
    .B(net362),
    .Y(_1512_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(net399),
    .A1(net1627),
    .S(_1512_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(net394),
    .A1(net1359),
    .S(_1512_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(net388),
    .A1(net1464),
    .S(_1512_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(net383),
    .A1(net1434),
    .S(_1512_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net379),
    .A1(net1193),
    .S(_1512_),
    .X(_0266_));
 sky130_fd_sc_hd__nand2_4 _4196_ (.A(_1078_),
    .B(net362),
    .Y(_1513_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(net399),
    .A1(net1639),
    .S(_1513_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(net394),
    .A1(net1402),
    .S(_1513_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net388),
    .A1(net1494),
    .S(_1513_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(net383),
    .A1(net1495),
    .S(_1513_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net379),
    .A1(net1283),
    .S(_1513_),
    .X(_0271_));
 sky130_fd_sc_hd__o221a_4 _4202_ (.A1(_0917_),
    .A2(net413),
    .B1(_1477_),
    .B2(_0918_),
    .C1(net366),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net1418),
    .A1(net1347),
    .S(_0918_),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _4204_ (.A0(net1415),
    .A1(_1515_),
    .S(_1514_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net779),
    .A1(net398),
    .S(_0918_),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(net1189),
    .A1(_1516_),
    .S(_1514_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(net1016),
    .A1(net392),
    .S(_0918_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(net1349),
    .A1(_1517_),
    .S(_1514_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net1103),
    .A1(net386),
    .S(_0918_),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(net1378),
    .A1(_1518_),
    .S(_1514_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net920),
    .A1(net382),
    .S(_0918_),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(net1702),
    .A1(net921),
    .S(_1514_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(net1698),
    .A1(net540),
    .S(_0918_),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(net735),
    .A1(_1520_),
    .S(_1514_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(net983),
    .A1(net373),
    .S(_0918_),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(net1336),
    .A1(_1521_),
    .S(_1514_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(net1701),
    .A1(net476),
    .S(_0918_),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(net716),
    .A1(_1522_),
    .S(_1514_),
    .X(_0279_));
 sky130_fd_sc_hd__o221a_4 _4219_ (.A1(_0932_),
    .A2(net412),
    .B1(_1477_),
    .B2(_0950_),
    .C1(net509),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(net1425),
    .A1(net399),
    .S(_0950_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(net1688),
    .A1(_1524_),
    .S(_1523_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _4222_ (.A0(net1374),
    .A1(net394),
    .S(_0950_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(net1543),
    .A1(_1525_),
    .S(_1523_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(net1149),
    .A1(net389),
    .S(_0950_),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(net1383),
    .A1(_1526_),
    .S(_1523_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(net1700),
    .A1(net598),
    .S(_0950_),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net908),
    .A1(_1527_),
    .S(_1523_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _4228_ (.A0(net755),
    .A1(net631),
    .S(_0950_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(net1010),
    .A1(_1528_),
    .S(_1523_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net1162),
    .A1(net375),
    .S(_0950_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(net1392),
    .A1(_1529_),
    .S(_1523_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _4232_ (.A0(net708),
    .A1(net592),
    .S(_0950_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _4233_ (.A0(net985),
    .A1(_1530_),
    .S(_1523_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(net891),
    .A1(net369),
    .S(_0950_),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(net1309),
    .A1(_1531_),
    .S(_1523_),
    .X(_0287_));
 sky130_fd_sc_hd__nor3_4 _4236_ (.A(\wbbd_state[8] ),
    .B(\wbbd_state[7] ),
    .C(\wbbd_state[9] ),
    .Y(_1532_));
 sky130_fd_sc_hd__or4_2 _4237_ (.A(\wbbd_state[2] ),
    .B(\wbbd_state[1] ),
    .C(\wbbd_state[3] ),
    .D(\wbbd_state[4] ),
    .X(_1533_));
 sky130_fd_sc_hd__and2b_4 _4238_ (.A_N(\wbbd_state[5] ),
    .B(_1532_),
    .X(_1534_));
 sky130_fd_sc_hd__or4_4 _4239_ (.A(\wbbd_state[5] ),
    .B(\wbbd_state[8] ),
    .C(\wbbd_state[7] ),
    .D(\wbbd_state[9] ),
    .X(_1535_));
 sky130_fd_sc_hd__a2111o_1 _4240_ (.A1(_0816_),
    .A2(net406),
    .B1(\wbbd_state[6] ),
    .C1(_1533_),
    .D1(_1535_),
    .X(_0288_));
 sky130_fd_sc_hd__or4_4 _4241_ (.A(net358),
    .B(_0917_),
    .C(net413),
    .D(net1275),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(net403),
    .A1(net1418),
    .S(_1536_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(net398),
    .A1(net779),
    .S(_1536_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net392),
    .A1(net1016),
    .S(_1536_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(net386),
    .A1(net1103),
    .S(_1536_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(net381),
    .A1(net920),
    .S(_1536_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(net469),
    .A1(net1698),
    .S(_1536_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(net373),
    .A1(net983),
    .S(_1536_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(net465),
    .A1(net1701),
    .S(_1536_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_4 _4250_ (.A(_1123_),
    .B(net365),
    .Y(_1537_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(net400),
    .A1(net1625),
    .S(_1537_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(net395),
    .A1(net951),
    .S(_1537_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net389),
    .A1(net1152),
    .S(_1537_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(net384),
    .A1(net1234),
    .S(_1537_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(net378),
    .A1(net1508),
    .S(_1537_),
    .X(_0301_));
 sky130_fd_sc_hd__and2_4 _4256_ (.A(_1046_),
    .B(net509),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(net1679),
    .A1(net400),
    .S(_1538_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(net989),
    .A1(net395),
    .S(_1538_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(net1329),
    .A1(net391),
    .S(_1538_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(net1204),
    .A1(net384),
    .S(_1538_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net1498),
    .A1(net378),
    .S(_1538_),
    .X(_0306_));
 sky130_fd_sc_hd__and2_4 _4262_ (.A(_1118_),
    .B(net365),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net1612),
    .A1(net403),
    .S(_1539_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(net1073),
    .A1(net395),
    .S(_1539_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net1631),
    .A1(net390),
    .S(_1539_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(net1303),
    .A1(net384),
    .S(_1539_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net1664),
    .A1(net378),
    .S(_1539_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_4 _4268_ (.A(_1124_),
    .B(net562),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net1531),
    .A1(net403),
    .S(_1540_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(net1071),
    .A1(net395),
    .S(_1540_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(net1404),
    .A1(net391),
    .S(_1540_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(net1332),
    .A1(net384),
    .S(_1540_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(net1334),
    .A1(net379),
    .S(_1540_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_4 _4274_ (.A(_1077_),
    .B(net362),
    .Y(_1541_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(net399),
    .A1(net1637),
    .S(_1541_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(net394),
    .A1(net1396),
    .S(_1541_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(net388),
    .A1(net1497),
    .S(_1541_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(net383),
    .A1(net1479),
    .S(_1541_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(net379),
    .A1(net1250),
    .S(_1541_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_8 _4280_ (.A(_1104_),
    .B(net562),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(net403),
    .A1(net1367),
    .S(_1542_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(net395),
    .A1(net1028),
    .S(_1542_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(net390),
    .A1(net1409),
    .S(_1542_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(net384),
    .A1(net1327),
    .S(_1542_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(net378),
    .A1(net1387),
    .S(_1542_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_4 _4286_ (.A(_1090_),
    .B(net362),
    .Y(_1543_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(net400),
    .A1(net1656),
    .S(_1543_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(net395),
    .A1(net875),
    .S(_1543_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(net388),
    .A1(net1466),
    .S(_1543_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(net383),
    .A1(net1452),
    .S(_1543_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(net379),
    .A1(net1201),
    .S(_1543_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_8 _4292_ (.A(_1108_),
    .B(net365),
    .Y(_1544_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(net403),
    .A1(net1581),
    .S(_1544_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(net395),
    .A1(net1030),
    .S(_1544_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(net390),
    .A1(net1624),
    .S(_1544_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net384),
    .A1(net1297),
    .S(_1544_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(net378),
    .A1(net1566),
    .S(_1544_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _4298_ (.A(_1051_),
    .B(net362),
    .Y(_1545_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(net399),
    .A1(net1654),
    .S(_1545_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(net394),
    .A1(net1369),
    .S(_1545_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(net388),
    .A1(net1470),
    .S(_1545_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(net383),
    .A1(net1455),
    .S(_1545_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(net379),
    .A1(net1210),
    .S(_1545_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_4 _4304_ (.A(_1092_),
    .B(net362),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(net1682),
    .A1(net400),
    .S(_1546_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(net959),
    .A1(net395),
    .S(_1546_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(net1552),
    .A1(net388),
    .S(_1546_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(net1550),
    .A1(net383),
    .S(_1546_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(net1293),
    .A1(net379),
    .S(_1546_),
    .X(_0346_));
 sky130_fd_sc_hd__and2_4 _4310_ (.A(_1054_),
    .B(net509),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(net1673),
    .A1(net400),
    .S(_1547_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(net915),
    .A1(net395),
    .S(_1547_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(net1507),
    .A1(net388),
    .S(_1547_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(net1260),
    .A1(net384),
    .S(_1547_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(net1225),
    .A1(net379),
    .S(_1547_),
    .X(_0351_));
 sky130_fd_sc_hd__and2_4 _4316_ (.A(_1043_),
    .B(net362),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(net1694),
    .A1(net399),
    .S(_1548_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(net1376),
    .A1(net394),
    .S(_1548_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(net1490),
    .A1(net388),
    .S(_1548_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(net1474),
    .A1(net383),
    .S(_1548_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(net1484),
    .A1(net378),
    .S(_1548_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_4 _4322_ (.A(_1098_),
    .B(net362),
    .Y(_1549_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(net400),
    .A1(net1677),
    .S(_1549_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(net395),
    .A1(net963),
    .S(_1549_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(net388),
    .A1(net1558),
    .S(_1549_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(net384),
    .A1(net1262),
    .S(_1549_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(net379),
    .A1(net1252),
    .S(_1549_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_4 _4328_ (.A(_1044_),
    .B(net509),
    .Y(_1550_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(net399),
    .A1(net1576),
    .S(_1550_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(net394),
    .A1(net1390),
    .S(_1550_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(net389),
    .A1(net1131),
    .S(_1550_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(net383),
    .A1(net1462),
    .S(_1550_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(net378),
    .A1(net1516),
    .S(_1550_),
    .X(_0366_));
 sky130_fd_sc_hd__and2_4 _4334_ (.A(net459),
    .B(net125),
    .X(_1551_));
 sky130_fd_sc_hd__nand2_8 _4335_ (.A(net459),
    .B(net125),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_8 _4336_ (.A(net124),
    .B(net121),
    .Y(_1553_));
 sky130_fd_sc_hd__and3_4 _4337_ (.A(net110),
    .B(net124),
    .C(net121),
    .X(_1554_));
 sky130_fd_sc_hd__or2_4 _4338_ (.A(_0831_),
    .B(_1553_),
    .X(_1555_));
 sky130_fd_sc_hd__nand2_8 _4339_ (.A(_1551_),
    .B(_1554_),
    .Y(_1556_));
 sky130_fd_sc_hd__xor2_4 _4340_ (.A(net127),
    .B(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__a31o_2 _4341_ (.A1(net127),
    .A2(_1551_),
    .A3(_1554_),
    .B1(_0835_),
    .X(_1558_));
 sky130_fd_sc_hd__nand2_4 _4342_ (.A(net127),
    .B(_0835_),
    .Y(_1559_));
 sky130_fd_sc_hd__o21ai_4 _4343_ (.A1(_1556_),
    .A2(_1559_),
    .B1(_1558_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2b_4 _4344_ (.A_N(_1560_),
    .B(_1557_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _4345_ (.A(net114),
    .B(net113),
    .Y(_1562_));
 sky130_fd_sc_hd__mux2_8 _4346_ (.A0(_1436_),
    .A1(_1562_),
    .S(_1434_),
    .X(_1563_));
 sky130_fd_sc_hd__nor2_4 _4347_ (.A(net112),
    .B(_1436_),
    .Y(_1564_));
 sky130_fd_sc_hd__or2_4 _4348_ (.A(net112),
    .B(_1436_),
    .X(_1565_));
 sky130_fd_sc_hd__and4_1 _4349_ (.A(net107),
    .B(net106),
    .C(net109),
    .D(net108),
    .X(_1566_));
 sky130_fd_sc_hd__and4_1 _4350_ (.A(net103),
    .B(net102),
    .C(net105),
    .D(net104),
    .X(_1567_));
 sky130_fd_sc_hd__and4_1 _4351_ (.A(net130),
    .B(net129),
    .C(net101),
    .D(net100),
    .X(_1568_));
 sky130_fd_sc_hd__and3_4 _4352_ (.A(_1566_),
    .B(_1567_),
    .C(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__and2_4 _4353_ (.A(net127),
    .B(net128),
    .X(_1570_));
 sky130_fd_sc_hd__and3_4 _4354_ (.A(_1551_),
    .B(_1554_),
    .C(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__a21bo_4 _4355_ (.A1(_1569_),
    .A2(_1571_),
    .B1_N(net111),
    .X(_1572_));
 sky130_fd_sc_hd__nand3b_4 _4356_ (.A_N(net111),
    .B(_1569_),
    .C(_1571_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_2 _4357_ (.A(_1572_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__or3b_4 _4358_ (.A(_1561_),
    .B(_1565_),
    .C_N(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__nand2b_4 _4359_ (.A_N(net99),
    .B(net110),
    .Y(_1576_));
 sky130_fd_sc_hd__nor2_8 _4360_ (.A(_1553_),
    .B(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__or2_4 _4361_ (.A(_1553_),
    .B(_1576_),
    .X(_1578_));
 sky130_fd_sc_hd__nor2_2 _4362_ (.A(net125),
    .B(_1554_),
    .Y(_1579_));
 sky130_fd_sc_hd__and2_2 _4363_ (.A(net125),
    .B(_1554_),
    .X(_1580_));
 sky130_fd_sc_hd__or2_4 _4364_ (.A(_1579_),
    .B(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__o21a_1 _4365_ (.A1(net459),
    .A2(_1580_),
    .B1(_1556_),
    .X(_1582_));
 sky130_fd_sc_hd__o21bai_4 _4366_ (.A1(_1579_),
    .A2(_1580_),
    .B1_N(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__o31a_2 _4367_ (.A1(_1552_),
    .A2(_1575_),
    .A3(_1578_),
    .B1(\wbbd_state[7] ),
    .X(_1584_));
 sky130_fd_sc_hd__or2_4 _4368_ (.A(net112),
    .B(net111),
    .X(_1585_));
 sky130_fd_sc_hd__nand2_4 _4369_ (.A(_1435_),
    .B(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__inv_2 _4370_ (.A(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__and4b_4 _4371_ (.A_N(_1563_),
    .B(_1572_),
    .C(_1573_),
    .D(_1586_),
    .X(_1588_));
 sky130_fd_sc_hd__nand4b_4 _4372_ (.A_N(_1563_),
    .B(_1572_),
    .C(_1573_),
    .D(_1586_),
    .Y(_1589_));
 sky130_fd_sc_hd__nor2_4 _4373_ (.A(_0836_),
    .B(_1581_),
    .Y(_1590_));
 sky130_fd_sc_hd__nand2_4 _4374_ (.A(_1588_),
    .B(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__or2_4 _4375_ (.A(_1561_),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__inv_2 _4376_ (.A(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__nand2_8 _4377_ (.A(net110),
    .B(net99),
    .Y(_1594_));
 sky130_fd_sc_hd__nor2_8 _4378_ (.A(net124),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__or2_4 _4379_ (.A(net124),
    .B(_1594_),
    .X(_1596_));
 sky130_fd_sc_hd__nand2_8 _4380_ (.A(_0833_),
    .B(net121),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_8 _4381_ (.A(net121),
    .B(_1595_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_8 _4382_ (.A(net124),
    .B(_0834_),
    .Y(_1599_));
 sky130_fd_sc_hd__nor2_8 _4383_ (.A(_1594_),
    .B(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__or2_4 _4384_ (.A(_1594_),
    .B(_1599_),
    .X(_1601_));
 sky130_fd_sc_hd__and2_4 _4385_ (.A(_1598_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__nor2_1 _4386_ (.A(_1592_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__or2_4 _4387_ (.A(net128),
    .B(_1557_),
    .X(_1604_));
 sky130_fd_sc_hd__and2_4 _4388_ (.A(_1581_),
    .B(_1582_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_8 _4389_ (.A(_1588_),
    .B(_1605_),
    .Y(_1606_));
 sky130_fd_sc_hd__nor2_8 _4390_ (.A(_1604_),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__or2_4 _4391_ (.A(_1604_),
    .B(_1606_),
    .X(_1608_));
 sky130_fd_sc_hd__or2_4 _4392_ (.A(net124),
    .B(net121),
    .X(_1609_));
 sky130_fd_sc_hd__nor2_8 _4393_ (.A(_1594_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__or2_4 _4394_ (.A(_1594_),
    .B(_1609_),
    .X(_1611_));
 sky130_fd_sc_hd__and4_4 _4395_ (.A(net110),
    .B(net99),
    .C(net124),
    .D(net121),
    .X(_1612_));
 sky130_fd_sc_hd__nand2_8 _4396_ (.A(net99),
    .B(_1554_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_4 _4397_ (.A(_1611_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__inv_2 _4398_ (.A(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__nor2_4 _4399_ (.A(_1591_),
    .B(_1604_),
    .Y(_1616_));
 sky130_fd_sc_hd__or2_4 _4400_ (.A(_1591_),
    .B(_1604_),
    .X(_1617_));
 sky130_fd_sc_hd__nor3_4 _4401_ (.A(_1583_),
    .B(_1589_),
    .C(_1604_),
    .Y(_1618_));
 sky130_fd_sc_hd__or3_4 _4402_ (.A(_1583_),
    .B(_1589_),
    .C(_1604_),
    .X(_1619_));
 sky130_fd_sc_hd__nor2_2 _4403_ (.A(_1613_),
    .B(_1617_),
    .Y(_1620_));
 sky130_fd_sc_hd__nor2_2 _4404_ (.A(_1561_),
    .B(_1606_),
    .Y(_1621_));
 sky130_fd_sc_hd__or2_4 _4405_ (.A(_1561_),
    .B(_1606_),
    .X(_1622_));
 sky130_fd_sc_hd__or3_4 _4406_ (.A(net459),
    .B(_1581_),
    .C(_1589_),
    .X(_1623_));
 sky130_fd_sc_hd__and2_4 _4407_ (.A(_1557_),
    .B(_1560_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_4 _4408_ (.A(_1557_),
    .B(_1560_),
    .Y(_1625_));
 sky130_fd_sc_hd__nor2_4 _4409_ (.A(_1623_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__or4_4 _4410_ (.A(net459),
    .B(_1581_),
    .C(_1589_),
    .D(_1625_),
    .X(_1627_));
 sky130_fd_sc_hd__nor2_1 _4411_ (.A(_1601_),
    .B(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__nor2_2 _4412_ (.A(_1613_),
    .B(_1627_),
    .Y(_1629_));
 sky130_fd_sc_hd__and4_4 _4413_ (.A(net99),
    .B(_1551_),
    .C(_1554_),
    .D(_1570_),
    .X(_1630_));
 sky130_fd_sc_hd__nand2_8 _4414_ (.A(_1569_),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__a31o_2 _4415_ (.A1(_1435_),
    .A2(_1569_),
    .A3(_1630_),
    .B1(_1563_),
    .X(_1632_));
 sky130_fd_sc_hd__xor2_4 _4416_ (.A(net111),
    .B(_1631_),
    .X(_1633_));
 sky130_fd_sc_hd__a21oi_4 _4417_ (.A1(_1585_),
    .A2(_1631_),
    .B1(_1632_),
    .Y(_1634_));
 sky130_fd_sc_hd__xor2_4 _4418_ (.A(net125),
    .B(_1612_),
    .X(_1635_));
 sky130_fd_sc_hd__nand2_2 _4419_ (.A(net459),
    .B(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__and3_2 _4420_ (.A(net127),
    .B(net459),
    .C(net125),
    .X(_1637_));
 sky130_fd_sc_hd__nor2_2 _4421_ (.A(_1552_),
    .B(_1613_),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_2 _4422_ (.A(_1612_),
    .B(_1637_),
    .Y(_1639_));
 sky130_fd_sc_hd__a21o_1 _4423_ (.A1(_1551_),
    .A2(_1612_),
    .B1(net127),
    .X(_1640_));
 sky130_fd_sc_hd__a21oi_2 _4424_ (.A1(_1612_),
    .A2(_1637_),
    .B1(net128),
    .Y(_1641_));
 sky130_fd_sc_hd__a211o_4 _4425_ (.A1(_1639_),
    .A2(_1640_),
    .B1(_1641_),
    .C1(_1630_),
    .X(_1642_));
 sky130_fd_sc_hd__nor2_4 _4426_ (.A(_1636_),
    .B(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_2 _4427_ (.A(_1634_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__and3_2 _4428_ (.A(_1612_),
    .B(_1634_),
    .C(_1643_),
    .X(_1645_));
 sky130_fd_sc_hd__and3_4 _4429_ (.A(_1588_),
    .B(_1605_),
    .C(_1624_),
    .X(_1646_));
 sky130_fd_sc_hd__and4_2 _4430_ (.A(_1588_),
    .B(_1600_),
    .C(_1605_),
    .D(_1624_),
    .X(_1647_));
 sky130_fd_sc_hd__o211a_2 _4431_ (.A1(_1590_),
    .A2(_1605_),
    .B1(_1624_),
    .C1(_1588_),
    .X(_1648_));
 sky130_fd_sc_hd__nor2_4 _4432_ (.A(net110),
    .B(net99),
    .Y(_1649_));
 sky130_fd_sc_hd__or2_4 _4433_ (.A(net110),
    .B(net99),
    .X(_1650_));
 sky130_fd_sc_hd__o211a_4 _4434_ (.A1(net110),
    .A2(net99),
    .B1(net124),
    .C1(net121),
    .X(_1651_));
 sky130_fd_sc_hd__nand2_4 _4435_ (.A(_1551_),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__and3_4 _4436_ (.A(_1551_),
    .B(_1570_),
    .C(_1651_),
    .X(_1653_));
 sky130_fd_sc_hd__nand2_4 _4437_ (.A(_1569_),
    .B(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__xor2_4 _4438_ (.A(net111),
    .B(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__or2_4 _4439_ (.A(_1565_),
    .B(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__xor2_4 _4440_ (.A(net127),
    .B(_1652_),
    .X(_1657_));
 sky130_fd_sc_hd__a31o_2 _4441_ (.A1(net127),
    .A2(_1551_),
    .A3(_1651_),
    .B1(net128),
    .X(_1658_));
 sky130_fd_sc_hd__nand2b_4 _4442_ (.A_N(_1653_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__and2_4 _4443_ (.A(_1657_),
    .B(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__nand2_8 _4444_ (.A(_1657_),
    .B(_1659_),
    .Y(_1661_));
 sky130_fd_sc_hd__o2111a_2 _4445_ (.A1(net110),
    .A2(net99),
    .B1(net124),
    .C1(net121),
    .D1(net125),
    .X(_1662_));
 sky130_fd_sc_hd__xnor2_4 _4446_ (.A(net125),
    .B(_1651_),
    .Y(_1663_));
 sky130_fd_sc_hd__o2bb2a_1 _4447_ (.A1_N(_1551_),
    .A2_N(_1651_),
    .B1(_1662_),
    .B2(net459),
    .X(_1664_));
 sky130_fd_sc_hd__o21ai_2 _4448_ (.A1(net459),
    .A2(_1662_),
    .B1(_1652_),
    .Y(_1665_));
 sky130_fd_sc_hd__nand2_2 _4449_ (.A(_1663_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__or2_2 _4450_ (.A(_1661_),
    .B(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__or2_4 _4451_ (.A(_1656_),
    .B(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__inv_2 _4452_ (.A(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nor2_8 _4453_ (.A(_1599_),
    .B(_1650_),
    .Y(_1670_));
 sky130_fd_sc_hd__or2_4 _4454_ (.A(_1599_),
    .B(_1650_),
    .X(_1671_));
 sky130_fd_sc_hd__nor2_2 _4455_ (.A(_1668_),
    .B(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__or2_4 _4456_ (.A(net124),
    .B(_1576_),
    .X(_1673_));
 sky130_fd_sc_hd__nor2_8 _4457_ (.A(_1576_),
    .B(_1597_),
    .Y(_1674_));
 sky130_fd_sc_hd__or2_4 _4458_ (.A(_1576_),
    .B(_1597_),
    .X(_1675_));
 sky130_fd_sc_hd__nor2_1 _4459_ (.A(_1668_),
    .B(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__or2_4 _4460_ (.A(_1668_),
    .B(_1675_),
    .X(_1677_));
 sky130_fd_sc_hd__nor2_1 _4461_ (.A(net459),
    .B(net125),
    .Y(_1678_));
 sky130_fd_sc_hd__or2_4 _4462_ (.A(net459),
    .B(net125),
    .X(_1679_));
 sky130_fd_sc_hd__or2_4 _4463_ (.A(net127),
    .B(net128),
    .X(_1680_));
 sky130_fd_sc_hd__nor2_8 _4464_ (.A(_1679_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__or2_4 _4465_ (.A(_1679_),
    .B(_1680_),
    .X(_1682_));
 sky130_fd_sc_hd__and2_4 _4466_ (.A(net111),
    .B(_1564_),
    .X(_1683_));
 sky130_fd_sc_hd__nand2_8 _4467_ (.A(net111),
    .B(_1564_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_4 _4468_ (.A(_1681_),
    .B(_1683_),
    .Y(_1685_));
 sky130_fd_sc_hd__nor2_8 _4469_ (.A(net124),
    .B(_1650_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_0833_),
    .B(_1649_),
    .Y(_1687_));
 sky130_fd_sc_hd__or2_4 _4471_ (.A(_1597_),
    .B(_1650_),
    .X(_1688_));
 sky130_fd_sc_hd__nor2_8 _4472_ (.A(net459),
    .B(_1663_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_8 _4473_ (.A(_1656_),
    .B(_1661_),
    .Y(_1690_));
 sky130_fd_sc_hd__nand2_8 _4474_ (.A(_1689_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__nor2_8 _4475_ (.A(_1576_),
    .B(_1599_),
    .Y(_1692_));
 sky130_fd_sc_hd__or2_4 _4476_ (.A(_1576_),
    .B(_1599_),
    .X(_1693_));
 sky130_fd_sc_hd__nor2_1 _4477_ (.A(_1691_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__or3_4 _4478_ (.A(net459),
    .B(_1575_),
    .C(_1581_),
    .X(_1695_));
 sky130_fd_sc_hd__nor2_2 _4479_ (.A(_1611_),
    .B(_1622_),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_4 _4480_ (.A(_1576_),
    .B(_1609_),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_4 _4481_ (.A(_1576_),
    .B(_1609_),
    .X(_1698_));
 sky130_fd_sc_hd__nor2_2 _4482_ (.A(_1668_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_2 _4483_ (.A(_1563_),
    .B(_1586_),
    .Y(_1700_));
 sky130_fd_sc_hd__or3_2 _4484_ (.A(_1563_),
    .B(_1574_),
    .C(_1586_),
    .X(_1701_));
 sky130_fd_sc_hd__clkinv_2 _4485_ (.A(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__and3_2 _4486_ (.A(_0832_),
    .B(_1571_),
    .C(_1588_),
    .X(_1703_));
 sky130_fd_sc_hd__or2_4 _4487_ (.A(_0836_),
    .B(net125),
    .X(_1704_));
 sky130_fd_sc_hd__or2_1 _4488_ (.A(_0836_),
    .B(_1680_),
    .X(_1705_));
 sky130_fd_sc_hd__nor2_8 _4489_ (.A(_1680_),
    .B(_1704_),
    .Y(_1706_));
 sky130_fd_sc_hd__or2_1 _4490_ (.A(_1680_),
    .B(_1704_),
    .X(_1707_));
 sky130_fd_sc_hd__nand2_8 _4491_ (.A(_1683_),
    .B(_1706_),
    .Y(_1708_));
 sky130_fd_sc_hd__or2_4 _4492_ (.A(_1553_),
    .B(_1650_),
    .X(_1709_));
 sky130_fd_sc_hd__nor2_2 _4493_ (.A(_1708_),
    .B(net368),
    .Y(_1710_));
 sky130_fd_sc_hd__nor2_2 _4494_ (.A(_1555_),
    .B(_1708_),
    .Y(_1711_));
 sky130_fd_sc_hd__or3b_4 _4495_ (.A(_1680_),
    .B(net459),
    .C_N(net125),
    .X(_1712_));
 sky130_fd_sc_hd__or2_4 _4496_ (.A(_1684_),
    .B(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__nor2_4 _4497_ (.A(net368),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__nor2_4 _4498_ (.A(_1578_),
    .B(_1713_),
    .Y(_1715_));
 sky130_fd_sc_hd__and3b_4 _4499_ (.A_N(_1583_),
    .B(_1588_),
    .C(_1624_),
    .X(_1716_));
 sky130_fd_sc_hd__and2_2 _4500_ (.A(_1600_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__nor2_2 _4501_ (.A(_1555_),
    .B(_1682_),
    .Y(_1718_));
 sky130_fd_sc_hd__nor2_4 _4502_ (.A(_1578_),
    .B(_1682_),
    .Y(_1719_));
 sky130_fd_sc_hd__inv_2 _4503_ (.A(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__nor2_2 _4504_ (.A(_1682_),
    .B(net368),
    .Y(_1721_));
 sky130_fd_sc_hd__or2_4 _4505_ (.A(_1682_),
    .B(_1709_),
    .X(_1722_));
 sky130_fd_sc_hd__a31o_1 _4506_ (.A1(_1578_),
    .A2(_1693_),
    .A3(_1709_),
    .B1(_1682_),
    .X(_1723_));
 sky130_fd_sc_hd__and3_4 _4507_ (.A(_1588_),
    .B(_1612_),
    .C(_1706_),
    .X(_1724_));
 sky130_fd_sc_hd__and2_2 _4508_ (.A(_1612_),
    .B(_1646_),
    .X(_1725_));
 sky130_fd_sc_hd__nor2_1 _4509_ (.A(_1592_),
    .B(_1611_),
    .Y(_1726_));
 sky130_fd_sc_hd__and2_4 _4510_ (.A(_1663_),
    .B(_1664_),
    .X(_1727_));
 sky130_fd_sc_hd__nand2_4 _4511_ (.A(_1690_),
    .B(_1727_),
    .Y(_1728_));
 sky130_fd_sc_hd__nor2_8 _4512_ (.A(_1604_),
    .B(_1623_),
    .Y(_1729_));
 sky130_fd_sc_hd__or2_4 _4513_ (.A(_1604_),
    .B(_1623_),
    .X(_1730_));
 sky130_fd_sc_hd__nor2_1 _4514_ (.A(_1613_),
    .B(_1619_),
    .Y(_1731_));
 sky130_fd_sc_hd__nor2_2 _4515_ (.A(_1592_),
    .B(_1601_),
    .Y(_1732_));
 sky130_fd_sc_hd__nor2_2 _4516_ (.A(_1601_),
    .B(_1622_),
    .Y(_1733_));
 sky130_fd_sc_hd__and2_1 _4517_ (.A(_1612_),
    .B(_1716_),
    .X(_1734_));
 sky130_fd_sc_hd__nor2_2 _4518_ (.A(_1601_),
    .B(_1730_),
    .Y(_1735_));
 sky130_fd_sc_hd__nor2_1 _4519_ (.A(_1601_),
    .B(_1619_),
    .Y(_1736_));
 sky130_fd_sc_hd__a2111o_4 _4520_ (.A1(_1587_),
    .A2(_1720_),
    .B1(_1723_),
    .C1(_1574_),
    .D1(_1563_),
    .X(_1737_));
 sky130_fd_sc_hd__nor2_1 _4521_ (.A(_1601_),
    .B(_1617_),
    .Y(_1738_));
 sky130_fd_sc_hd__a21oi_2 _4522_ (.A1(_1598_),
    .A2(_1601_),
    .B1(_1617_),
    .Y(_1739_));
 sky130_fd_sc_hd__nor2_4 _4523_ (.A(_1613_),
    .B(_1730_),
    .Y(_1740_));
 sky130_fd_sc_hd__nor2_2 _4524_ (.A(_1608_),
    .B(_1613_),
    .Y(_1741_));
 sky130_fd_sc_hd__or3b_4 _4525_ (.A(_1656_),
    .B(_1661_),
    .C_N(_1727_),
    .X(_1742_));
 sky130_fd_sc_hd__nor2_1 _4526_ (.A(_1693_),
    .B(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__nor2_1 _4527_ (.A(_1578_),
    .B(_1708_),
    .Y(_1744_));
 sky130_fd_sc_hd__and2b_4 _4528_ (.A_N(_1659_),
    .B(_1657_),
    .X(_1745_));
 sky130_fd_sc_hd__and3_4 _4529_ (.A(_1435_),
    .B(_1569_),
    .C(_1653_),
    .X(_1746_));
 sky130_fd_sc_hd__a21boi_4 _4530_ (.A1(_1569_),
    .A2(_1653_),
    .B1_N(_1585_),
    .Y(_1747_));
 sky130_fd_sc_hd__a21bo_1 _4531_ (.A1(_1569_),
    .A2(_1653_),
    .B1_N(_1585_),
    .X(_1748_));
 sky130_fd_sc_hd__nor3_4 _4532_ (.A(_1563_),
    .B(_1746_),
    .C(_1747_),
    .Y(_1749_));
 sky130_fd_sc_hd__or3_4 _4533_ (.A(_1563_),
    .B(_1746_),
    .C(_1747_),
    .X(_1750_));
 sky130_fd_sc_hd__nor2_2 _4534_ (.A(_0836_),
    .B(_1663_),
    .Y(_1751_));
 sky130_fd_sc_hd__and4bb_4 _4535_ (.A_N(_1563_),
    .B_N(_1746_),
    .C(_1748_),
    .D(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__and2_4 _4536_ (.A(_1745_),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__and4bb_4 _4537_ (.A_N(_1563_),
    .B_N(_1746_),
    .C(_1748_),
    .D(_1727_),
    .X(_1754_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(_1727_),
    .B(_1745_),
    .Y(_1755_));
 sky130_fd_sc_hd__and4_1 _4539_ (.A(net110),
    .B(net99),
    .C(_0833_),
    .D(_1648_),
    .X(_1756_));
 sky130_fd_sc_hd__or3b_1 _4540_ (.A(_1645_),
    .B(_1647_),
    .C_N(_1737_),
    .X(_1757_));
 sky130_fd_sc_hd__a21oi_1 _4541_ (.A1(_1598_),
    .A2(_1601_),
    .B1(_1627_),
    .Y(_1758_));
 sky130_fd_sc_hd__or4_1 _4542_ (.A(_1725_),
    .B(_1756_),
    .C(_1757_),
    .D(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__a211o_1 _4543_ (.A1(_1610_),
    .A2(_1626_),
    .B1(_1629_),
    .C1(_1717_),
    .X(_1760_));
 sky130_fd_sc_hd__a211o_1 _4544_ (.A1(_1595_),
    .A2(_1716_),
    .B1(_1759_),
    .C1(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _4545_ (.A1(_1600_),
    .A2(_1607_),
    .B1(_1610_),
    .B2(_1616_),
    .C1(_1620_),
    .X(_1762_));
 sky130_fd_sc_hd__or4_1 _4546_ (.A(_1734_),
    .B(_1739_),
    .C(_1761_),
    .D(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__nor2_1 _4547_ (.A(_1596_),
    .B(_1608_),
    .Y(_1764_));
 sky130_fd_sc_hd__or4_1 _4548_ (.A(_1735_),
    .B(_1741_),
    .C(_1763_),
    .D(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__a211o_1 _4549_ (.A1(_1595_),
    .A2(_1729_),
    .B1(_1740_),
    .C1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__a211o_1 _4550_ (.A1(_1595_),
    .A2(_1618_),
    .B1(_1736_),
    .C1(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__or3_1 _4551_ (.A(_1731_),
    .B(_1732_),
    .C(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__a2111o_1 _4552_ (.A1(_1593_),
    .A2(_1595_),
    .B1(_1724_),
    .C1(_1733_),
    .D1(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__nor3_2 _4553_ (.A(_1561_),
    .B(_1583_),
    .C(_1698_),
    .Y(_1770_));
 sky130_fd_sc_hd__and2_2 _4554_ (.A(_1702_),
    .B(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__a211o_1 _4555_ (.A1(_1595_),
    .A2(_1621_),
    .B1(_1769_),
    .C1(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__or4_1 _4556_ (.A(_1703_),
    .B(_1710_),
    .C(_1744_),
    .D(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__or4_1 _4557_ (.A(_1694_),
    .B(_1715_),
    .C(_1743_),
    .D(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__or3_1 _4558_ (.A(_0834_),
    .B(_1576_),
    .C(_1695_),
    .X(_1775_));
 sky130_fd_sc_hd__or4b_2 _4559_ (.A(_1672_),
    .B(_1714_),
    .C(_1774_),
    .D_N(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__or2_4 _4560_ (.A(_1682_),
    .B(_1688_),
    .X(_1777_));
 sky130_fd_sc_hd__inv_2 _4561_ (.A(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nor2_8 _4562_ (.A(_1684_),
    .B(_1777_),
    .Y(_1779_));
 sky130_fd_sc_hd__o41a_4 _4563_ (.A1(_1676_),
    .A2(_1699_),
    .A3(_1776_),
    .A4(_1779_),
    .B1(_1584_),
    .X(_1780_));
 sky130_fd_sc_hd__nand2_8 _4564_ (.A(_0831_),
    .B(net99),
    .Y(_1781_));
 sky130_fd_sc_hd__nor2_4 _4565_ (.A(_1553_),
    .B(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__or2_4 _4566_ (.A(_1553_),
    .B(_1781_),
    .X(_1783_));
 sky130_fd_sc_hd__o21a_2 _4567_ (.A1(_1668_),
    .A2(_1783_),
    .B1(\wbbd_state[9] ),
    .X(_1784_));
 sky130_fd_sc_hd__nand2_4 _4568_ (.A(_1674_),
    .B(_1729_),
    .Y(_1785_));
 sky130_fd_sc_hd__nor2_4 _4569_ (.A(_1693_),
    .B(_1730_),
    .Y(_1786_));
 sky130_fd_sc_hd__inv_2 _4570_ (.A(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__nor2_4 _4571_ (.A(_1666_),
    .B(_1750_),
    .Y(_1788_));
 sky130_fd_sc_hd__or3_4 _4572_ (.A(_1661_),
    .B(_1666_),
    .C(_1750_),
    .X(_1789_));
 sky130_fd_sc_hd__nor2_2 _4573_ (.A(_1783_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_1577_),
    .B(_1618_),
    .Y(_1792_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(_1601_),
    .B(_1728_),
    .Y(_1793_));
 sky130_fd_sc_hd__nor2_8 _4577_ (.A(_1597_),
    .B(_1781_),
    .Y(_1794_));
 sky130_fd_sc_hd__or2_4 _4578_ (.A(_1597_),
    .B(_1781_),
    .X(_1795_));
 sky130_fd_sc_hd__or2_4 _4579_ (.A(_1685_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a22oi_4 _4580_ (.A1(_1646_),
    .A2(_1692_),
    .B1(_1753_),
    .B2(_1577_),
    .Y(_1797_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_1577_),
    .B(_1646_),
    .Y(_1798_));
 sky130_fd_sc_hd__nor2_1 _4582_ (.A(_1608_),
    .B(_1693_),
    .Y(_1799_));
 sky130_fd_sc_hd__nor2_8 _4583_ (.A(_1599_),
    .B(_1781_),
    .Y(_1800_));
 sky130_fd_sc_hd__or2_4 _4584_ (.A(_1599_),
    .B(_1781_),
    .X(_1801_));
 sky130_fd_sc_hd__nand2_4 _4585_ (.A(_1692_),
    .B(_1716_),
    .Y(_1802_));
 sky130_fd_sc_hd__nand2_4 _4586_ (.A(_1674_),
    .B(_1716_),
    .Y(_1803_));
 sky130_fd_sc_hd__nor2_8 _4587_ (.A(_1609_),
    .B(_1781_),
    .Y(_1804_));
 sky130_fd_sc_hd__or2_4 _4588_ (.A(_1609_),
    .B(_1781_),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_1 _4589_ (.A(_1655_),
    .B(_1700_),
    .Y(_1806_));
 sky130_fd_sc_hd__or2_4 _4590_ (.A(_1667_),
    .B(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__or2_1 _4591_ (.A(net361),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nor2_4 _4592_ (.A(_1682_),
    .B(_1783_),
    .Y(_1809_));
 sky130_fd_sc_hd__nand3_2 _4593_ (.A(_1655_),
    .B(_1700_),
    .C(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__a21oi_4 _4594_ (.A1(_1601_),
    .A2(_1783_),
    .B1(_1682_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _4595_ (.A(_1749_),
    .B(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__nor2_8 _4596_ (.A(_1713_),
    .B(_1783_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor2_4 _4597_ (.A(_1708_),
    .B(_1783_),
    .Y(_1814_));
 sky130_fd_sc_hd__nor2_4 _4598_ (.A(_1627_),
    .B(_1693_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand2_4 _4599_ (.A(_1607_),
    .B(_1674_),
    .Y(_1816_));
 sky130_fd_sc_hd__nor2_2 _4600_ (.A(_1617_),
    .B(_1693_),
    .Y(_1817_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_1691_),
    .B(_1795_),
    .Y(_1818_));
 sky130_fd_sc_hd__nor2_1 _4602_ (.A(_1691_),
    .B(_1783_),
    .Y(_1819_));
 sky130_fd_sc_hd__nor2_4 _4603_ (.A(_1601_),
    .B(_1691_),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(_1668_),
    .B(net361),
    .Y(_1821_));
 sky130_fd_sc_hd__nor2_1 _4605_ (.A(_1598_),
    .B(_1668_),
    .Y(_1822_));
 sky130_fd_sc_hd__or2_2 _4606_ (.A(_1611_),
    .B(_1668_),
    .X(_1823_));
 sky130_fd_sc_hd__inv_2 _4607_ (.A(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__o21ai_1 _4608_ (.A1(_1596_),
    .A2(_1668_),
    .B1(_1796_),
    .Y(_1825_));
 sky130_fd_sc_hd__o21ai_1 _4609_ (.A1(_1577_),
    .A2(_1697_),
    .B1(_1716_),
    .Y(_1826_));
 sky130_fd_sc_hd__o2111ai_4 _4610_ (.A1(_1752_),
    .A2(_1754_),
    .B1(_0832_),
    .C1(_0833_),
    .D1(_1745_),
    .Y(_1827_));
 sky130_fd_sc_hd__o221a_1 _4611_ (.A1(_1789_),
    .A2(_1801_),
    .B1(_1827_),
    .B2(_0831_),
    .C1(_1810_),
    .X(_1828_));
 sky130_fd_sc_hd__and4_4 _4612_ (.A(_1797_),
    .B(_1798_),
    .C(_1812_),
    .D(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__nor2_4 _4613_ (.A(_1627_),
    .B(_1675_),
    .Y(_1830_));
 sky130_fd_sc_hd__or2_1 _4614_ (.A(_1627_),
    .B(_1673_),
    .X(_1831_));
 sky130_fd_sc_hd__and3b_1 _4615_ (.A_N(_1815_),
    .B(_1829_),
    .C(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__o211a_1 _4616_ (.A1(_1578_),
    .A2(_1627_),
    .B1(_1802_),
    .C1(_1803_),
    .X(_1833_));
 sky130_fd_sc_hd__nor2_2 _4617_ (.A(_1617_),
    .B(_1675_),
    .Y(_1834_));
 sky130_fd_sc_hd__a21o_1 _4618_ (.A1(_1673_),
    .A2(_1693_),
    .B1(_1617_),
    .X(_1835_));
 sky130_fd_sc_hd__and4_1 _4619_ (.A(_1826_),
    .B(_1832_),
    .C(_1833_),
    .D(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__o221a_1 _4620_ (.A1(_1578_),
    .A2(_1617_),
    .B1(_1693_),
    .B2(_1608_),
    .C1(_1816_),
    .X(_1837_));
 sky130_fd_sc_hd__o211a_1 _4621_ (.A1(_1608_),
    .A2(_1698_),
    .B1(_1836_),
    .C1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__nand2_1 _4622_ (.A(_1577_),
    .B(_1607_),
    .Y(_1839_));
 sky130_fd_sc_hd__and4_1 _4623_ (.A(_1785_),
    .B(_1787_),
    .C(_1838_),
    .D(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__nand2_1 _4624_ (.A(_1577_),
    .B(_1729_),
    .Y(_1841_));
 sky130_fd_sc_hd__nor2_4 _4625_ (.A(_1619_),
    .B(_1693_),
    .Y(_1842_));
 sky130_fd_sc_hd__inv_2 _4626_ (.A(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__o2111a_2 _4627_ (.A1(_1698_),
    .A2(_1730_),
    .B1(_1840_),
    .C1(_1841_),
    .D1(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__nor2_1 _4628_ (.A(_1619_),
    .B(_1675_),
    .Y(_1845_));
 sky130_fd_sc_hd__nor2_2 _4629_ (.A(_1592_),
    .B(_1693_),
    .Y(_1846_));
 sky130_fd_sc_hd__inv_2 _4630_ (.A(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__o2111a_1 _4631_ (.A1(_1619_),
    .A2(_1673_),
    .B1(_1792_),
    .C1(_1844_),
    .D1(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__nor2_2 _4632_ (.A(_1592_),
    .B(_1675_),
    .Y(_1849_));
 sky130_fd_sc_hd__or2_2 _4633_ (.A(_1578_),
    .B(_1592_),
    .X(_1850_));
 sky130_fd_sc_hd__nand2_1 _4634_ (.A(_1621_),
    .B(_1692_),
    .Y(_1851_));
 sky130_fd_sc_hd__o2111a_1 _4635_ (.A1(_1592_),
    .A2(_1673_),
    .B1(_1848_),
    .C1(_1850_),
    .D1(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__nor2_4 _4636_ (.A(_1622_),
    .B(_1675_),
    .Y(_1853_));
 sky130_fd_sc_hd__o211a_1 _4637_ (.A1(_1622_),
    .A2(_1673_),
    .B1(_1808_),
    .C1(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__or3_4 _4638_ (.A(_1684_),
    .B(_1707_),
    .C(_1783_),
    .X(_1855_));
 sky130_fd_sc_hd__o2111a_1 _4639_ (.A1(_1601_),
    .A2(_1742_),
    .B1(_1791_),
    .C1(_1854_),
    .D1(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__o21ba_1 _4640_ (.A1(_1691_),
    .A2(_1801_),
    .B1_N(_1813_),
    .X(_1857_));
 sky130_fd_sc_hd__o211a_1 _4641_ (.A1(_1742_),
    .A2(_1801_),
    .B1(_1856_),
    .C1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__or4b_2 _4642_ (.A(_1818_),
    .B(_1819_),
    .C(_1820_),
    .D_N(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__or3_4 _4643_ (.A(_1682_),
    .B(_1684_),
    .C(_1795_),
    .X(_1860_));
 sky130_fd_sc_hd__nand2_1 _4644_ (.A(_1823_),
    .B(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__o41a_4 _4645_ (.A1(_1821_),
    .A2(_1822_),
    .A3(_1859_),
    .A4(_1861_),
    .B1(_1784_),
    .X(_1862_));
 sky130_fd_sc_hd__or2_2 _4646_ (.A(_1565_),
    .B(_1633_),
    .X(_1863_));
 sky130_fd_sc_hd__o31a_4 _4647_ (.A1(_0835_),
    .A2(_1639_),
    .A3(_1863_),
    .B1(\wbbd_state[8] ),
    .X(_1864_));
 sky130_fd_sc_hd__nor2_1 _4648_ (.A(_1613_),
    .B(_1708_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_8 _4649_ (.A(_1436_),
    .B(_1585_),
    .Y(_1866_));
 sky130_fd_sc_hd__or2_4 _4650_ (.A(_1436_),
    .B(_1585_),
    .X(_1867_));
 sky130_fd_sc_hd__nor2_8 _4651_ (.A(_1552_),
    .B(_1680_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_8 _4652_ (.A(net367),
    .B(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__nor2_4 _4653_ (.A(net368),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__nor2_8 _4654_ (.A(net127),
    .B(_0835_),
    .Y(_1871_));
 sky130_fd_sc_hd__and3_4 _4655_ (.A(_0836_),
    .B(net125),
    .C(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__and2_4 _4656_ (.A(net367),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_8 _4657_ (.A(net367),
    .B(_1872_),
    .Y(_1874_));
 sky130_fd_sc_hd__a2111o_1 _4658_ (.A1(_1649_),
    .A2(_1873_),
    .B1(_1870_),
    .C1(_1814_),
    .D1(_1813_),
    .X(_1875_));
 sky130_fd_sc_hd__nand2_8 _4659_ (.A(_1706_),
    .B(net367),
    .Y(_1876_));
 sky130_fd_sc_hd__and2_4 _4660_ (.A(_1671_),
    .B(_1688_),
    .X(_1877_));
 sky130_fd_sc_hd__nand2_2 _4661_ (.A(_1671_),
    .B(_1688_),
    .Y(_1878_));
 sky130_fd_sc_hd__nor2_8 _4662_ (.A(_1609_),
    .B(_1650_),
    .Y(_1879_));
 sky130_fd_sc_hd__or2_4 _4663_ (.A(_1609_),
    .B(_1650_),
    .X(_1880_));
 sky130_fd_sc_hd__o22a_1 _4664_ (.A1(net368),
    .A2(_1876_),
    .B1(_1880_),
    .B2(_1869_),
    .X(_1881_));
 sky130_fd_sc_hd__nand2_8 _4665_ (.A(net459),
    .B(_1871_),
    .Y(_1882_));
 sky130_fd_sc_hd__nor2_8 _4666_ (.A(net125),
    .B(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__or2_4 _4667_ (.A(net125),
    .B(_1882_),
    .X(_1884_));
 sky130_fd_sc_hd__nand2_8 _4668_ (.A(net367),
    .B(_1883_),
    .Y(_1885_));
 sky130_fd_sc_hd__a31o_1 _4669_ (.A1(_1688_),
    .A2(net368),
    .A3(_1880_),
    .B1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__o211a_1 _4670_ (.A1(_1876_),
    .A2(_1877_),
    .B1(_1881_),
    .C1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_2 _4671_ (.A(_1613_),
    .B(_1713_),
    .Y(_1888_));
 sky130_fd_sc_hd__and3_1 _4672_ (.A(net99),
    .B(_1718_),
    .C(net367),
    .X(_1889_));
 sky130_fd_sc_hd__nor2_1 _4673_ (.A(_1688_),
    .B(_1869_),
    .Y(_1890_));
 sky130_fd_sc_hd__nor2_4 _4674_ (.A(_1671_),
    .B(_1869_),
    .Y(_1891_));
 sky130_fd_sc_hd__and3_4 _4675_ (.A(_1678_),
    .B(net367),
    .C(_1871_),
    .X(_1892_));
 sky130_fd_sc_hd__or3b_4 _4676_ (.A(_1679_),
    .B(_1867_),
    .C_N(_1871_),
    .X(_1893_));
 sky130_fd_sc_hd__or2_4 _4677_ (.A(_1559_),
    .B(_1867_),
    .X(_1894_));
 sky130_fd_sc_hd__a21oi_2 _4678_ (.A1(_1893_),
    .A2(_1894_),
    .B1(_1650_),
    .Y(_1895_));
 sky130_fd_sc_hd__or3_1 _4679_ (.A(_1890_),
    .B(_1891_),
    .C(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__or4b_1 _4680_ (.A(_1888_),
    .B(_1889_),
    .C(_1896_),
    .D_N(_1887_),
    .X(_1897_));
 sky130_fd_sc_hd__nor2_1 _4681_ (.A(_1688_),
    .B(_1885_),
    .Y(_1898_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(_1688_),
    .B(_1876_),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_2 _4683_ (.A(_1671_),
    .B(_1876_),
    .Y(_1900_));
 sky130_fd_sc_hd__nor2_4 _4684_ (.A(_1679_),
    .B(_1894_),
    .Y(_1901_));
 sky130_fd_sc_hd__or2_4 _4685_ (.A(_1679_),
    .B(_1894_),
    .X(_1902_));
 sky130_fd_sc_hd__nor2_1 _4686_ (.A(_1880_),
    .B(_1893_),
    .Y(_1903_));
 sky130_fd_sc_hd__nor2_4 _4687_ (.A(_1709_),
    .B(_1893_),
    .Y(_1904_));
 sky130_fd_sc_hd__or3_4 _4688_ (.A(_1552_),
    .B(_1559_),
    .C(_1867_),
    .X(_1905_));
 sky130_fd_sc_hd__inv_6 _4689_ (.A(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__or3_4 _4690_ (.A(_1559_),
    .B(_1704_),
    .C(_1867_),
    .X(_1907_));
 sky130_fd_sc_hd__or3b_4 _4691_ (.A(_1894_),
    .B(net459),
    .C_N(net125),
    .X(_1908_));
 sky130_fd_sc_hd__and3_2 _4692_ (.A(_1612_),
    .B(_1681_),
    .C(net367),
    .X(_1909_));
 sky130_fd_sc_hd__and2_4 _4693_ (.A(_1633_),
    .B(_1700_),
    .X(_1910_));
 sky130_fd_sc_hd__nor2_8 _4694_ (.A(_1668_),
    .B(_1801_),
    .Y(_1911_));
 sky130_fd_sc_hd__and2_4 _4695_ (.A(_1551_),
    .B(_1871_),
    .X(_1912_));
 sky130_fd_sc_hd__nand2_8 _4696_ (.A(_1551_),
    .B(_1871_),
    .Y(_1913_));
 sky130_fd_sc_hd__nor2_1 _4697_ (.A(_1688_),
    .B(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__nor2_2 _4698_ (.A(_1671_),
    .B(_1884_),
    .Y(_1915_));
 sky130_fd_sc_hd__o31a_1 _4699_ (.A1(_1811_),
    .A2(_1914_),
    .A3(_1915_),
    .B1(_1634_),
    .X(_1916_));
 sky130_fd_sc_hd__o2bb2a_2 _4700_ (.A1_N(_1639_),
    .A2_N(_1640_),
    .B1(_1641_),
    .B2(_1630_),
    .X(_1917_));
 sky130_fd_sc_hd__a21oi_1 _4701_ (.A1(net125),
    .A2(_1612_),
    .B1(net459),
    .Y(_1918_));
 sky130_fd_sc_hd__or2_1 _4702_ (.A(_1638_),
    .B(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__and3b_2 _4703_ (.A_N(_1635_),
    .B(_1917_),
    .C(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__and3_4 _4704_ (.A(_1610_),
    .B(_1910_),
    .C(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__nor2_2 _4705_ (.A(_1644_),
    .B(_1880_),
    .Y(_1922_));
 sky130_fd_sc_hd__a31o_1 _4706_ (.A1(_1634_),
    .A2(_1670_),
    .A3(_1912_),
    .B1(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__or4bb_4 _4707_ (.A(_1863_),
    .B(net459),
    .C_N(_1635_),
    .D_N(_1917_),
    .X(_1924_));
 sky130_fd_sc_hd__or4_1 _4708_ (.A(_1793_),
    .B(_1865_),
    .C(_1875_),
    .D(_1897_),
    .X(_1925_));
 sky130_fd_sc_hd__a311o_1 _4709_ (.A1(_1570_),
    .A2(_1634_),
    .A3(_1638_),
    .B1(_1921_),
    .C1(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__a21oi_1 _4710_ (.A1(_1598_),
    .A2(_1613_),
    .B1(_1924_),
    .Y(_1927_));
 sky130_fd_sc_hd__and3_1 _4711_ (.A(_1612_),
    .B(_1681_),
    .C(_1910_),
    .X(_1928_));
 sky130_fd_sc_hd__or4_1 _4712_ (.A(_1820_),
    .B(_1825_),
    .C(_1911_),
    .D(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__or4_1 _4713_ (.A(_1916_),
    .B(_1926_),
    .C(_1927_),
    .D(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__or2_1 _4714_ (.A(_1867_),
    .B(_1882_),
    .X(_1931_));
 sky130_fd_sc_hd__a31o_1 _4715_ (.A1(_1670_),
    .A2(net367),
    .A3(_1912_),
    .B1(_1922_),
    .X(_1932_));
 sky130_fd_sc_hd__nor2_1 _4716_ (.A(_1874_),
    .B(_1880_),
    .Y(_1933_));
 sky130_fd_sc_hd__nor2_1 _4717_ (.A(net368),
    .B(_1905_),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_4 _4718_ (.A(_1671_),
    .B(_1907_),
    .Y(_1935_));
 sky130_fd_sc_hd__and3b_4 _4719_ (.A_N(_1559_),
    .B(_1678_),
    .C(_1866_),
    .X(_1936_));
 sky130_fd_sc_hd__o21a_1 _4720_ (.A1(_1923_),
    .A2(_1930_),
    .B1(_1864_),
    .X(_1937_));
 sky130_fd_sc_hd__o21a_4 _4721_ (.A1(_1685_),
    .A2(_1880_),
    .B1(_1532_),
    .X(_1938_));
 sky130_fd_sc_hd__or3b_4 _4722_ (.A(net111),
    .B(_1436_),
    .C_N(net112),
    .X(_1939_));
 sky130_fd_sc_hd__a21o_1 _4723_ (.A1(_1783_),
    .A2(net361),
    .B1(_1885_),
    .X(_1940_));
 sky130_fd_sc_hd__nor3_4 _4724_ (.A(_1712_),
    .B(_1880_),
    .C(_1939_),
    .Y(_1941_));
 sky130_fd_sc_hd__inv_2 _4725_ (.A(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__nor2_1 _4726_ (.A(_1781_),
    .B(_1869_),
    .Y(_1943_));
 sky130_fd_sc_hd__a21oi_1 _4727_ (.A1(_1609_),
    .A2(_1943_),
    .B1(_1941_),
    .Y(_1944_));
 sky130_fd_sc_hd__or2_4 _4728_ (.A(_1552_),
    .B(_1894_),
    .X(_1945_));
 sky130_fd_sc_hd__and3_1 _4729_ (.A(_0833_),
    .B(_0834_),
    .C(_1943_),
    .X(_1946_));
 sky130_fd_sc_hd__o21ba_1 _4730_ (.A1(_1781_),
    .A2(_1902_),
    .B1_N(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__o221a_1 _4731_ (.A1(net361),
    .A2(_1908_),
    .B1(_1945_),
    .B2(_1783_),
    .C1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__o2111a_1 _4732_ (.A1(_1777_),
    .A2(_1939_),
    .B1(_1940_),
    .C1(_1944_),
    .D1(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__o31a_1 _4733_ (.A1(net99),
    .A2(_1553_),
    .A3(_1708_),
    .B1(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__o21a_1 _4734_ (.A1(_1712_),
    .A2(_1880_),
    .B1(_1720_),
    .X(_1951_));
 sky130_fd_sc_hd__or3b_2 _4735_ (.A(net110),
    .B(_0832_),
    .C_N(_1553_),
    .X(_1952_));
 sky130_fd_sc_hd__nor2_2 _4736_ (.A(_1794_),
    .B(_1800_),
    .Y(_1953_));
 sky130_fd_sc_hd__nor2_4 _4737_ (.A(net361),
    .B(_1913_),
    .Y(_1954_));
 sky130_fd_sc_hd__a21oi_1 _4738_ (.A1(_1681_),
    .A2(_1879_),
    .B1(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__o2111a_1 _4739_ (.A1(_1882_),
    .A2(_1953_),
    .B1(_1955_),
    .C1(_1951_),
    .D1(_1722_),
    .X(_1956_));
 sky130_fd_sc_hd__or3_4 _4740_ (.A(_0833_),
    .B(_1781_),
    .C(_1893_),
    .X(_1957_));
 sky130_fd_sc_hd__nand2_4 _4741_ (.A(_1804_),
    .B(_1892_),
    .Y(_1958_));
 sky130_fd_sc_hd__o311a_1 _4742_ (.A1(_0833_),
    .A2(_1781_),
    .A3(_1876_),
    .B1(_1957_),
    .C1(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__a211o_1 _4743_ (.A1(_1705_),
    .A2(_1712_),
    .B1(_1880_),
    .C1(_1684_),
    .X(_1960_));
 sky130_fd_sc_hd__o311a_1 _4744_ (.A1(net99),
    .A2(_1553_),
    .A3(_1713_),
    .B1(_1959_),
    .C1(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__or2_1 _4745_ (.A(_1671_),
    .B(_1713_),
    .X(_1962_));
 sky130_fd_sc_hd__or2_4 _4746_ (.A(_1704_),
    .B(_1894_),
    .X(_1963_));
 sky130_fd_sc_hd__o221a_1 _4747_ (.A1(_1945_),
    .A2(_1952_),
    .B1(_1963_),
    .B2(_1781_),
    .C1(_1962_),
    .X(_1964_));
 sky130_fd_sc_hd__nand2_2 _4748_ (.A(_1794_),
    .B(_1892_),
    .Y(_1965_));
 sky130_fd_sc_hd__or3_4 _4749_ (.A(_1682_),
    .B(_1684_),
    .C(_1693_),
    .X(_1966_));
 sky130_fd_sc_hd__or2_4 _4750_ (.A(_1795_),
    .B(_1876_),
    .X(_1967_));
 sky130_fd_sc_hd__o2111a_1 _4751_ (.A1(_1874_),
    .A2(_1952_),
    .B1(_1965_),
    .C1(_1966_),
    .D1(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__a21o_1 _4752_ (.A1(_1783_),
    .A2(_1953_),
    .B1(_1908_),
    .X(_1969_));
 sky130_fd_sc_hd__and4_1 _4753_ (.A(_1961_),
    .B(_1964_),
    .C(_1968_),
    .D(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__nor2_4 _4754_ (.A(net361),
    .B(_1874_),
    .Y(_1971_));
 sky130_fd_sc_hd__or2_4 _4755_ (.A(net361),
    .B(_1907_),
    .X(_1972_));
 sky130_fd_sc_hd__nor2_1 _4756_ (.A(_1795_),
    .B(_1908_),
    .Y(_1973_));
 sky130_fd_sc_hd__nor2_1 _4757_ (.A(_1795_),
    .B(_1907_),
    .Y(_1974_));
 sky130_fd_sc_hd__and3_1 _4758_ (.A(_1681_),
    .B(net367),
    .C(_1879_),
    .X(_1975_));
 sky130_fd_sc_hd__o211ai_2 _4759_ (.A1(_1867_),
    .A2(_1956_),
    .B1(_1970_),
    .C1(_1950_),
    .Y(_1976_));
 sky130_fd_sc_hd__nor2_1 _4760_ (.A(_1783_),
    .B(_1869_),
    .Y(_1977_));
 sky130_fd_sc_hd__nor2_1 _4761_ (.A(_1795_),
    .B(_1869_),
    .Y(_1978_));
 sky130_fd_sc_hd__a31o_2 _4762_ (.A1(_1745_),
    .A2(_1754_),
    .A3(_1782_),
    .B1(_1976_),
    .X(_1979_));
 sky130_fd_sc_hd__or4_2 _4763_ (.A(_1672_),
    .B(_1676_),
    .C(_1779_),
    .D(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__a211o_4 _4764_ (.A1(_1938_),
    .A2(_1980_),
    .B1(_1534_),
    .C1(_1937_),
    .X(_1981_));
 sky130_fd_sc_hd__o32a_1 _4765_ (.A1(_1780_),
    .A2(_1862_),
    .A3(_1981_),
    .B1(_1535_),
    .B2(\wbbd_addr[0] ),
    .X(_0367_));
 sky130_fd_sc_hd__or2_4 _4766_ (.A(_1696_),
    .B(_1900_),
    .X(_1982_));
 sky130_fd_sc_hd__o22a_1 _4767_ (.A1(_1601_),
    .A2(_1627_),
    .B1(_1880_),
    .B2(_1885_),
    .X(_1983_));
 sky130_fd_sc_hd__a22o_1 _4768_ (.A1(_1610_),
    .A2(_1626_),
    .B1(_1670_),
    .B2(_1873_),
    .X(_1984_));
 sky130_fd_sc_hd__or2_4 _4769_ (.A(_1714_),
    .B(_1813_),
    .X(_1985_));
 sky130_fd_sc_hd__o21a_2 _4770_ (.A1(_1719_),
    .A2(_1809_),
    .B1(_1634_),
    .X(_1986_));
 sky130_fd_sc_hd__nor2_1 _4771_ (.A(_1596_),
    .B(_1924_),
    .Y(_1987_));
 sky130_fd_sc_hd__and3_1 _4772_ (.A(_1610_),
    .B(_1634_),
    .C(_1920_),
    .X(_1988_));
 sky130_fd_sc_hd__or2_4 _4773_ (.A(_1635_),
    .B(_1919_),
    .X(_1989_));
 sky130_fd_sc_hd__or4b_4 _4774_ (.A(_1565_),
    .B(_1989_),
    .C(_1633_),
    .D_N(_1917_),
    .X(_1990_));
 sky130_fd_sc_hd__nor2_1 _4775_ (.A(_1611_),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__nor2_2 _4776_ (.A(_1642_),
    .B(_1989_),
    .Y(_1992_));
 sky130_fd_sc_hd__a21o_1 _4777_ (.A1(_1610_),
    .A2(_1992_),
    .B1(_1915_),
    .X(_1993_));
 sky130_fd_sc_hd__and2_1 _4778_ (.A(_1634_),
    .B(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__o21bai_1 _4779_ (.A1(_1880_),
    .A2(_1907_),
    .B1_N(_1735_),
    .Y(_1995_));
 sky130_fd_sc_hd__a22o_1 _4780_ (.A1(_1610_),
    .A2(_1716_),
    .B1(_1892_),
    .B2(_1670_),
    .X(_1996_));
 sky130_fd_sc_hd__a21o_1 _4781_ (.A1(_1607_),
    .A2(_1610_),
    .B1(_1935_),
    .X(_1997_));
 sky130_fd_sc_hd__o22ai_2 _4782_ (.A1(_1611_),
    .A2(_1730_),
    .B1(_1908_),
    .B2(_1671_),
    .Y(_1998_));
 sky130_fd_sc_hd__or2_1 _4783_ (.A(_1726_),
    .B(_1891_),
    .X(_1999_));
 sky130_fd_sc_hd__o21bai_1 _4784_ (.A1(_1880_),
    .A2(_1908_),
    .B1_N(_1736_),
    .Y(_2000_));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(_1600_),
    .A2(_1607_),
    .B1(_1879_),
    .B2(_1906_),
    .X(_2001_));
 sky130_fd_sc_hd__a22o_1 _4786_ (.A1(_1610_),
    .A2(_1616_),
    .B1(_1670_),
    .B2(_1906_),
    .X(_2002_));
 sky130_fd_sc_hd__or2_4 _4787_ (.A(_1672_),
    .B(_1822_),
    .X(_2003_));
 sky130_fd_sc_hd__a31o_1 _4788_ (.A1(net367),
    .A2(_1868_),
    .A3(_1879_),
    .B1(_1733_),
    .X(_2004_));
 sky130_fd_sc_hd__a22o_1 _4789_ (.A1(_1610_),
    .A2(_1618_),
    .B1(_1670_),
    .B2(_1936_),
    .X(_2005_));
 sky130_fd_sc_hd__a31o_1 _4790_ (.A1(net367),
    .A2(_1879_),
    .A3(_1883_),
    .B1(_1628_),
    .X(_2006_));
 sky130_fd_sc_hd__a31o_1 _4791_ (.A1(_1610_),
    .A2(_1634_),
    .A3(_1920_),
    .B1(_1928_),
    .X(_2007_));
 sky130_fd_sc_hd__o32a_1 _4792_ (.A1(_1611_),
    .A2(_1642_),
    .A3(_1989_),
    .B1(_1884_),
    .B2(_1671_),
    .X(_2008_));
 sky130_fd_sc_hd__inv_2 _4793_ (.A(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__a211o_1 _4794_ (.A1(_1634_),
    .A2(_2009_),
    .B1(_2007_),
    .C1(_1986_),
    .X(_2010_));
 sky130_fd_sc_hd__a31o_1 _4795_ (.A1(_1610_),
    .A2(_1634_),
    .A3(_1643_),
    .B1(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__or4_1 _4796_ (.A(_1647_),
    .B(_1984_),
    .C(_2006_),
    .D(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__or4_1 _4797_ (.A(_1717_),
    .B(_1932_),
    .C(_1933_),
    .D(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__or4_1 _4798_ (.A(_1738_),
    .B(_1903_),
    .C(_2002_),
    .D(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__or4_1 _4799_ (.A(_1995_),
    .B(_1996_),
    .C(_2001_),
    .D(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__or4_1 _4800_ (.A(_1997_),
    .B(_1998_),
    .C(_2000_),
    .D(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__a2111o_1 _4801_ (.A1(_1879_),
    .A2(_1936_),
    .B1(_2005_),
    .C1(_2016_),
    .D1(_1732_),
    .X(_2017_));
 sky130_fd_sc_hd__or4_2 _4802_ (.A(_1982_),
    .B(_1999_),
    .C(_2004_),
    .D(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__a41o_1 _4803_ (.A1(net127),
    .A2(net128),
    .A3(_1634_),
    .A4(_1638_),
    .B1(_1921_),
    .X(_2019_));
 sky130_fd_sc_hd__a41o_1 _4804_ (.A1(net127),
    .A2(net128),
    .A3(_1638_),
    .A4(_1910_),
    .B1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__or4b_1 _4805_ (.A(_1744_),
    .B(_2018_),
    .C(_2020_),
    .D_N(_1855_),
    .X(_2021_));
 sky130_fd_sc_hd__or4_1 _4806_ (.A(_1985_),
    .B(_1987_),
    .C(_1991_),
    .D(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__o41a_4 _4807_ (.A1(_1779_),
    .A2(_1824_),
    .A3(_2003_),
    .A4(_2022_),
    .B1(_1864_),
    .X(_2023_));
 sky130_fd_sc_hd__or2_2 _4808_ (.A(_1672_),
    .B(_1911_),
    .X(_2024_));
 sky130_fd_sc_hd__a21o_1 _4809_ (.A1(_1688_),
    .A2(_1801_),
    .B1(_1963_),
    .X(_2025_));
 sky130_fd_sc_hd__o21ai_1 _4810_ (.A1(_1713_),
    .A2(_1877_),
    .B1(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__a311o_1 _4811_ (.A1(_1800_),
    .A2(net367),
    .A3(_1912_),
    .B1(_1975_),
    .C1(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__or3_4 _4812_ (.A(_1682_),
    .B(_1687_),
    .C(_1939_),
    .X(_2028_));
 sky130_fd_sc_hd__a31o_1 _4813_ (.A1(net121),
    .A2(_1649_),
    .A3(_1873_),
    .B1(_1711_),
    .X(_2029_));
 sky130_fd_sc_hd__or4b_1 _4814_ (.A(_1904_),
    .B(_1971_),
    .C(_2029_),
    .D_N(_2028_),
    .X(_2030_));
 sky130_fd_sc_hd__o21ai_4 _4815_ (.A1(_1709_),
    .A2(_1945_),
    .B1(_1958_),
    .Y(_2031_));
 sky130_fd_sc_hd__o21bai_1 _4816_ (.A1(_1709_),
    .A2(_1876_),
    .B1_N(_1946_),
    .Y(_2032_));
 sky130_fd_sc_hd__or4_1 _4817_ (.A(_2027_),
    .B(_2030_),
    .C(_2031_),
    .D(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__or3_4 _4818_ (.A(net110),
    .B(_1597_),
    .C(_1685_),
    .X(_2034_));
 sky130_fd_sc_hd__or4_1 _4819_ (.A(_0834_),
    .B(_1684_),
    .C(_1687_),
    .D(_1707_),
    .X(_2035_));
 sky130_fd_sc_hd__nand2_1 _4820_ (.A(_2034_),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__or2_2 _4821_ (.A(_1715_),
    .B(_1813_),
    .X(_2037_));
 sky130_fd_sc_hd__a21o_2 _4822_ (.A1(_1804_),
    .A2(_1901_),
    .B1(_1870_),
    .X(_2038_));
 sky130_fd_sc_hd__o22a_1 _4823_ (.A1(net368),
    .A2(_1902_),
    .B1(_1908_),
    .B2(net361),
    .X(_2039_));
 sky130_fd_sc_hd__o22a_1 _4824_ (.A1(net368),
    .A2(_1908_),
    .B1(_1963_),
    .B2(net361),
    .X(_2040_));
 sky130_fd_sc_hd__o221a_1 _4825_ (.A1(net361),
    .A2(_1945_),
    .B1(_1963_),
    .B2(net368),
    .C1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__o2111a_1 _4826_ (.A1(_1777_),
    .A2(_1867_),
    .B1(_1942_),
    .C1(_2039_),
    .D1(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__or4b_1 _4827_ (.A(_2036_),
    .B(_2037_),
    .C(_2038_),
    .D_N(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__a21oi_1 _4828_ (.A1(_1709_),
    .A2(net361),
    .B1(_1884_),
    .Y(_2044_));
 sky130_fd_sc_hd__a211o_1 _4829_ (.A1(_1800_),
    .A2(_1872_),
    .B1(_1914_),
    .C1(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__o31a_1 _4830_ (.A1(_1718_),
    .A2(_1954_),
    .A3(_2045_),
    .B1(net367),
    .X(_2046_));
 sky130_fd_sc_hd__o211a_1 _4831_ (.A1(net459),
    .A2(_1894_),
    .B1(_1945_),
    .C1(_1885_),
    .X(_2047_));
 sky130_fd_sc_hd__and4_1 _4832_ (.A(_1869_),
    .B(_1876_),
    .C(_1893_),
    .D(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__a21oi_1 _4833_ (.A1(_1688_),
    .A2(_1801_),
    .B1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__or4_4 _4834_ (.A(_2033_),
    .B(_2043_),
    .C(_2046_),
    .D(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__o22a_1 _4835_ (.A1(net361),
    .A2(_1869_),
    .B1(_1876_),
    .B2(net368),
    .X(_2051_));
 sky130_fd_sc_hd__a21o_1 _4836_ (.A1(_1688_),
    .A2(_1801_),
    .B1(_1876_),
    .X(_2052_));
 sky130_fd_sc_hd__o22a_1 _4837_ (.A1(_1805_),
    .A2(_1905_),
    .B1(_1907_),
    .B2(net368),
    .X(_2053_));
 sky130_fd_sc_hd__or2_1 _4838_ (.A(_2024_),
    .B(_2050_),
    .X(_2054_));
 sky130_fd_sc_hd__o21a_4 _4839_ (.A1(_1721_),
    .A2(_1809_),
    .B1(_1866_),
    .X(_2055_));
 sky130_fd_sc_hd__or2_2 _4840_ (.A(_1710_),
    .B(_1814_),
    .X(_2056_));
 sky130_fd_sc_hd__nand2b_1 _4841_ (.A_N(_1629_),
    .B(_1802_),
    .Y(_2057_));
 sky130_fd_sc_hd__a22o_2 _4842_ (.A1(_1702_),
    .A2(_1719_),
    .B1(_1770_),
    .B2(_1588_),
    .X(_2058_));
 sky130_fd_sc_hd__nand2_8 _4843_ (.A(_1598_),
    .B(_1698_),
    .Y(_2059_));
 sky130_fd_sc_hd__nor2_1 _4844_ (.A(_1673_),
    .B(_1695_),
    .Y(_2060_));
 sky130_fd_sc_hd__and2_2 _4845_ (.A(_1621_),
    .B(_2059_),
    .X(_2061_));
 sky130_fd_sc_hd__or2_1 _4846_ (.A(_1725_),
    .B(_1815_),
    .X(_2062_));
 sky130_fd_sc_hd__or2_1 _4847_ (.A(_1620_),
    .B(_1799_),
    .X(_2063_));
 sky130_fd_sc_hd__a21o_1 _4848_ (.A1(_1621_),
    .A2(_1692_),
    .B1(_1724_),
    .X(_2064_));
 sky130_fd_sc_hd__or2_1 _4849_ (.A(_1741_),
    .B(_1786_),
    .X(_2065_));
 sky130_fd_sc_hd__or2_1 _4850_ (.A(_1734_),
    .B(_1817_),
    .X(_2066_));
 sky130_fd_sc_hd__nand2b_1 _4851_ (.A_N(_1575_),
    .B(_1605_),
    .Y(_2067_));
 sky130_fd_sc_hd__nor2_1 _4852_ (.A(_1698_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__a2111o_1 _4853_ (.A1(_1646_),
    .A2(_1692_),
    .B1(_2055_),
    .C1(_2058_),
    .D1(_1645_),
    .X(_2069_));
 sky130_fd_sc_hd__a21o_1 _4854_ (.A1(_1626_),
    .A2(_2059_),
    .B1(_2062_),
    .X(_2070_));
 sky130_fd_sc_hd__a211o_1 _4855_ (.A1(_1648_),
    .A2(_2059_),
    .B1(_2069_),
    .C1(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__a2111o_1 _4856_ (.A1(_1716_),
    .A2(_2059_),
    .B1(_2066_),
    .C1(_2071_),
    .D1(_2057_),
    .X(_2072_));
 sky130_fd_sc_hd__a211o_1 _4857_ (.A1(_1607_),
    .A2(_2059_),
    .B1(_1786_),
    .C1(_1741_),
    .X(_2073_));
 sky130_fd_sc_hd__a2111o_1 _4858_ (.A1(_1616_),
    .A2(_2059_),
    .B1(_2063_),
    .C1(_2072_),
    .D1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__a2111o_2 _4859_ (.A1(_1729_),
    .A2(_2059_),
    .B1(_2074_),
    .C1(_1740_),
    .D1(_1842_),
    .X(_2075_));
 sky130_fd_sc_hd__a211o_1 _4860_ (.A1(_1618_),
    .A2(_2059_),
    .B1(_1846_),
    .C1(_1731_),
    .X(_2076_));
 sky130_fd_sc_hd__a2111o_2 _4861_ (.A1(_1593_),
    .A2(_2059_),
    .B1(_2064_),
    .C1(_2075_),
    .D1(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__a31o_1 _4862_ (.A1(_0832_),
    .A2(_1571_),
    .A3(_1702_),
    .B1(_1771_),
    .X(_2078_));
 sky130_fd_sc_hd__or4_1 _4863_ (.A(_1703_),
    .B(_2061_),
    .C(_2077_),
    .D(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__o21ai_1 _4864_ (.A1(_1708_),
    .A2(net368),
    .B1(_1855_),
    .Y(_2080_));
 sky130_fd_sc_hd__or3_1 _4865_ (.A(_2068_),
    .B(_2079_),
    .C(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__or4_1 _4866_ (.A(_1714_),
    .B(_1820_),
    .C(_2060_),
    .D(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__a31o_1 _4867_ (.A1(net110),
    .A2(_0833_),
    .A3(_1669_),
    .B1(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__and3_2 _4868_ (.A(_1674_),
    .B(_1745_),
    .C(_1751_),
    .X(_2084_));
 sky130_fd_sc_hd__o21ai_2 _4869_ (.A1(_1954_),
    .A2(_2084_),
    .B1(_1749_),
    .Y(_2085_));
 sky130_fd_sc_hd__inv_2 _4870_ (.A(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__and2_4 _4871_ (.A(_1601_),
    .B(net368),
    .X(_2087_));
 sky130_fd_sc_hd__nor2_2 _4872_ (.A(_1728_),
    .B(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__a21oi_1 _4873_ (.A1(_1783_),
    .A2(net361),
    .B1(_1807_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_1677_),
    .B(_1796_),
    .Y(_2090_));
 sky130_fd_sc_hd__nor2_4 _4875_ (.A(_1789_),
    .B(_2087_),
    .Y(_2091_));
 sky130_fd_sc_hd__o22a_1 _4876_ (.A1(_1675_),
    .A2(_1755_),
    .B1(net361),
    .B2(_1884_),
    .X(_2092_));
 sky130_fd_sc_hd__or2_2 _4877_ (.A(_1750_),
    .B(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__inv_2 _4878_ (.A(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__o21ai_2 _4879_ (.A1(_1801_),
    .A2(_1876_),
    .B1(_1850_),
    .Y(_2095_));
 sky130_fd_sc_hd__o21ai_1 _4880_ (.A1(_1789_),
    .A2(_1805_),
    .B1(_1810_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(_1803_),
    .B(_1958_),
    .Y(_2097_));
 sky130_fd_sc_hd__a32o_2 _4882_ (.A1(_1800_),
    .A2(net367),
    .A3(_1872_),
    .B1(_1646_),
    .B2(_1577_),
    .X(_2098_));
 sky130_fd_sc_hd__or2_2 _4883_ (.A(_1694_),
    .B(_1820_),
    .X(_2099_));
 sky130_fd_sc_hd__o21ai_4 _4884_ (.A1(net361),
    .A2(_1908_),
    .B1(_1785_),
    .Y(_2100_));
 sky130_fd_sc_hd__o22a_1 _4885_ (.A1(_1578_),
    .A2(_1627_),
    .B1(_1957_),
    .B2(net121),
    .X(_2101_));
 sky130_fd_sc_hd__nor2_1 _4886_ (.A(_1801_),
    .B(_1885_),
    .Y(_2102_));
 sky130_fd_sc_hd__or2_1 _4887_ (.A(_1699_),
    .B(_1821_),
    .X(_2103_));
 sky130_fd_sc_hd__a31o_1 _4888_ (.A1(_1804_),
    .A2(net367),
    .A3(_1868_),
    .B1(_1849_),
    .X(_2104_));
 sky130_fd_sc_hd__o21ai_2 _4889_ (.A1(_1801_),
    .A2(_1869_),
    .B1(_1792_),
    .Y(_2105_));
 sky130_fd_sc_hd__a31o_1 _4890_ (.A1(_1660_),
    .A2(_1754_),
    .A3(_1804_),
    .B1(_1853_),
    .X(_2106_));
 sky130_fd_sc_hd__o22ai_4 _4891_ (.A1(_1578_),
    .A2(_1617_),
    .B1(_1801_),
    .B2(_1907_),
    .Y(_2107_));
 sky130_fd_sc_hd__o21ai_2 _4892_ (.A1(_1801_),
    .A2(_1908_),
    .B1(_1839_),
    .Y(_2108_));
 sky130_fd_sc_hd__nand2_4 _4893_ (.A(_1816_),
    .B(_1972_),
    .Y(_2109_));
 sky130_fd_sc_hd__a21o_1 _4894_ (.A1(_1804_),
    .A2(_1906_),
    .B1(_1834_),
    .X(_2110_));
 sky130_fd_sc_hd__a22o_2 _4895_ (.A1(_1577_),
    .A2(_1626_),
    .B1(_1800_),
    .B2(_1892_),
    .X(_2111_));
 sky130_fd_sc_hd__a22o_4 _4896_ (.A1(_1577_),
    .A2(_1716_),
    .B1(_1800_),
    .B2(_1906_),
    .X(_2112_));
 sky130_fd_sc_hd__nand2_1 _4897_ (.A(_1677_),
    .B(_1860_),
    .Y(_2113_));
 sky130_fd_sc_hd__nor2_1 _4898_ (.A(_1742_),
    .B(net361),
    .Y(_2114_));
 sky130_fd_sc_hd__nor2_1 _4899_ (.A(_1742_),
    .B(_2087_),
    .Y(_2115_));
 sky130_fd_sc_hd__a21oi_1 _4900_ (.A1(_1783_),
    .A2(net361),
    .B1(_1807_),
    .Y(_2116_));
 sky130_fd_sc_hd__a22o_2 _4901_ (.A1(_1577_),
    .A2(_1729_),
    .B1(_1800_),
    .B2(_1936_),
    .X(_2117_));
 sky130_fd_sc_hd__a211o_1 _4902_ (.A1(_1577_),
    .A2(_1753_),
    .B1(_2096_),
    .C1(_2102_),
    .X(_2118_));
 sky130_fd_sc_hd__or4b_1 _4903_ (.A(_2086_),
    .B(_2091_),
    .C(_2098_),
    .D_N(_2093_),
    .X(_2119_));
 sky130_fd_sc_hd__or4_1 _4904_ (.A(_1830_),
    .B(_2111_),
    .C(_2118_),
    .D(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__or4_4 _4905_ (.A(_1971_),
    .B(_2097_),
    .C(_2112_),
    .D(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__or4_1 _4906_ (.A(_2107_),
    .B(_2109_),
    .C(_2110_),
    .D(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__or4_2 _4907_ (.A(_2100_),
    .B(_2108_),
    .C(_2117_),
    .D(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__a2111o_2 _4908_ (.A1(_1804_),
    .A2(_1936_),
    .B1(_2105_),
    .C1(_2123_),
    .D1(_1845_),
    .X(_2124_));
 sky130_fd_sc_hd__or4_1 _4909_ (.A(_2095_),
    .B(_2104_),
    .C(_2106_),
    .D(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__or3_1 _4910_ (.A(_1790_),
    .B(_2116_),
    .C(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__or4_1 _4911_ (.A(_2099_),
    .B(_2114_),
    .C(_2115_),
    .D(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__a21oi_1 _4912_ (.A1(_1795_),
    .A2(net361),
    .B1(_1691_),
    .Y(_2128_));
 sky130_fd_sc_hd__or4_1 _4913_ (.A(_2103_),
    .B(_2113_),
    .C(_2127_),
    .D(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__a221o_1 _4914_ (.A1(_1938_),
    .A2(_2054_),
    .B1(_2129_),
    .B2(_1784_),
    .C1(_1534_),
    .X(_2130_));
 sky130_fd_sc_hd__a21o_2 _4915_ (.A1(_1584_),
    .A2(_2083_),
    .B1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__o22a_1 _4916_ (.A1(\wbbd_addr[1] ),
    .A2(_1535_),
    .B1(_2023_),
    .B2(_2131_),
    .X(_0368_));
 sky130_fd_sc_hd__and3_2 _4917_ (.A(_1823_),
    .B(_1864_),
    .C(_2034_),
    .X(_2132_));
 sky130_fd_sc_hd__nor2_4 _4918_ (.A(_1911_),
    .B(_2003_),
    .Y(_2133_));
 sky130_fd_sc_hd__a311o_2 _4919_ (.A1(net121),
    .A2(_1686_),
    .A3(_1873_),
    .B1(_1984_),
    .C1(_1629_),
    .X(_2134_));
 sky130_fd_sc_hd__or4_1 _4920_ (.A(_1724_),
    .B(_1726_),
    .C(_1890_),
    .D(_1891_),
    .X(_2135_));
 sky130_fd_sc_hd__a22o_1 _4921_ (.A1(_1614_),
    .A2(_1618_),
    .B1(_1878_),
    .B2(_1901_),
    .X(_2136_));
 sky130_fd_sc_hd__or2_2 _4922_ (.A(_1820_),
    .B(_1985_),
    .X(_2137_));
 sky130_fd_sc_hd__a311o_1 _4923_ (.A1(net99),
    .A2(_1718_),
    .A3(_1910_),
    .B1(_1988_),
    .C1(_2091_),
    .X(_2138_));
 sky130_fd_sc_hd__a2bb2o_1 _4924_ (.A1_N(_1908_),
    .A2_N(_1877_),
    .B1(_1729_),
    .B2(_1614_),
    .X(_2139_));
 sky130_fd_sc_hd__a22o_1 _4925_ (.A1(_1614_),
    .A2(_1716_),
    .B1(_1878_),
    .B2(_1892_),
    .X(_2140_));
 sky130_fd_sc_hd__o22a_2 _4926_ (.A1(_1608_),
    .A2(_1615_),
    .B1(_1877_),
    .B2(_1963_),
    .X(_2141_));
 sky130_fd_sc_hd__nor2_2 _4927_ (.A(_1598_),
    .B(_1990_),
    .Y(_2142_));
 sky130_fd_sc_hd__inv_2 _4928_ (.A(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__a31o_1 _4929_ (.A1(_1600_),
    .A2(_1681_),
    .A3(_1910_),
    .B1(_1899_),
    .X(_2144_));
 sky130_fd_sc_hd__and4bb_1 _4930_ (.A_N(_1636_),
    .B_N(_1863_),
    .C(_1917_),
    .D(_1614_),
    .X(_2145_));
 sky130_fd_sc_hd__a211o_1 _4931_ (.A1(_0832_),
    .A2(_1711_),
    .B1(_1814_),
    .C1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__or3_2 _4932_ (.A(_2142_),
    .B(_2144_),
    .C(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__nand2_1 _4933_ (.A(_1634_),
    .B(_1878_),
    .Y(_2148_));
 sky130_fd_sc_hd__o22a_1 _4934_ (.A1(_1615_),
    .A2(_1644_),
    .B1(_1913_),
    .B2(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nand4b_1 _4935_ (.A_N(_1982_),
    .B(_2133_),
    .C(_2149_),
    .D(_1966_),
    .Y(_2150_));
 sky130_fd_sc_hd__or3_2 _4936_ (.A(_1928_),
    .B(_1988_),
    .C(_2091_),
    .X(_2151_));
 sky130_fd_sc_hd__or4_1 _4937_ (.A(_1725_),
    .B(_1898_),
    .C(_1994_),
    .D(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__a21oi_1 _4938_ (.A1(_1671_),
    .A2(_1688_),
    .B1(_1907_),
    .Y(_2153_));
 sky130_fd_sc_hd__a211o_2 _4939_ (.A1(_1607_),
    .A2(_1610_),
    .B1(_1741_),
    .C1(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__or4_1 _4940_ (.A(_2137_),
    .B(_2147_),
    .C(_2152_),
    .D(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__or4_1 _4941_ (.A(_2135_),
    .B(_2136_),
    .C(_2150_),
    .D(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__a311o_1 _4942_ (.A1(net121),
    .A2(_1686_),
    .A3(_1906_),
    .B1(_2002_),
    .C1(_1620_),
    .X(_2157_));
 sky130_fd_sc_hd__a21oi_1 _4943_ (.A1(_1671_),
    .A2(_1688_),
    .B1(_1908_),
    .Y(_2158_));
 sky130_fd_sc_hd__a211o_1 _4944_ (.A1(_1610_),
    .A2(_1729_),
    .B1(_1740_),
    .C1(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__or4_1 _4945_ (.A(_2134_),
    .B(_2140_),
    .C(_2157_),
    .D(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__or2_1 _4946_ (.A(_2156_),
    .B(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__nand2_8 _4947_ (.A(_1698_),
    .B(_1783_),
    .Y(_2162_));
 sky130_fd_sc_hd__a31o_2 _4948_ (.A1(_1745_),
    .A2(_1754_),
    .A3(_2162_),
    .B1(_2094_),
    .X(_2163_));
 sky130_fd_sc_hd__and4_1 _4949_ (.A(_1689_),
    .B(_1745_),
    .C(_1749_),
    .D(_2162_),
    .X(_2164_));
 sky130_fd_sc_hd__or3_4 _4950_ (.A(_1830_),
    .B(_1971_),
    .C(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__a31o_1 _4951_ (.A1(_1745_),
    .A2(_1752_),
    .A3(_2162_),
    .B1(_2086_),
    .X(_2166_));
 sky130_fd_sc_hd__a31o_2 _4952_ (.A1(_1689_),
    .A2(_1690_),
    .A3(_1800_),
    .B1(_2099_),
    .X(_2167_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(_1728_),
    .B(_1795_),
    .Y(_2168_));
 sky130_fd_sc_hd__o22ai_4 _4954_ (.A1(_1622_),
    .A2(_1698_),
    .B1(_1801_),
    .B2(_1807_),
    .Y(_2169_));
 sky130_fd_sc_hd__a311o_1 _4955_ (.A1(_1660_),
    .A2(_1754_),
    .A3(_1804_),
    .B1(_1853_),
    .C1(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__and3_2 _4956_ (.A(_1690_),
    .B(_1751_),
    .C(_1804_),
    .X(_2171_));
 sky130_fd_sc_hd__or3_1 _4957_ (.A(_1814_),
    .B(_2088_),
    .C(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__nor2_4 _4958_ (.A(net128),
    .B(_1657_),
    .Y(_2173_));
 sky130_fd_sc_hd__and2_4 _4959_ (.A(_2162_),
    .B(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__a31o_4 _4960_ (.A1(_1689_),
    .A2(_1749_),
    .A3(_2174_),
    .B1(_2100_),
    .X(_2175_));
 sky130_fd_sc_hd__a21oi_1 _4961_ (.A1(_1693_),
    .A2(_1801_),
    .B1(_1789_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_2 _4962_ (.A(_2096_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__inv_2 _4963_ (.A(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__a21o_2 _4964_ (.A1(_1752_),
    .A2(_2174_),
    .B1(_2110_),
    .X(_2179_));
 sky130_fd_sc_hd__nor2_1 _4965_ (.A(_1742_),
    .B(_1795_),
    .Y(_2180_));
 sky130_fd_sc_hd__a31o_1 _4966_ (.A1(_1660_),
    .A2(_1752_),
    .A3(_2162_),
    .B1(_2104_),
    .X(_2181_));
 sky130_fd_sc_hd__a221o_2 _4967_ (.A1(_1804_),
    .A2(_1936_),
    .B1(_2174_),
    .B2(_1788_),
    .C1(_1845_),
    .X(_2182_));
 sky130_fd_sc_hd__a31o_4 _4968_ (.A1(_1754_),
    .A2(_2162_),
    .A3(_2173_),
    .B1(_2109_),
    .X(_2183_));
 sky130_fd_sc_hd__a31o_2 _4969_ (.A1(_1745_),
    .A2(_1788_),
    .A3(_2162_),
    .B1(_2097_),
    .X(_2184_));
 sky130_fd_sc_hd__or3b_2 _4970_ (.A(_1750_),
    .B(_1755_),
    .C_N(_2162_),
    .X(_2185_));
 sky130_fd_sc_hd__or3b_2 _4971_ (.A(_2094_),
    .B(_2177_),
    .C_N(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__a2111o_4 _4972_ (.A1(_1753_),
    .A2(_2162_),
    .B1(_2165_),
    .C1(_2186_),
    .D1(_2086_),
    .X(_2187_));
 sky130_fd_sc_hd__or4_1 _4973_ (.A(_2179_),
    .B(_2183_),
    .C(_2184_),
    .D(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__or4_1 _4974_ (.A(_2175_),
    .B(_2181_),
    .C(_2182_),
    .D(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__or3_1 _4975_ (.A(_2106_),
    .B(_2169_),
    .C(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__or4b_1 _4976_ (.A(_2115_),
    .B(_2190_),
    .C(_2171_),
    .D_N(_1855_),
    .X(_2191_));
 sky130_fd_sc_hd__or4_2 _4977_ (.A(_2003_),
    .B(_2167_),
    .C(_2180_),
    .D(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__or3b_2 _4978_ (.A(_1824_),
    .B(_2103_),
    .C_N(_1784_),
    .X(_2193_));
 sky130_fd_sc_hd__o21ba_4 _4979_ (.A1(_2113_),
    .A2(_2192_),
    .B1_N(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__or4b_4 _4980_ (.A(_1699_),
    .B(_1779_),
    .C(_1824_),
    .D_N(_1584_),
    .X(_2195_));
 sky130_fd_sc_hd__nand2_2 _4981_ (.A(_1677_),
    .B(_2133_),
    .Y(_2196_));
 sky130_fd_sc_hd__a311o_2 _4982_ (.A1(_1681_),
    .A2(_1692_),
    .A3(_1702_),
    .B1(_2061_),
    .C1(_1696_),
    .X(_2197_));
 sky130_fd_sc_hd__or2_2 _4983_ (.A(_1714_),
    .B(_2099_),
    .X(_2198_));
 sky130_fd_sc_hd__a21oi_4 _4984_ (.A1(_1601_),
    .A2(_1693_),
    .B1(_1682_),
    .Y(_2199_));
 sky130_fd_sc_hd__a21oi_1 _4985_ (.A1(_1588_),
    .A2(_2199_),
    .B1(_2058_),
    .Y(_2200_));
 sky130_fd_sc_hd__and3_4 _4986_ (.A(_1578_),
    .B(_1596_),
    .C(_1698_),
    .X(_2201_));
 sky130_fd_sc_hd__or3_4 _4987_ (.A(_1577_),
    .B(_1595_),
    .C(_1697_),
    .X(_2202_));
 sky130_fd_sc_hd__nor2_2 _4988_ (.A(_1608_),
    .B(_2201_),
    .Y(_2203_));
 sky130_fd_sc_hd__nor2_1 _4989_ (.A(_1675_),
    .B(_2067_),
    .Y(_2204_));
 sky130_fd_sc_hd__nor2_1 _4990_ (.A(_1730_),
    .B(_2201_),
    .Y(_2205_));
 sky130_fd_sc_hd__a211o_2 _4991_ (.A1(net110),
    .A2(net99),
    .B1(_1553_),
    .C1(_1708_),
    .X(_2206_));
 sky130_fd_sc_hd__nand2_1 _4992_ (.A(_1590_),
    .B(_1697_),
    .Y(_2207_));
 sky130_fd_sc_hd__o21ai_2 _4993_ (.A1(_1575_),
    .A2(_2207_),
    .B1(_2206_),
    .Y(_2208_));
 sky130_fd_sc_hd__o31a_1 _4994_ (.A1(_1616_),
    .A2(_1648_),
    .A3(_1716_),
    .B1(_2202_),
    .X(_2209_));
 sky130_fd_sc_hd__nor2_2 _4995_ (.A(_1619_),
    .B(_2201_),
    .Y(_2210_));
 sky130_fd_sc_hd__nor2_1 _4996_ (.A(_1592_),
    .B(_2201_),
    .Y(_2211_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_1627_),
    .B(_2201_),
    .Y(_2212_));
 sky130_fd_sc_hd__or2_2 _4998_ (.A(_2205_),
    .B(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__or4b_1 _4999_ (.A(_2204_),
    .B(_2208_),
    .C(_2210_),
    .D_N(_2200_),
    .X(_2214_));
 sky130_fd_sc_hd__or4_1 _5000_ (.A(_2196_),
    .B(_2203_),
    .C(_2209_),
    .D(_2211_),
    .X(_2215_));
 sky130_fd_sc_hd__or4_1 _5001_ (.A(_2198_),
    .B(_2213_),
    .C(_2214_),
    .D(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__o21ba_1 _5002_ (.A1(_2197_),
    .A2(_2216_),
    .B1_N(_2195_),
    .X(_2217_));
 sky130_fd_sc_hd__and3_1 _5003_ (.A(_1677_),
    .B(_1938_),
    .C(_2034_),
    .X(_2218_));
 sky130_fd_sc_hd__and2_1 _5004_ (.A(_1683_),
    .B(_2199_),
    .X(_2219_));
 sky130_fd_sc_hd__and3_4 _5005_ (.A(_1687_),
    .B(_1795_),
    .C(_1801_),
    .X(_2220_));
 sky130_fd_sc_hd__a21o_1 _5006_ (.A1(_1869_),
    .A2(_1945_),
    .B1(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__o32a_1 _5007_ (.A1(net126),
    .A2(_1894_),
    .A3(_2220_),
    .B1(_1671_),
    .B2(_1708_),
    .X(_2222_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_2221_),
    .B(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__a31o_1 _5009_ (.A1(_1683_),
    .A2(_1686_),
    .A3(_1868_),
    .B1(_1711_),
    .X(_2224_));
 sky130_fd_sc_hd__o22a_1 _5010_ (.A1(_1688_),
    .A2(_1876_),
    .B1(_1939_),
    .B2(_1722_),
    .X(_2225_));
 sky130_fd_sc_hd__o211a_1 _5011_ (.A1(_1801_),
    .A2(_1876_),
    .B1(_1967_),
    .C1(_2225_),
    .X(_2226_));
 sky130_fd_sc_hd__or3b_1 _5012_ (.A(_2223_),
    .B(_2224_),
    .C_N(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__or2_4 _5013_ (.A(_1714_),
    .B(_2037_),
    .X(_2228_));
 sky130_fd_sc_hd__a211o_2 _5014_ (.A1(_1778_),
    .A2(net367),
    .B1(_1941_),
    .C1(_2055_),
    .X(_2229_));
 sky130_fd_sc_hd__a41o_1 _5015_ (.A1(_1874_),
    .A2(_1893_),
    .A3(_1931_),
    .A4(_1963_),
    .B1(_2220_),
    .X(_2230_));
 sky130_fd_sc_hd__or4b_2 _5016_ (.A(_2227_),
    .B(_2228_),
    .C(_2229_),
    .D_N(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__nor2_1 _5017_ (.A(_1902_),
    .B(_2220_),
    .Y(_2232_));
 sky130_fd_sc_hd__or3_1 _5018_ (.A(_2024_),
    .B(_2219_),
    .C(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__a21o_1 _5019_ (.A1(_2218_),
    .A2(_2233_),
    .B1(_1534_),
    .X(_2234_));
 sky130_fd_sc_hd__a211o_4 _5020_ (.A1(_2132_),
    .A2(_2161_),
    .B1(_2217_),
    .C1(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__o22a_1 _5021_ (.A1(\wbbd_addr[2] ),
    .A2(_1535_),
    .B1(_2194_),
    .B2(_2235_),
    .X(_0369_));
 sky130_fd_sc_hd__or4_2 _5022_ (.A(_1739_),
    .B(_1903_),
    .C(_1934_),
    .D(_2140_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5023_ (.A(_1598_),
    .B(_1644_),
    .Y(_2237_));
 sky130_fd_sc_hd__or4_2 _5024_ (.A(_1889_),
    .B(_1986_),
    .C(_2138_),
    .D(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__o22a_2 _5025_ (.A1(net368),
    .A2(_1908_),
    .B1(_1963_),
    .B2(_1880_),
    .X(_2239_));
 sky130_fd_sc_hd__o211ai_4 _5026_ (.A1(_1602_),
    .A2(_1730_),
    .B1(_2141_),
    .C1(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__a2111o_1 _5027_ (.A1(_1879_),
    .A2(_1901_),
    .B1(_2136_),
    .C1(_1870_),
    .D1(_1603_),
    .X(_2241_));
 sky130_fd_sc_hd__or4_1 _5028_ (.A(_2236_),
    .B(_2238_),
    .C(_2240_),
    .D(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__a2111o_1 _5029_ (.A1(_1630_),
    .A2(_1910_),
    .B1(_1921_),
    .C1(_1982_),
    .D1(_2144_),
    .X(_2243_));
 sky130_fd_sc_hd__a311o_1 _5030_ (.A1(_1600_),
    .A2(_1681_),
    .A3(_1683_),
    .B1(_2088_),
    .C1(_2142_),
    .X(_2244_));
 sky130_fd_sc_hd__or3b_1 _5031_ (.A(_1594_),
    .B(_1924_),
    .C_N(_1599_),
    .X(_2245_));
 sky130_fd_sc_hd__o221a_1 _5032_ (.A1(_1598_),
    .A2(_1627_),
    .B1(net368),
    .B2(_1874_),
    .C1(_1983_),
    .X(_2246_));
 sky130_fd_sc_hd__or4b_2 _5033_ (.A(_1725_),
    .B(_1898_),
    .C(_1994_),
    .D_N(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__or4b_1 _5034_ (.A(_2137_),
    .B(_2244_),
    .C(_2247_),
    .D_N(_2245_),
    .X(_2248_));
 sky130_fd_sc_hd__or4_1 _5035_ (.A(_1909_),
    .B(_1986_),
    .C(_2151_),
    .D(_2237_),
    .X(_2249_));
 sky130_fd_sc_hd__or3_1 _5036_ (.A(_2242_),
    .B(_2243_),
    .C(_2248_),
    .X(_2250_));
 sky130_fd_sc_hd__or3b_4 _5037_ (.A(_2024_),
    .B(_2219_),
    .C_N(_2218_),
    .X(_2251_));
 sky130_fd_sc_hd__nor2_1 _5038_ (.A(_1534_),
    .B(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__a2bb2o_1 _5039_ (.A1_N(_1893_),
    .A2_N(_2220_),
    .B1(_1906_),
    .B2(_1670_),
    .X(_2253_));
 sky130_fd_sc_hd__a211o_1 _5040_ (.A1(_1782_),
    .A2(_1906_),
    .B1(_2031_),
    .C1(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__a21o_1 _5041_ (.A1(net124),
    .A2(_1649_),
    .B1(_1782_),
    .X(_2255_));
 sky130_fd_sc_hd__o21ai_2 _5042_ (.A1(_1671_),
    .A2(_1913_),
    .B1(_1951_),
    .Y(_2256_));
 sky130_fd_sc_hd__o31a_2 _5043_ (.A1(net110),
    .A2(_1553_),
    .A3(_1908_),
    .B1(_1972_),
    .X(_2257_));
 sky130_fd_sc_hd__o221ai_2 _5044_ (.A1(_1671_),
    .A2(_1908_),
    .B1(_2220_),
    .B2(_1907_),
    .C1(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__a211o_1 _5045_ (.A1(net367),
    .A2(_2256_),
    .B1(_2229_),
    .C1(_1909_),
    .X(_2259_));
 sky130_fd_sc_hd__or3_1 _5046_ (.A(_2056_),
    .B(_2258_),
    .C(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__or4_1 _5047_ (.A(_1891_),
    .B(_1977_),
    .C(_2038_),
    .D(_2232_),
    .X(_2261_));
 sky130_fd_sc_hd__or2_1 _5048_ (.A(_2254_),
    .B(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__a22o_1 _5049_ (.A1(_1804_),
    .A2(_1883_),
    .B1(_2255_),
    .B2(_1872_),
    .X(_2263_));
 sky130_fd_sc_hd__or3_1 _5050_ (.A(net125),
    .B(_1931_),
    .C(_2220_),
    .X(_2264_));
 sky130_fd_sc_hd__a21bo_1 _5051_ (.A1(net367),
    .A2(_2263_),
    .B1_N(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__a211o_1 _5052_ (.A1(_1877_),
    .A2(_1880_),
    .B1(_1684_),
    .C1(_1712_),
    .X(_2266_));
 sky130_fd_sc_hd__o221ai_2 _5053_ (.A1(_1671_),
    .A2(_1708_),
    .B1(net368),
    .B2(_1685_),
    .C1(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__o2111ai_4 _5054_ (.A1(_1722_),
    .A2(_1939_),
    .B1(_1967_),
    .C1(_2028_),
    .D1(_2052_),
    .Y(_2268_));
 sky130_fd_sc_hd__or2_1 _5055_ (.A(_2228_),
    .B(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__or4_1 _5056_ (.A(_2262_),
    .B(_2265_),
    .C(_2267_),
    .D(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__or2_2 _5057_ (.A(_2260_),
    .B(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__a22o_1 _5058_ (.A1(\wbbd_addr[3] ),
    .A2(_1534_),
    .B1(_2252_),
    .B2(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__a41o_1 _5059_ (.A1(_1966_),
    .A2(_2132_),
    .A3(_2133_),
    .A4(_2250_),
    .B1(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__or2_4 _5060_ (.A(_2090_),
    .B(_2193_),
    .X(_2274_));
 sky130_fd_sc_hd__nor2_1 _5061_ (.A(_2003_),
    .B(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__or3_1 _5062_ (.A(_1795_),
    .B(_1867_),
    .C(_1913_),
    .X(_2276_));
 sky130_fd_sc_hd__o2111a_2 _5063_ (.A1(_1722_),
    .A2(_1867_),
    .B1(_2178_),
    .C1(_2276_),
    .D1(_1812_),
    .X(_2277_));
 sky130_fd_sc_hd__a311o_4 _5064_ (.A1(_1749_),
    .A2(_1794_),
    .A3(_1872_),
    .B1(_2098_),
    .C1(_1815_),
    .X(_2278_));
 sky130_fd_sc_hd__nor2_4 _5065_ (.A(_2163_),
    .B(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_2 _5066_ (.A(_2277_),
    .B(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__a211o_1 _5067_ (.A1(net124),
    .A2(_0834_),
    .B1(_1691_),
    .C1(_1781_),
    .X(_2281_));
 sky130_fd_sc_hd__or3b_1 _5068_ (.A(_1911_),
    .B(_2168_),
    .C_N(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__or4_1 _5069_ (.A(_1819_),
    .B(_1911_),
    .C(_2128_),
    .D(_2180_),
    .X(_2283_));
 sky130_fd_sc_hd__a21oi_1 _5070_ (.A1(_1693_),
    .A2(_1801_),
    .B1(_1742_),
    .Y(_2284_));
 sky130_fd_sc_hd__or4_4 _5071_ (.A(_1786_),
    .B(_1973_),
    .C(_2108_),
    .D(_2183_),
    .X(_2285_));
 sky130_fd_sc_hd__a2111o_1 _5072_ (.A1(_1794_),
    .A2(_1906_),
    .B1(_2112_),
    .C1(_2184_),
    .D1(_1817_),
    .X(_2286_));
 sky130_fd_sc_hd__or4_2 _5073_ (.A(_1846_),
    .B(_1978_),
    .C(_2105_),
    .D(_2182_),
    .X(_2287_));
 sky130_fd_sc_hd__or4_1 _5074_ (.A(_2280_),
    .B(_2285_),
    .C(_2286_),
    .D(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__or4_1 _5075_ (.A(_2106_),
    .B(_2116_),
    .C(_2169_),
    .D(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__or4_2 _5076_ (.A(_2167_),
    .B(_2283_),
    .C(_2284_),
    .D(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__nor2_1 _5077_ (.A(_2195_),
    .B(_2196_),
    .Y(_2291_));
 sky130_fd_sc_hd__or3_1 _5078_ (.A(_1732_),
    .B(_1849_),
    .C(_2210_),
    .X(_2292_));
 sky130_fd_sc_hd__or3_1 _5079_ (.A(_1731_),
    .B(_1846_),
    .C(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__a2111o_1 _5080_ (.A1(_1716_),
    .A2(_2202_),
    .B1(_2066_),
    .C1(_1834_),
    .D1(_1738_),
    .X(_2294_));
 sky130_fd_sc_hd__or4b_2 _5081_ (.A(_1735_),
    .B(_2065_),
    .C(_2203_),
    .D_N(_1785_),
    .X(_2295_));
 sky130_fd_sc_hd__a2111o_2 _5082_ (.A1(_1646_),
    .A2(_2202_),
    .B1(_1830_),
    .C1(_1628_),
    .D1(_2062_),
    .X(_2296_));
 sky130_fd_sc_hd__or4_2 _5083_ (.A(_2293_),
    .B(_2294_),
    .C(_2295_),
    .D(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__or2_1 _5084_ (.A(_2078_),
    .B(_2197_),
    .X(_2298_));
 sky130_fd_sc_hd__o21ai_1 _5085_ (.A1(_1578_),
    .A2(_1695_),
    .B1(_1966_),
    .Y(_2299_));
 sky130_fd_sc_hd__or2_1 _5086_ (.A(_2060_),
    .B(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__or4_4 _5087_ (.A(_1719_),
    .B(_1721_),
    .C(_1809_),
    .D(_2084_),
    .X(_2301_));
 sky130_fd_sc_hd__a21bo_1 _5088_ (.A1(_1588_),
    .A2(_2301_),
    .B1_N(_2200_),
    .X(_2302_));
 sky130_fd_sc_hd__a21oi_1 _5089_ (.A1(_1601_),
    .A2(_1693_),
    .B1(_1728_),
    .Y(_2303_));
 sky130_fd_sc_hd__or4_1 _5090_ (.A(_2204_),
    .B(_2300_),
    .C(_2302_),
    .D(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__or3_1 _5091_ (.A(_2198_),
    .B(_2298_),
    .C(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__o21a_1 _5092_ (.A1(_2297_),
    .A2(_2305_),
    .B1(_2291_),
    .X(_2306_));
 sky130_fd_sc_hd__a211o_1 _5093_ (.A1(_2275_),
    .A2(_2290_),
    .B1(_2306_),
    .C1(_2273_),
    .X(_0370_));
 sky130_fd_sc_hd__a311o_1 _5094_ (.A1(net121),
    .A2(_1595_),
    .A3(_1716_),
    .B1(_1717_),
    .C1(_1933_),
    .X(_2307_));
 sky130_fd_sc_hd__or4_2 _5095_ (.A(_1904_),
    .B(_2134_),
    .C(_2247_),
    .D(_2307_),
    .X(_2308_));
 sky130_fd_sc_hd__o22a_1 _5096_ (.A1(net368),
    .A2(_1902_),
    .B1(_1908_),
    .B2(_1880_),
    .X(_2309_));
 sky130_fd_sc_hd__o21ai_1 _5097_ (.A1(_1602_),
    .A2(_1619_),
    .B1(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__or3_2 _5098_ (.A(_2139_),
    .B(_2240_),
    .C(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__or3_1 _5099_ (.A(_1888_),
    .B(_1991_),
    .C(_2088_),
    .X(_2312_));
 sky130_fd_sc_hd__a211o_1 _5100_ (.A1(_1630_),
    .A2(_1634_),
    .B1(_1715_),
    .C1(_2146_),
    .X(_2313_));
 sky130_fd_sc_hd__or4_1 _5101_ (.A(_2243_),
    .B(_2311_),
    .C(_2312_),
    .D(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__and4b_1 _5102_ (.A_N(_2219_),
    .B(_2245_),
    .C(_2132_),
    .D(_2133_),
    .X(_2315_));
 sky130_fd_sc_hd__o211a_1 _5103_ (.A1(_2308_),
    .A2(_2314_),
    .B1(_2315_),
    .C1(_2143_),
    .X(_2316_));
 sky130_fd_sc_hd__a21oi_1 _5104_ (.A1(net361),
    .A2(_2220_),
    .B1(_1874_),
    .Y(_2317_));
 sky130_fd_sc_hd__or3_2 _5105_ (.A(_1975_),
    .B(_2224_),
    .C(_2268_),
    .X(_2318_));
 sky130_fd_sc_hd__a21oi_1 _5106_ (.A1(_1671_),
    .A2(_1783_),
    .B1(_1902_),
    .Y(_2319_));
 sky130_fd_sc_hd__o21ai_2 _5107_ (.A1(_1908_),
    .A2(_2220_),
    .B1(_2039_),
    .Y(_2320_));
 sky130_fd_sc_hd__or3_2 _5108_ (.A(_2258_),
    .B(_2319_),
    .C(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__a211o_1 _5109_ (.A1(_1892_),
    .A2(_2255_),
    .B1(_2265_),
    .C1(_2317_),
    .X(_2322_));
 sky130_fd_sc_hd__a311o_1 _5110_ (.A1(_1683_),
    .A2(_1686_),
    .A3(_1706_),
    .B1(_1888_),
    .C1(_2056_),
    .X(_2323_));
 sky130_fd_sc_hd__or4_4 _5111_ (.A(_2318_),
    .B(_2321_),
    .C(_2322_),
    .D(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__a221o_4 _5112_ (.A1(\wbbd_addr[4] ),
    .A2(_1534_),
    .B1(_2252_),
    .B2(_2324_),
    .C1(_2316_),
    .X(_2325_));
 sky130_fd_sc_hd__a21oi_1 _5113_ (.A1(_1601_),
    .A2(_1675_),
    .B1(_1619_),
    .Y(_2326_));
 sky130_fd_sc_hd__or4_1 _5114_ (.A(_1740_),
    .B(_1842_),
    .C(_2205_),
    .D(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__or2_2 _5115_ (.A(_2295_),
    .B(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__or4b_1 _5116_ (.A(_1717_),
    .B(_2057_),
    .C(_2212_),
    .D_N(_1803_),
    .X(_2329_));
 sky130_fd_sc_hd__or2_2 _5117_ (.A(_2296_),
    .B(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__or4_1 _5118_ (.A(_1703_),
    .B(_2068_),
    .C(_2208_),
    .D(_2303_),
    .X(_2331_));
 sky130_fd_sc_hd__or3_1 _5119_ (.A(_1715_),
    .B(_2298_),
    .C(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__or4_2 _5120_ (.A(_1813_),
    .B(_2328_),
    .C(_2330_),
    .D(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__or4_1 _5121_ (.A(_2195_),
    .B(_2196_),
    .C(_2204_),
    .D(_2300_),
    .X(_2334_));
 sky130_fd_sc_hd__a31o_2 _5122_ (.A1(_1693_),
    .A2(_1801_),
    .A3(net361),
    .B1(_1728_),
    .X(_2335_));
 sky130_fd_sc_hd__and4b_4 _5123_ (.A_N(_2165_),
    .B(_1965_),
    .C(_1802_),
    .D(_2101_),
    .X(_2336_));
 sky130_fd_sc_hd__nand4b_4 _5124_ (.A_N(_1985_),
    .B(_2279_),
    .C(_2335_),
    .D(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__a2111o_1 _5125_ (.A1(_1794_),
    .A2(_1936_),
    .B1(_2117_),
    .C1(_2175_),
    .D1(_1842_),
    .X(_2338_));
 sky130_fd_sc_hd__nor2_1 _5126_ (.A(_2285_),
    .B(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__inv_2 _5127_ (.A(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__or4_4 _5128_ (.A(_1790_),
    .B(_2089_),
    .C(_2170_),
    .D(_2172_),
    .X(_2341_));
 sky130_fd_sc_hd__or4bb_1 _5129_ (.A(_2111_),
    .B(_2165_),
    .C_N(_1802_),
    .D_N(_1965_),
    .X(_2342_));
 sky130_fd_sc_hd__or4b_4 _5130_ (.A(_2094_),
    .B(_2278_),
    .C(_2342_),
    .D_N(_2185_),
    .X(_2343_));
 sky130_fd_sc_hd__nor3_2 _5131_ (.A(_2337_),
    .B(_2340_),
    .C(_2341_),
    .Y(_2344_));
 sky130_fd_sc_hd__or3_1 _5132_ (.A(_2003_),
    .B(_2274_),
    .C(_2282_),
    .X(_2345_));
 sky130_fd_sc_hd__nor2_2 _5133_ (.A(_2274_),
    .B(_2344_),
    .Y(_2346_));
 sky130_fd_sc_hd__a211o_4 _5134_ (.A1(_2291_),
    .A2(_2333_),
    .B1(_2346_),
    .C1(_2325_),
    .X(_0371_));
 sky130_fd_sc_hd__or4_2 _5135_ (.A(_1813_),
    .B(_2198_),
    .C(_2332_),
    .D(_2334_),
    .X(_2347_));
 sky130_fd_sc_hd__or4_1 _5136_ (.A(_1733_),
    .B(_1853_),
    .C(_2064_),
    .D(_2211_),
    .X(_2348_));
 sky130_fd_sc_hd__or3_1 _5137_ (.A(_2293_),
    .B(_2328_),
    .C(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__o21ai_1 _5138_ (.A1(_1674_),
    .A2(_1692_),
    .B1(_1646_),
    .Y(_2350_));
 sky130_fd_sc_hd__o31a_1 _5139_ (.A1(_1591_),
    .A2(_1625_),
    .A3(_2201_),
    .B1(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__or4b_4 _5140_ (.A(_1645_),
    .B(_1647_),
    .C(_2302_),
    .D_N(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__o21ba_1 _5141_ (.A1(_2349_),
    .A2(_2352_),
    .B1_N(_2347_),
    .X(_2353_));
 sky130_fd_sc_hd__or3b_2 _5142_ (.A(_1985_),
    .B(_2167_),
    .C_N(_2335_),
    .X(_2354_));
 sky130_fd_sc_hd__nor3_2 _5143_ (.A(_2341_),
    .B(_2345_),
    .C(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_1851_),
    .B(_1967_),
    .Y(_2356_));
 sky130_fd_sc_hd__or4_2 _5145_ (.A(_2095_),
    .B(_2181_),
    .C(_2287_),
    .D(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__nor2_1 _5146_ (.A(_2340_),
    .B(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__nor3_1 _5147_ (.A(_1750_),
    .B(_1884_),
    .C(_1953_),
    .Y(_2359_));
 sky130_fd_sc_hd__or4bb_4 _5148_ (.A(_2166_),
    .B(_2359_),
    .C_N(_2277_),
    .D_N(_1797_),
    .X(_2360_));
 sky130_fd_sc_hd__o31a_1 _5149_ (.A1(_2340_),
    .A2(_2357_),
    .A3(_2360_),
    .B1(_2355_),
    .X(_2361_));
 sky130_fd_sc_hd__o221a_1 _5150_ (.A1(_1783_),
    .A2(_1876_),
    .B1(_2220_),
    .B2(_1869_),
    .C1(_2051_),
    .X(_2362_));
 sky130_fd_sc_hd__or3b_1 _5151_ (.A(_1900_),
    .B(_2261_),
    .C_N(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__a2bb2o_1 _5152_ (.A1_N(_1913_),
    .A2_N(_2220_),
    .B1(_2255_),
    .B2(_1883_),
    .X(_2364_));
 sky130_fd_sc_hd__o21a_1 _5153_ (.A1(_1954_),
    .A2(_2364_),
    .B1(net367),
    .X(_2365_));
 sky130_fd_sc_hd__or2_1 _5154_ (.A(_2259_),
    .B(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__or3_2 _5155_ (.A(_2321_),
    .B(_2363_),
    .C(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__or3_1 _5156_ (.A(_1534_),
    .B(_2228_),
    .C(_2323_),
    .X(_2368_));
 sky130_fd_sc_hd__or3_4 _5157_ (.A(_2267_),
    .B(_2318_),
    .C(_2368_),
    .X(_2369_));
 sky130_fd_sc_hd__nor2_2 _5158_ (.A(_2251_),
    .B(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__a2111o_1 _5159_ (.A1(_1630_),
    .A2(_1634_),
    .B1(_1820_),
    .C1(_1921_),
    .D1(_2228_),
    .X(_2371_));
 sky130_fd_sc_hd__a211oi_2 _5160_ (.A1(_1630_),
    .A2(_1910_),
    .B1(_1982_),
    .C1(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__and4bb_2 _5161_ (.A_N(_2147_),
    .B_N(_2312_),
    .C(_2315_),
    .D(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__o21ai_1 _5162_ (.A1(_1602_),
    .A2(_1622_),
    .B1(_1881_),
    .Y(_2374_));
 sky130_fd_sc_hd__or3_1 _5163_ (.A(_2135_),
    .B(_2241_),
    .C(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__nand2_1 _5164_ (.A(_1602_),
    .B(net368),
    .Y(_2376_));
 sky130_fd_sc_hd__and3_1 _5165_ (.A(_1634_),
    .B(_1992_),
    .C(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__or4b_2 _5166_ (.A(_1922_),
    .B(_2377_),
    .C(_2249_),
    .D_N(_2149_),
    .X(_2378_));
 sky130_fd_sc_hd__o31a_1 _5167_ (.A1(_2311_),
    .A2(_2375_),
    .A3(_2378_),
    .B1(_2373_),
    .X(_2379_));
 sky130_fd_sc_hd__a221o_2 _5168_ (.A1(\wbbd_addr[5] ),
    .A2(_1534_),
    .B1(_2367_),
    .B2(_2370_),
    .C1(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__or3_2 _5169_ (.A(_2353_),
    .B(_2361_),
    .C(_2380_),
    .X(_0372_));
 sky130_fd_sc_hd__o221a_1 _5170_ (.A1(_1601_),
    .A2(_1608_),
    .B1(_1617_),
    .B2(_2201_),
    .C1(_1816_),
    .X(_2381_));
 sky130_fd_sc_hd__or4b_1 _5171_ (.A(_2063_),
    .B(_2294_),
    .C(_2352_),
    .D_N(_2381_),
    .X(_2382_));
 sky130_fd_sc_hd__nor2_1 _5172_ (.A(_2347_),
    .B(_2349_),
    .Y(_2383_));
 sky130_fd_sc_hd__o21a_1 _5173_ (.A1(_2330_),
    .A2(_2382_),
    .B1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__or4_2 _5174_ (.A(_1799_),
    .B(_1974_),
    .C(_2107_),
    .D(_2179_),
    .X(_2385_));
 sky130_fd_sc_hd__or4_1 _5175_ (.A(_2286_),
    .B(_2343_),
    .C(_2360_),
    .D(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__o221a_1 _5176_ (.A1(_1783_),
    .A2(_1907_),
    .B1(_2220_),
    .B2(_1905_),
    .C1(_2053_),
    .X(_2387_));
 sky130_fd_sc_hd__nand2b_1 _5177_ (.A_N(_2254_),
    .B(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__or4_4 _5178_ (.A(_1935_),
    .B(_2322_),
    .C(_2366_),
    .D(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__o22a_1 _5179_ (.A1(_1598_),
    .A2(_1608_),
    .B1(net368),
    .B2(_1907_),
    .X(_2390_));
 sky130_fd_sc_hd__or4b_2 _5180_ (.A(_2001_),
    .B(_2157_),
    .C(_2236_),
    .D_N(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__o31a_1 _5181_ (.A1(_2308_),
    .A2(_2378_),
    .A3(_2391_),
    .B1(_2373_),
    .X(_2392_));
 sky130_fd_sc_hd__a221o_4 _5182_ (.A1(\wbbd_addr[6] ),
    .A2(_1534_),
    .B1(_2370_),
    .B2(_2389_),
    .C1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__a31o_1 _5183_ (.A1(_2355_),
    .A2(_2358_),
    .A3(_2386_),
    .B1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__or2_2 _5184_ (.A(_2384_),
    .B(_2394_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_4 _5185_ (.A(_1075_),
    .B(net362),
    .Y(_2395_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(net399),
    .A1(net1647),
    .S(_2395_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(net394),
    .A1(net1363),
    .S(_2395_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _5188_ (.A0(net388),
    .A1(net1458),
    .S(_2395_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(net383),
    .A1(net1432),
    .S(_2395_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(net379),
    .A1(net1195),
    .S(_2395_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _5191_ (.A(_1254_),
    .B(net362),
    .Y(_2396_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(net399),
    .A1(net1669),
    .S(_2396_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net394),
    .A1(net1389),
    .S(_2396_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_4 _5194_ (.A(_1099_),
    .B(net362),
    .Y(_2397_));
 sky130_fd_sc_hd__mux2_1 _5195_ (.A0(net399),
    .A1(net1658),
    .S(_2397_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _5196_ (.A0(net394),
    .A1(net1394),
    .S(_2397_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(net388),
    .A1(net1522),
    .S(_2397_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _5198_ (.A0(net383),
    .A1(net1476),
    .S(_2397_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(net379),
    .A1(net1285),
    .S(_2397_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_8 _5200_ (.A(_1008_),
    .B(net362),
    .Y(_2398_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(net399),
    .A1(net1651),
    .S(_2398_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(net394),
    .A1(net1381),
    .S(_2398_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _5203_ (.A0(net388),
    .A1(net1488),
    .S(_2398_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _5204_ (.A0(net383),
    .A1(net1442),
    .S(_2398_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _5205_ (.A0(net379),
    .A1(net1249),
    .S(_2398_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _5206_ (.A0(net375),
    .A1(net1067),
    .S(_2398_),
    .X(_0399_));
 sky130_fd_sc_hd__and2_4 _5207_ (.A(_0922_),
    .B(net363),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(net1633),
    .A1(net400),
    .S(_2399_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(net834),
    .A1(net396),
    .S(_2399_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(net1503),
    .A1(net388),
    .S(_2399_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(net1365),
    .A1(net383),
    .S(_2399_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(net928),
    .A1(net379),
    .S(_2399_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _5213_ (.A0(net1076),
    .A1(net375),
    .S(_2399_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(net1141),
    .A1(net372),
    .S(_2399_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(net879),
    .A1(net369),
    .S(_2399_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_1311_),
    .B(net363),
    .Y(_2400_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(net401),
    .A1(net1546),
    .S(_2400_),
    .X(_0408_));
 sky130_fd_sc_hd__and2_4 _5218_ (.A(net640),
    .B(net363),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(net1535),
    .A1(net401),
    .S(_2401_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(net815),
    .A1(net396),
    .S(_2401_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(net1142),
    .A1(net389),
    .S(_2401_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(net1723),
    .A1(net598),
    .S(_2401_),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(_1310_),
    .B(net362),
    .Y(_2402_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(net399),
    .A1(net1662),
    .S(_2402_),
    .X(_0413_));
 sky130_fd_sc_hd__or3_1 _5225_ (.A(net356),
    .B(net587),
    .C(net399),
    .X(_2403_));
 sky130_fd_sc_hd__o211a_1 _5226_ (.A1(net1595),
    .A2(_1314_),
    .B1(net363),
    .C1(_2403_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_8 _5227_ (.A(_0972_),
    .B(net363),
    .Y(_2404_));
 sky130_fd_sc_hd__mux2_1 _5228_ (.A0(net631),
    .A1(net1718),
    .S(_2404_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _5229_ (.A0(net598),
    .A1(net1707),
    .S(_2404_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(net389),
    .A1(net1166),
    .S(_2404_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(net375),
    .A1(net1037),
    .S(_2404_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(net372),
    .A1(net1134),
    .S(_2404_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(net396),
    .A1(serial_bb_enable),
    .S(_2404_),
    .X(_0420_));
 sky130_fd_sc_hd__or3_4 _5234_ (.A(net569),
    .B(_0971_),
    .C(net399),
    .X(_2405_));
 sky130_fd_sc_hd__o211a_1 _5235_ (.A1(net1660),
    .A2(_0972_),
    .B1(net363),
    .C1(_2405_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(_1312_),
    .B(net365),
    .Y(_2406_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(net403),
    .A1(net1645),
    .S(_2406_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_2 _5238_ (.A(_1191_),
    .B(net366),
    .Y(_2407_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(net392),
    .A1(net1187),
    .S(_2407_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(net398),
    .A1(net887),
    .S(_2407_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(net402),
    .A1(net1529),
    .S(_2407_),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_1253_),
    .B(net362),
    .Y(_2408_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(net399),
    .A1(net1686),
    .S(_2408_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(net394),
    .A1(net1398),
    .S(_2408_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_8 _5245_ (.A(_1006_),
    .B(net366),
    .Y(_2409_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(net400),
    .A1(net1671),
    .S(_2409_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(net395),
    .A1(net953),
    .S(_2409_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(net392),
    .A1(net1003),
    .S(_2409_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(net383),
    .A1(net1472),
    .S(_2409_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _5250_ (.A0(net381),
    .A1(net1342),
    .S(_2409_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(net540),
    .A1(net557),
    .S(_2409_),
    .X(_0433_));
 sky130_fd_sc_hd__or4_4 _5252_ (.A(net359),
    .B(_0932_),
    .C(net412),
    .D(net677),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(net399),
    .A1(net1425),
    .S(net678),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net394),
    .A1(net1374),
    .S(net678),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(net389),
    .A1(net1149),
    .S(net678),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net598),
    .A1(net1700),
    .S(net678),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(net647),
    .A1(net755),
    .S(net678),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(net375),
    .A1(net1162),
    .S(net678),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _5259_ (.A0(net671),
    .A1(net708),
    .S(net678),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(net369),
    .A1(net891),
    .S(net678),
    .X(_0441_));
 sky130_fd_sc_hd__and2_4 _5261_ (.A(net570),
    .B(net363),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(net1538),
    .A1(net401),
    .S(_2411_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(net857),
    .A1(net396),
    .S(_2411_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(net1218),
    .A1(net389),
    .S(_2411_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(net660),
    .A1(net598),
    .S(_2411_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(net739),
    .A1(net631),
    .S(_2411_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _5267_ (.A0(net1111),
    .A1(net375),
    .S(_2411_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _5268_ (.A0(net1168),
    .A1(net372),
    .S(_2411_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(net1709),
    .A1(net476),
    .S(_2411_),
    .X(_0449_));
 sky130_fd_sc_hd__nand2_8 _5270_ (.A(net490),
    .B(net366),
    .Y(_2412_));
 sky130_fd_sc_hd__mux2_1 _5271_ (.A0(net402),
    .A1(net1447),
    .S(net491),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net397),
    .A1(net854),
    .S(net491),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _5273_ (.A0(net390),
    .A1(net1547),
    .S(net491),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(net533),
    .A1(net633),
    .S(net491),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(net381),
    .A1(net1082),
    .S(net491),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(net540),
    .A1(net1717),
    .S(net491),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(net671),
    .A1(net718),
    .S(net491),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(net476),
    .A1(net1704),
    .S(net491),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_8 _5279_ (.A(_0963_),
    .B(net365),
    .Y(_2413_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(net402),
    .A1(net1436),
    .S(_2413_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net397),
    .A1(net1018),
    .S(_2413_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(net390),
    .A1(net1622),
    .S(_2413_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net533),
    .A1(net802),
    .S(_2413_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net381),
    .A1(net1317),
    .S(_2413_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(net540),
    .A1(net726),
    .S(_2413_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _5286_ (.A0(net373),
    .A1(net1229),
    .S(_2413_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(net370),
    .A1(net981),
    .S(_2413_),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_8 _5288_ (.A(_0942_),
    .B(net366),
    .Y(_2414_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(net403),
    .A1(net1575),
    .S(_2414_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(net397),
    .A1(net1049),
    .S(_2414_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net390),
    .A1(net1610),
    .S(_2414_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(net386),
    .A1(net1098),
    .S(_2414_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net381),
    .A1(net1305),
    .S(_2414_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(net376),
    .A1(net855),
    .S(_2414_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(net373),
    .A1(net1061),
    .S(_2414_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(net370),
    .A1(net839),
    .S(_2414_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_8 _5297_ (.A(_0936_),
    .B(net366),
    .Y(_2415_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(net402),
    .A1(net1491),
    .S(_2415_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net397),
    .A1(net969),
    .S(_2415_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net391),
    .A1(net1407),
    .S(_2415_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(net386),
    .A1(net1034),
    .S(_2415_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net381),
    .A1(net1313),
    .S(_2415_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net376),
    .A1(net930),
    .S(_2415_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(net373),
    .A1(net1001),
    .S(_2415_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net370),
    .A1(net828),
    .S(_2415_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_8 _5306_ (.A(_0941_),
    .B(net365),
    .Y(_2416_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net402),
    .A1(net1427),
    .S(_2416_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net397),
    .A1(net1089),
    .S(_2416_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net390),
    .A1(net1598),
    .S(_2416_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net386),
    .A1(net1045),
    .S(_2416_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(net381),
    .A1(net1289),
    .S(_2416_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net376),
    .A1(net1014),
    .S(_2416_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(net373),
    .A1(net1121),
    .S(_2416_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(net370),
    .A1(net848),
    .S(_2416_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_8 _5315_ (.A(_0927_),
    .B(net365),
    .Y(_2417_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(net402),
    .A1(net1537),
    .S(_2417_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _5317_ (.A0(net397),
    .A1(net1203),
    .S(_2417_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _5318_ (.A0(net390),
    .A1(net1618),
    .S(_2417_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(net386),
    .A1(net1240),
    .S(_2417_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(net382),
    .A1(net906),
    .S(_2417_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net376),
    .A1(net1043),
    .S(_2417_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _5322_ (.A0(net373),
    .A1(net1199),
    .S(_2417_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(net370),
    .A1(net991),
    .S(_2417_),
    .X(_0497_));
 sky130_fd_sc_hd__nand2_8 _5324_ (.A(_0914_),
    .B(net366),
    .Y(_2418_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net402),
    .A1(net1487),
    .S(_2418_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(net398),
    .A1(net777),
    .S(_2418_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5327_ (.A0(net392),
    .A1(net973),
    .S(_2418_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(net386),
    .A1(net1035),
    .S(_2418_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(net381),
    .A1(net1197),
    .S(_2418_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(net376),
    .A1(net911),
    .S(_2418_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net373),
    .A1(net1047),
    .S(_2418_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(net370),
    .A1(net809),
    .S(_2418_),
    .X(_0505_));
 sky130_fd_sc_hd__and2_4 _5333_ (.A(_0913_),
    .B(net366),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net1422),
    .A1(net402),
    .S(_2419_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net1021),
    .A1(net397),
    .S(_2419_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(net1614),
    .A1(net390),
    .S(_2419_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net1125),
    .A1(net386),
    .S(_2419_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(net1299),
    .A1(net381),
    .S(_2419_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _5339_ (.A0(net866),
    .A1(net376),
    .S(_2419_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _5340_ (.A0(net1051),
    .A1(net373),
    .S(_2419_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(net799),
    .A1(net370),
    .S(_2419_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_8 _5342_ (.A(_0895_),
    .B(net366),
    .Y(_2420_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net402),
    .A1(net1424),
    .S(_2420_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(net398),
    .A1(net773),
    .S(_2420_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(net390),
    .A1(net1585),
    .S(_2420_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net386),
    .A1(net1053),
    .S(_2420_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(net382),
    .A1(net763),
    .S(_2420_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(net376),
    .A1(net836),
    .S(_2420_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(net373),
    .A1(net1007),
    .S(_2420_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net370),
    .A1(net797),
    .S(_2420_),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_8 _5351_ (.A(_0945_),
    .B(net366),
    .Y(_2421_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(net402),
    .A1(net1504),
    .S(_2421_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(net398),
    .A1(net794),
    .S(_2421_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(net390),
    .A1(net1608),
    .S(_2421_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(net386),
    .A1(net1255),
    .S(_2421_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net381),
    .A1(net1307),
    .S(_2421_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(net376),
    .A1(net904),
    .S(_2421_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(net373),
    .A1(net1086),
    .S(_2421_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(net370),
    .A1(net1055),
    .S(_2421_),
    .X(_0529_));
 sky130_fd_sc_hd__nand2_8 _5360_ (.A(_0951_),
    .B(net363),
    .Y(_2422_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net401),
    .A1(net1534),
    .S(_2422_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(net396),
    .A1(net841),
    .S(_2422_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net505),
    .A1(net1724),
    .S(_2422_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(net598),
    .A1(net724),
    .S(_2422_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net647),
    .A1(net699),
    .S(_2422_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(net375),
    .A1(net1172),
    .S(_2422_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net372),
    .A1(net1084),
    .S(_2422_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net369),
    .A1(net860),
    .S(_2422_),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_8 _5369_ (.A(_0964_),
    .B(net366),
    .Y(_2423_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(net402),
    .A1(net1486),
    .S(_2423_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net397),
    .A1(net1157),
    .S(_2423_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(net390),
    .A1(net1643),
    .S(_2423_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net386),
    .A1(net1258),
    .S(_2423_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(net381),
    .A1(net1311),
    .S(_2423_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(net376),
    .A1(net1024),
    .S(_2423_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(net373),
    .A1(net1214),
    .S(_2423_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(net370),
    .A1(net961),
    .S(_2423_),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_8 _5378_ (.A(_0894_),
    .B(net366),
    .Y(_2424_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net1347),
    .A1(\gpio_configure[13][0] ),
    .S(net563),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(net398),
    .A1(net844),
    .S(net563),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net390),
    .A1(net1649),
    .S(net563),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(net533),
    .A1(net757),
    .S(net563),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net382),
    .A1(net895),
    .S(net563),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _5384_ (.A0(net376),
    .A1(net1041),
    .S(net563),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(net671),
    .A1(net753),
    .S(net563),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _5386_ (.A0(net476),
    .A1(net1714),
    .S(net563),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_8 _5387_ (.A(_0916_),
    .B(net366),
    .Y(_2425_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(net402),
    .A1(net1483),
    .S(_2425_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(net398),
    .A1(net795),
    .S(_2425_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(net392),
    .A1(net1012),
    .S(_2425_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(net386),
    .A1(net1092),
    .S(_2425_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(net382),
    .A1(net745),
    .S(_2425_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(net376),
    .A1(net938),
    .S(_2425_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _5394_ (.A0(net373),
    .A1(net1208),
    .S(_2425_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(net370),
    .A1(net830),
    .S(_2425_),
    .X(_0561_));
 sky130_fd_sc_hd__and2_4 _5396_ (.A(_0958_),
    .B(net366),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(net1380),
    .A1(net1347),
    .S(_2426_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(net970),
    .A1(net397),
    .S(_2426_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(net1246),
    .A1(net392),
    .S(_2426_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(net1244),
    .A1(net386),
    .S(_2426_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(net940),
    .A1(net382),
    .S(_2426_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(net649),
    .A1(net540),
    .S(_2426_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(net722),
    .A1(net671),
    .S(_2426_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(net955),
    .A1(net370),
    .S(_2426_),
    .X(_0569_));
 sky130_fd_sc_hd__and2_4 _5405_ (.A(_0961_),
    .B(net366),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(net1437),
    .A1(net402),
    .S(_2427_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(net776),
    .A1(net398),
    .S(_2427_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(net977),
    .A1(net392),
    .S(_2427_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(net1079),
    .A1(net386),
    .S(_2427_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(net741),
    .A1(net382),
    .S(_2427_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(net871),
    .A1(net376),
    .S(_2427_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _5412_ (.A0(net1022),
    .A1(net373),
    .S(_2427_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(net832),
    .A1(net370),
    .S(_2427_),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_8 _5414_ (.A(net579),
    .B(net363),
    .Y(_2428_));
 sky130_fd_sc_hd__mux2_1 _5415_ (.A0(net401),
    .A1(net1557),
    .S(_2428_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(net396),
    .A1(net859),
    .S(_2428_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(net389),
    .A1(net1138),
    .S(_2428_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(net598),
    .A1(net682),
    .S(_2428_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(net647),
    .A1(net692),
    .S(_2428_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _5420_ (.A0(net540),
    .A1(net1715),
    .S(_2428_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(net372),
    .A1(net1236),
    .S(_2428_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _5422_ (.A0(net369),
    .A1(net944),
    .S(_2428_),
    .X(_0585_));
 sky130_fd_sc_hd__nand2_8 _5423_ (.A(_0938_),
    .B(net509),
    .Y(_2429_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(net401),
    .A1(net1533),
    .S(net510),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(net396),
    .A1(net813),
    .S(net510),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(net505),
    .A1(net1722),
    .S(net510),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(net386),
    .A1(net1091),
    .S(net510),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(net382),
    .A1(net765),
    .S(net510),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(net375),
    .A1(net1032),
    .S(net510),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(net373),
    .A1(net1090),
    .S(net510),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(net370),
    .A1(net842),
    .S(net510),
    .X(_0593_));
 sky130_fd_sc_hd__nand2_8 _5432_ (.A(_0863_),
    .B(net363),
    .Y(_2430_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net401),
    .A1(net1545),
    .S(_2430_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _5434_ (.A0(net396),
    .A1(net910),
    .S(_2430_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net389),
    .A1(net1179),
    .S(_2430_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(net598),
    .A1(net720),
    .S(_2430_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(net647),
    .A1(net737),
    .S(_2430_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(net540),
    .A1(net600),
    .S(_2430_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(net372),
    .A1(net1158),
    .S(_2430_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(net369),
    .A1(net936),
    .S(_2430_),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_8 _5441_ (.A(net610),
    .B(net363),
    .Y(_2431_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(net401),
    .A1(net1542),
    .S(net611),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(net396),
    .A1(net823),
    .S(net611),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(net389),
    .A1(net1127),
    .S(net611),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(net598),
    .A1(\gpio_configure[20][3] ),
    .S(net611),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(net647),
    .A1(net651),
    .S(net611),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _5447_ (.A0(net375),
    .A1(net1094),
    .S(net611),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(net372),
    .A1(net1147),
    .S(net611),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(net369),
    .A1(net883),
    .S(net611),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_8 _5450_ (.A(_0890_),
    .B(net509),
    .Y(_2432_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(net401),
    .A1(net1524),
    .S(_2432_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(net396),
    .A1(net903),
    .S(_2432_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(net495),
    .A1(net1725),
    .S(_2432_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(net598),
    .A1(net690),
    .S(_2432_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(net647),
    .A1(net759),
    .S(_2432_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(net375),
    .A1(net1153),
    .S(_2432_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _5457_ (.A0(net372),
    .A1(net1191),
    .S(_2432_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(net369),
    .A1(net934),
    .S(_2432_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_8 _5459_ (.A(_0928_),
    .B(net363),
    .Y(_2433_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(net401),
    .A1(net1574),
    .S(_2433_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(net396),
    .A1(net835),
    .S(_2433_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(net389),
    .A1(net1238),
    .S(_2433_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(net598),
    .A1(net702),
    .S(_2433_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(net379),
    .A1(net1319),
    .S(_2433_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(net375),
    .A1(net1077),
    .S(_2433_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(net372),
    .A1(net1115),
    .S(_2433_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(net369),
    .A1(net868),
    .S(_2433_),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_8 _5468_ (.A(net658),
    .B(net363),
    .Y(_2434_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net401),
    .A1(net1540),
    .S(_2434_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(net396),
    .A1(net808),
    .S(_2434_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(net389),
    .A1(net1145),
    .S(_2434_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(net598),
    .A1(\gpio_configure[23][3] ),
    .S(_2434_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(net647),
    .A1(net1720),
    .S(_2434_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(net375),
    .A1(net1039),
    .S(_2434_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(net372),
    .A1(net1105),
    .S(_2434_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(net369),
    .A1(net885),
    .S(_2434_),
    .X(_0633_));
 sky130_fd_sc_hd__and2_4 _5477_ (.A(_0880_),
    .B(net363),
    .X(_2435_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(net1560),
    .A1(net401),
    .S(_2435_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _5479_ (.A0(net917),
    .A1(net396),
    .S(_2435_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(net1164),
    .A1(net389),
    .S(_2435_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _5481_ (.A0(net728),
    .A1(net598),
    .S(_2435_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(net733),
    .A1(net647),
    .S(_2435_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(net1117),
    .A1(net375),
    .S(_2435_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(net1183),
    .A1(net372),
    .S(_2435_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(net967),
    .A1(net369),
    .S(_2435_),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_8 _5486_ (.A(_0887_),
    .B(net562),
    .Y(_2436_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(net402),
    .A1(net1386),
    .S(_2436_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(net398),
    .A1(net827),
    .S(_2436_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(net390),
    .A1(net1400),
    .S(_2436_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(net533),
    .A1(net1726),
    .S(_2436_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(net381),
    .A1(net1315),
    .S(_2436_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _5492_ (.A0(net376),
    .A1(net918),
    .S(_2436_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _5493_ (.A0(net373),
    .A1(net1059),
    .S(_2436_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(net370),
    .A1(net825),
    .S(_2436_),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_8 _5495_ (.A(net750),
    .B(net366),
    .Y(_2437_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(net401),
    .A1(net1539),
    .S(_2437_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _5497_ (.A0(net398),
    .A1(\gpio_configure[26][1] ),
    .S(_2437_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(net392),
    .A1(net893),
    .S(_2437_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(net533),
    .A1(net625),
    .S(_2437_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(net382),
    .A1(net924),
    .S(_2437_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _5501_ (.A0(net376),
    .A1(net864),
    .S(_2437_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(net372),
    .A1(net1155),
    .S(_2437_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _5503_ (.A0(net370),
    .A1(net946),
    .S(_2437_),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_8 _5504_ (.A(net554),
    .B(net509),
    .Y(_2438_));
 sky130_fd_sc_hd__mux2_1 _5505_ (.A0(net401),
    .A1(net1568),
    .S(net555),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(net396),
    .A1(net882),
    .S(net555),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _5507_ (.A0(net505),
    .A1(net1712),
    .S(net555),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(net598),
    .A1(net701),
    .S(net555),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(net647),
    .A1(net710),
    .S(net555),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(net375),
    .A1(net1227),
    .S(net555),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(net671),
    .A1(net769),
    .S(net555),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(net369),
    .A1(net948),
    .S(net555),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_8 _5513_ (.A(_0953_),
    .B(net363),
    .Y(_2439_));
 sky130_fd_sc_hd__mux2_1 _5514_ (.A0(net401),
    .A1(net1573),
    .S(_2439_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(net396),
    .A1(net877),
    .S(_2439_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _5516_ (.A0(net505),
    .A1(net619),
    .S(_2439_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _5517_ (.A0(net598),
    .A1(net697),
    .S(_2439_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(net647),
    .A1(net761),
    .S(_2439_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(net375),
    .A1(net1132),
    .S(_2439_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _5520_ (.A0(net372),
    .A1(net1175),
    .S(_2439_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(net369),
    .A1(net862),
    .S(_2439_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_8 _5522_ (.A(net516),
    .B(net363),
    .Y(_2440_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(net401),
    .A1(net1541),
    .S(net517),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _5524_ (.A0(net396),
    .A1(net801),
    .S(net517),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(net505),
    .A1(net1719),
    .S(net517),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _5526_ (.A0(net598),
    .A1(net752),
    .S(net517),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(net647),
    .A1(net712),
    .S(net517),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(net375),
    .A1(net1129),
    .S(net517),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(net372),
    .A1(net1109),
    .S(net517),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(net369),
    .A1(net897),
    .S(net517),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_8 _5531_ (.A(net588),
    .B(net363),
    .Y(_2441_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(net401),
    .A1(net1549),
    .S(_2441_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _5533_ (.A0(net396),
    .A1(net822),
    .S(_2441_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(net505),
    .A1(net1713),
    .S(_2441_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _5535_ (.A0(net598),
    .A1(net683),
    .S(_2441_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(net631),
    .A1(net731),
    .S(_2441_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(net375),
    .A1(net1096),
    .S(_2441_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(net372),
    .A1(net1170),
    .S(_2441_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(net369),
    .A1(net880),
    .S(_2441_),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_8 _5540_ (.A(net483),
    .B(net363),
    .Y(_2442_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(net401),
    .A1(net1554),
    .S(net484),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _5542_ (.A0(net529),
    .A1(\gpio_configure[31][1] ),
    .S(net484),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net389),
    .A1(net1321),
    .S(net484),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _5544_ (.A0(net598),
    .A1(net696),
    .S(net484),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(net378),
    .A1(net1569),
    .S(net484),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(net540),
    .A1(net581),
    .S(net484),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(net372),
    .A1(net1101),
    .S(net484),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _5548_ (.A0(net476),
    .A1(net1703),
    .S(net484),
    .X(_0697_));
 sky130_fd_sc_hd__and2_4 _5549_ (.A(net547),
    .B(net366),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _5550_ (.A0(net1438),
    .A1(net402),
    .S(net548),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(net1009),
    .A1(net397),
    .S(net548),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(net1005),
    .A1(net392),
    .S(net548),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(net1046),
    .A1(net386),
    .S(net548),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(net1281),
    .A1(net381),
    .S(net548),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _5555_ (.A0(net1708),
    .A1(net540),
    .S(net548),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(net1107),
    .A1(net373),
    .S(net548),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(net1705),
    .A1(net476),
    .S(_2443_),
    .X(_0705_));
 sky130_fd_sc_hd__nand2_8 _5558_ (.A(_0960_),
    .B(net365),
    .Y(_2444_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(net402),
    .A1(net1446),
    .S(_2444_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(net529),
    .A1(net1729),
    .S(_2444_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(net389),
    .A1(net1287),
    .S(_2444_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _5562_ (.A0(net386),
    .A1(net1026),
    .S(_2444_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _5563_ (.A0(net381),
    .A1(net1295),
    .S(_2444_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _5564_ (.A0(net540),
    .A1(net604),
    .S(_2444_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(net372),
    .A1(net1160),
    .S(_2444_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _5566_ (.A0(net369),
    .A1(net942),
    .S(_2444_),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_8 _5567_ (.A(_0947_),
    .B(net509),
    .Y(_2445_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(net402),
    .A1(net1423),
    .S(_2445_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _5569_ (.A0(net396),
    .A1(net803),
    .S(_2445_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(net392),
    .A1(net899),
    .S(_2445_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(net386),
    .A1(net1063),
    .S(_2445_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(net647),
    .A1(net680),
    .S(_2445_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(net376),
    .A1(net850),
    .S(_2445_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(net372),
    .A1(net1113),
    .S(_2445_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _5575_ (.A0(net369),
    .A1(net901),
    .S(_2445_),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_8 _5576_ (.A(net523),
    .B(net363),
    .Y(_2446_));
 sky130_fd_sc_hd__mux2_1 _5577_ (.A0(net1347),
    .A1(net1385),
    .S(net524),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(net396),
    .A1(net824),
    .S(net524),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(net505),
    .A1(net1716),
    .S(net524),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(net598),
    .A1(net706),
    .S(net524),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _5581_ (.A0(net382),
    .A1(net1330),
    .S(net524),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(net375),
    .A1(net1123),
    .S(net524),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net372),
    .A1(net1185),
    .S(net524),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _5584_ (.A0(net369),
    .A1(net889),
    .S(net524),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_8 _5585_ (.A(_0935_),
    .B(net366),
    .Y(_2447_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(net402),
    .A1(net1450),
    .S(_2447_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net397),
    .A1(net923),
    .S(_2447_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net390),
    .A1(net1593),
    .S(_2447_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(net533),
    .A1(\gpio_configure[36][3] ),
    .S(_2447_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(net381),
    .A1(net1301),
    .S(_2447_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net376),
    .A1(net913),
    .S(_2447_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(net671),
    .A1(net1721),
    .S(_2447_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net370),
    .A1(net811),
    .S(_2447_),
    .X(_0737_));
 sky130_fd_sc_hd__nand2_8 _5594_ (.A(_0939_),
    .B(net366),
    .Y(_2448_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(net402),
    .A1(net1465),
    .S(_2448_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(net398),
    .A1(net845),
    .S(_2448_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net392),
    .A1(net995),
    .S(_2448_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(net533),
    .A1(net602),
    .S(_2448_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net381),
    .A1(net1325),
    .S(_2448_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(net376),
    .A1(net926),
    .S(_2448_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net373),
    .A1(net1065),
    .S(_2448_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _5602_ (.A0(net370),
    .A1(net852),
    .S(_2448_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_4 _5603_ (.A(net407),
    .B(\xfer_state[2] ),
    .Y(_2449_));
 sky130_fd_sc_hd__o31a_4 _5604_ (.A1(net407),
    .A2(\xfer_state[3] ),
    .A3(\xfer_state[2] ),
    .B1(_1455_),
    .X(_2450_));
 sky130_fd_sc_hd__inv_2 _5605_ (.A(_2450_),
    .Y(_2451_));
 sky130_fd_sc_hd__or3_2 _5606_ (.A(\xfer_state[3] ),
    .B(_1456_),
    .C(_2449_),
    .X(_2452_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(\xfer_count[0] ),
    .B(_2450_),
    .Y(_2453_));
 sky130_fd_sc_hd__or2_1 _5608_ (.A(\xfer_count[0] ),
    .B(_2450_),
    .X(_2454_));
 sky130_fd_sc_hd__and3_1 _5609_ (.A(_2452_),
    .B(_2453_),
    .C(_2454_),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _5611_ (.A(net408),
    .B(\xfer_state[3] ),
    .Y(_2456_));
 sky130_fd_sc_hd__nor2_1 _5612_ (.A(_1448_),
    .B(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__a32o_1 _5613_ (.A1(_1455_),
    .A2(_2455_),
    .A3(_2457_),
    .B1(_2451_),
    .B2(\xfer_count[1] ),
    .X(_0747_));
 sky130_fd_sc_hd__a31o_1 _5614_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[1] ),
    .A3(_2450_),
    .B1(\xfer_count[2] ),
    .X(_2458_));
 sky130_fd_sc_hd__and4_2 _5615_ (.A(\xfer_count[0] ),
    .B(\xfer_count[1] ),
    .C(\xfer_count[2] ),
    .D(_2450_),
    .X(_2459_));
 sky130_fd_sc_hd__inv_2 _5616_ (.A(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__and3_1 _5617_ (.A(_2452_),
    .B(_2458_),
    .C(_2460_),
    .X(_0748_));
 sky130_fd_sc_hd__a21boi_1 _5618_ (.A1(\xfer_count[3] ),
    .A2(_2459_),
    .B1_N(_2452_),
    .Y(_2461_));
 sky130_fd_sc_hd__o21a_1 _5619_ (.A1(\xfer_count[3] ),
    .A2(_2459_),
    .B1(_2461_),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_2 _5620_ (.A(\xfer_state[0] ),
    .B(\xfer_state[2] ),
    .Y(_2462_));
 sky130_fd_sc_hd__or2_2 _5621_ (.A(\xfer_state[0] ),
    .B(\xfer_state[2] ),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _5622_ (.A0(\xfer_state[2] ),
    .A1(_2462_),
    .S(\pad_count_1[0] ),
    .X(_0750_));
 sky130_fd_sc_hd__nor2_8 _5623_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .Y(_2464_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(\xfer_state[2] ),
    .B(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__and2_4 _5625_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2466_));
 sky130_fd_sc_hd__nor2_4 _5626_ (.A(_0820_),
    .B(\xfer_state[2] ),
    .Y(_2467_));
 sky130_fd_sc_hd__nand2_4 _5627_ (.A(\xfer_state[0] ),
    .B(_0822_),
    .Y(_2468_));
 sky130_fd_sc_hd__o32a_1 _5628_ (.A1(_0822_),
    .A2(_2464_),
    .A3(_2466_),
    .B1(\pad_count_1[1] ),
    .B2(_2463_),
    .X(_0751_));
 sky130_fd_sc_hd__or2_2 _5629_ (.A(\pad_count_1[2] ),
    .B(_2465_),
    .X(_2469_));
 sky130_fd_sc_hd__inv_2 _5630_ (.A(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__a31o_1 _5631_ (.A1(\pad_count_1[2] ),
    .A2(_2465_),
    .A3(_2468_),
    .B1(_2470_),
    .X(_0752_));
 sky130_fd_sc_hd__nor2_8 _5632_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .Y(_2471_));
 sky130_fd_sc_hd__nor2_1 _5633_ (.A(\pad_count_1[3] ),
    .B(_2469_),
    .Y(_2472_));
 sky130_fd_sc_hd__a31o_1 _5634_ (.A1(\pad_count_1[3] ),
    .A2(_2468_),
    .A3(_2469_),
    .B1(_2472_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(net404),
    .B(_2468_),
    .Y(_2473_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(_2473_),
    .A1(_0830_),
    .S(_2472_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _5637_ (.A0(_2463_),
    .A1(_0822_),
    .S(\pad_count_2[0] ),
    .X(_0755_));
 sky130_fd_sc_hd__and2_4 _5638_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2474_));
 sky130_fd_sc_hd__and3_2 _5639_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .C(\xfer_state[2] ),
    .X(_2475_));
 sky130_fd_sc_hd__and2b_4 _5640_ (.A_N(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2476_));
 sky130_fd_sc_hd__o32a_1 _5641_ (.A1(_0822_),
    .A2(_1444_),
    .A3(_2476_),
    .B1(_2463_),
    .B2(\pad_count_2[1] ),
    .X(_0756_));
 sky130_fd_sc_hd__a21oi_1 _5642_ (.A1(\pad_count_2[2] ),
    .A2(_2468_),
    .B1(_2475_),
    .Y(_2477_));
 sky130_fd_sc_hd__a21oi_1 _5643_ (.A1(\pad_count_2[2] ),
    .A2(_2475_),
    .B1(_2477_),
    .Y(_0757_));
 sky130_fd_sc_hd__and2_4 _5644_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .X(_2478_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_2475_),
    .B(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__and3_1 _5646_ (.A(\xfer_state[2] ),
    .B(_1445_),
    .C(_2474_),
    .X(_2480_));
 sky130_fd_sc_hd__a31o_1 _5647_ (.A1(\pad_count_2[3] ),
    .A2(_2468_),
    .A3(_2479_),
    .B1(_2480_),
    .X(_0758_));
 sky130_fd_sc_hd__and3_1 _5648_ (.A(\pad_count_2[4] ),
    .B(_2475_),
    .C(_2478_),
    .X(_2481_));
 sky130_fd_sc_hd__nor2_1 _5649_ (.A(\pad_count_2[4] ),
    .B(_2467_),
    .Y(_2482_));
 sky130_fd_sc_hd__a21oi_1 _5650_ (.A1(_2479_),
    .A2(_2482_),
    .B1(_2481_),
    .Y(_0759_));
 sky130_fd_sc_hd__and2b_4 _5651_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .X(_2483_));
 sky130_fd_sc_hd__nand2b_4 _5652_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .Y(_2484_));
 sky130_fd_sc_hd__and3_4 _5653_ (.A(_2474_),
    .B(_2478_),
    .C(_2483_),
    .X(_2485_));
 sky130_fd_sc_hd__nor2_1 _5654_ (.A(_2467_),
    .B(_2481_),
    .Y(_2486_));
 sky130_fd_sc_hd__a22o_1 _5655_ (.A1(\xfer_state[2] ),
    .A2(_2485_),
    .B1(_2486_),
    .B2(\pad_count_2[5] ),
    .X(_0760_));
 sky130_fd_sc_hd__or3b_1 _5656_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C_N(_2455_),
    .X(_2487_));
 sky130_fd_sc_hd__a22o_1 _5657_ (.A1(_2456_),
    .A2(_2462_),
    .B1(_2487_),
    .B2(\xfer_state[3] ),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _5658_ (.A0(_1450_),
    .A1(serial_clock_pre),
    .S(_2488_),
    .X(_0761_));
 sky130_fd_sc_hd__or4b_1 _5659_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C(_0821_),
    .D_N(\xfer_count[0] ),
    .X(_2489_));
 sky130_fd_sc_hd__a2bb2o_1 _5660_ (.A1_N(\xfer_count[1] ),
    .A2_N(_2489_),
    .B1(_2488_),
    .B2(serial_load_pre),
    .X(_0762_));
 sky130_fd_sc_hd__a21o_1 _5661_ (.A1(\xfer_state[0] ),
    .A2(_0821_),
    .B1(serial_busy),
    .X(_2490_));
 sky130_fd_sc_hd__o311a_1 _5662_ (.A1(serial_xfer),
    .A2(_0820_),
    .A3(\xfer_state[3] ),
    .B1(_1454_),
    .C1(_2490_),
    .X(_0763_));
 sky130_fd_sc_hd__nor2_2 _5663_ (.A(net407),
    .B(_0822_),
    .Y(_2491_));
 sky130_fd_sc_hd__or2_4 _5664_ (.A(_1450_),
    .B(_2449_),
    .X(_2492_));
 sky130_fd_sc_hd__nor2_8 _5665_ (.A(_1450_),
    .B(_2449_),
    .Y(_2493_));
 sky130_fd_sc_hd__and2b_4 _5666_ (.A_N(\pad_count_1[0] ),
    .B(\pad_count_1[1] ),
    .X(_2494_));
 sky130_fd_sc_hd__and3_4 _5667_ (.A(\pad_count_1[4] ),
    .B(_2471_),
    .C(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__and2b_4 _5668_ (.A_N(\pad_count_1[2] ),
    .B(\pad_count_1[3] ),
    .X(_2496_));
 sky130_fd_sc_hd__and3_4 _5669_ (.A(\pad_count_1[4] ),
    .B(_2494_),
    .C(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__a22o_1 _5670_ (.A1(\gpio_configure[18][0] ),
    .A2(_2495_),
    .B1(_2497_),
    .B2(\gpio_configure[26][0] ),
    .X(_2498_));
 sky130_fd_sc_hd__and2b_4 _5671_ (.A_N(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2499_));
 sky130_fd_sc_hd__and2_4 _5672_ (.A(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .X(_2500_));
 sky130_fd_sc_hd__and3_4 _5673_ (.A(net404),
    .B(_2499_),
    .C(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__and3_4 _5674_ (.A(net404),
    .B(_2466_),
    .C(_2471_),
    .X(_2502_));
 sky130_fd_sc_hd__and3_4 _5675_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2500_),
    .X(_2503_));
 sky130_fd_sc_hd__and3_4 _5676_ (.A(net404),
    .B(_2466_),
    .C(_2500_),
    .X(_2504_));
 sky130_fd_sc_hd__a22o_1 _5677_ (.A1(\gpio_configure[31][0] ),
    .A2(_2503_),
    .B1(_2504_),
    .B2(\gpio_configure[15][0] ),
    .X(_2505_));
 sky130_fd_sc_hd__and3_4 _5678_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2471_),
    .X(_2506_));
 sky130_fd_sc_hd__and2b_4 _5679_ (.A_N(\pad_count_1[3] ),
    .B(\pad_count_1[2] ),
    .X(_2507_));
 sky130_fd_sc_hd__and3_4 _5680_ (.A(net404),
    .B(_2466_),
    .C(_2507_),
    .X(_2508_));
 sky130_fd_sc_hd__and3_4 _5681_ (.A(net404),
    .B(_2464_),
    .C(_2496_),
    .X(_2509_));
 sky130_fd_sc_hd__and3_4 _5682_ (.A(\pad_count_1[4] ),
    .B(_2464_),
    .C(_2507_),
    .X(_2510_));
 sky130_fd_sc_hd__and3_4 _5683_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2507_),
    .X(_2511_));
 sky130_fd_sc_hd__and3_4 _5684_ (.A(\pad_count_1[4] ),
    .B(_2471_),
    .C(_2499_),
    .X(_2512_));
 sky130_fd_sc_hd__and3_4 _5685_ (.A(\pad_count_1[4] ),
    .B(_2499_),
    .C(_2500_),
    .X(_2513_));
 sky130_fd_sc_hd__a22o_1 _5686_ (.A1(\gpio_configure[17][0] ),
    .A2(_2512_),
    .B1(_2513_),
    .B2(\gpio_configure[29][0] ),
    .X(_2514_));
 sky130_fd_sc_hd__and3_4 _5687_ (.A(\pad_count_1[4] ),
    .B(_2464_),
    .C(_2496_),
    .X(_2515_));
 sky130_fd_sc_hd__and3_4 _5688_ (.A(\pad_count_1[4] ),
    .B(_2494_),
    .C(_2507_),
    .X(_2516_));
 sky130_fd_sc_hd__and3_4 _5689_ (.A(net404),
    .B(_2494_),
    .C(_2507_),
    .X(_2517_));
 sky130_fd_sc_hd__and3_4 _5690_ (.A(\pad_count_1[4] ),
    .B(_2494_),
    .C(_2500_),
    .X(_2518_));
 sky130_fd_sc_hd__and3_4 _5691_ (.A(net404),
    .B(_2494_),
    .C(_2500_),
    .X(_2519_));
 sky130_fd_sc_hd__and3_4 _5692_ (.A(\pad_count_1[4] ),
    .B(_2466_),
    .C(_2496_),
    .X(_2520_));
 sky130_fd_sc_hd__and3_4 _5693_ (.A(\pad_count_1[4] ),
    .B(_2464_),
    .C(_2500_),
    .X(_2521_));
 sky130_fd_sc_hd__and3_4 _5694_ (.A(net404),
    .B(_2499_),
    .C(_2507_),
    .X(_2522_));
 sky130_fd_sc_hd__a22o_1 _5695_ (.A1(\gpio_configure[28][0] ),
    .A2(_2521_),
    .B1(_2522_),
    .B2(\gpio_configure[5][0] ),
    .X(_2523_));
 sky130_fd_sc_hd__and2_4 _5696_ (.A(_2464_),
    .B(_2471_),
    .X(_2524_));
 sky130_fd_sc_hd__and3_4 _5697_ (.A(net404),
    .B(_2464_),
    .C(_2471_),
    .X(_2525_));
 sky130_fd_sc_hd__nand2_8 _5698_ (.A(net404),
    .B(_2524_),
    .Y(_2526_));
 sky130_fd_sc_hd__and3_4 _5699_ (.A(net404),
    .B(_2496_),
    .C(_2499_),
    .X(_2527_));
 sky130_fd_sc_hd__and3_4 _5700_ (.A(net404),
    .B(_2471_),
    .C(_2499_),
    .X(_2528_));
 sky130_fd_sc_hd__and3_4 _5701_ (.A(net404),
    .B(_2464_),
    .C(_2500_),
    .X(_2529_));
 sky130_fd_sc_hd__and3_4 _5702_ (.A(net404),
    .B(_2464_),
    .C(_2507_),
    .X(_2530_));
 sky130_fd_sc_hd__and3_4 _5703_ (.A(net404),
    .B(_2471_),
    .C(_2494_),
    .X(_2531_));
 sky130_fd_sc_hd__and3_4 _5704_ (.A(net404),
    .B(_2494_),
    .C(_2496_),
    .X(_2532_));
 sky130_fd_sc_hd__and3_4 _5705_ (.A(net404),
    .B(_2466_),
    .C(_2496_),
    .X(_2533_));
 sky130_fd_sc_hd__and3_4 _5706_ (.A(\pad_count_1[4] ),
    .B(_2496_),
    .C(_2499_),
    .X(_2534_));
 sky130_fd_sc_hd__and3_4 _5707_ (.A(\pad_count_1[4] ),
    .B(_2499_),
    .C(_2507_),
    .X(_2535_));
 sky130_fd_sc_hd__a221o_1 _5708_ (.A1(\gpio_configure[22][0] ),
    .A2(_2516_),
    .B1(_2535_),
    .B2(\gpio_configure[21][0] ),
    .C1(_2498_),
    .X(_2536_));
 sky130_fd_sc_hd__a221o_2 _5709_ (.A1(\gpio_configure[24][0] ),
    .A2(_2515_),
    .B1(_2529_),
    .B2(\gpio_configure[12][0] ),
    .C1(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__a21o_1 _5710_ (.A1(\gpio_configure[13][0] ),
    .A2(_2501_),
    .B1(_2523_),
    .X(_2538_));
 sky130_fd_sc_hd__a22o_1 _5711_ (.A1(\gpio_configure[19][0] ),
    .A2(_2506_),
    .B1(_2530_),
    .B2(\gpio_configure[4][0] ),
    .X(_2539_));
 sky130_fd_sc_hd__a221o_2 _5712_ (.A1(\gpio_configure[3][0] ),
    .A2(_2502_),
    .B1(_2518_),
    .B2(\gpio_configure[30][0] ),
    .C1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__a211o_4 _5713_ (.A1(\gpio_configure[6][0] ),
    .A2(_2517_),
    .B1(_2538_),
    .C1(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__a221o_1 _5714_ (.A1(\gpio_configure[16][0] ),
    .A2(_2524_),
    .B1(_2533_),
    .B2(\gpio_configure[11][0] ),
    .C1(_2525_),
    .X(_2542_));
 sky130_fd_sc_hd__a221o_2 _5715_ (.A1(\gpio_configure[14][0] ),
    .A2(_2519_),
    .B1(_2532_),
    .B2(\gpio_configure[10][0] ),
    .C1(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__a221o_1 _5716_ (.A1(\gpio_configure[1][0] ),
    .A2(_2528_),
    .B1(_2534_),
    .B2(\gpio_configure[25][0] ),
    .C1(_2514_),
    .X(_2544_));
 sky130_fd_sc_hd__a22o_1 _5717_ (.A1(\gpio_configure[7][0] ),
    .A2(_2508_),
    .B1(_2531_),
    .B2(\gpio_configure[2][0] ),
    .X(_2545_));
 sky130_fd_sc_hd__a221o_2 _5718_ (.A1(\gpio_configure[23][0] ),
    .A2(_2511_),
    .B1(_2527_),
    .B2(\gpio_configure[9][0] ),
    .C1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__a221o_1 _5719_ (.A1(\gpio_configure[8][0] ),
    .A2(_2509_),
    .B1(_2510_),
    .B2(\gpio_configure[20][0] ),
    .C1(_2505_),
    .X(_2547_));
 sky130_fd_sc_hd__or4_4 _5720_ (.A(_2543_),
    .B(_2544_),
    .C(_2546_),
    .D(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a2111o_4 _5721_ (.A1(\gpio_configure[27][0] ),
    .A2(_2520_),
    .B1(_2537_),
    .C1(_2541_),
    .D1(_2548_),
    .X(_2549_));
 sky130_fd_sc_hd__or2_1 _5722_ (.A(\gpio_configure[0][0] ),
    .B(_2526_),
    .X(_2550_));
 sky130_fd_sc_hd__a32o_1 _5723_ (.A1(_2491_),
    .A2(_2549_),
    .A3(_2550_),
    .B1(net353),
    .B2(\serial_data_staging_1[0] ),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _5724_ (.A1(\gpio_configure[18][1] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][1] ),
    .X(_2551_));
 sky130_fd_sc_hd__a22o_1 _5725_ (.A1(\gpio_configure[5][1] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][1] ),
    .X(_2552_));
 sky130_fd_sc_hd__a22o_1 _5726_ (.A1(\gpio_configure[29][1] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][1] ),
    .X(_2553_));
 sky130_fd_sc_hd__a221o_1 _5727_ (.A1(\gpio_configure[23][1] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][1] ),
    .C1(_2551_),
    .X(_2554_));
 sky130_fd_sc_hd__a22o_1 _5728_ (.A1(\gpio_configure[14][1] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][1] ),
    .X(_2555_));
 sky130_fd_sc_hd__a221o_4 _5729_ (.A1(\gpio_configure[13][1] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][1] ),
    .C1(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__a22o_1 _5730_ (.A1(\gpio_configure[3][1] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][1] ),
    .X(_2557_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(\gpio_configure[31][1] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][1] ),
    .C1(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a221o_1 _5732_ (.A1(\gpio_configure[26][1] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(\gpio_configure[16][1] ),
    .C1(_2525_),
    .X(_2559_));
 sky130_fd_sc_hd__a221o_4 _5733_ (.A1(\gpio_configure[15][1] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][1] ),
    .C1(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__or4_2 _5734_ (.A(_2554_),
    .B(_2556_),
    .C(_2558_),
    .D(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(\gpio_configure[7][1] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][1] ),
    .C1(_2553_),
    .X(_2562_));
 sky130_fd_sc_hd__a211o_4 _5736_ (.A1(\gpio_configure[6][1] ),
    .A2(_2517_),
    .B1(_2552_),
    .C1(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a22o_1 _5737_ (.A1(\gpio_configure[20][1] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][1] ),
    .X(_2564_));
 sky130_fd_sc_hd__a221o_1 _5738_ (.A1(\gpio_configure[30][1] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][1] ),
    .C1(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__a22o_1 _5739_ (.A1(\gpio_configure[19][1] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][1] ),
    .X(_2566_));
 sky130_fd_sc_hd__a221o_1 _5740_ (.A1(\gpio_configure[11][1] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][1] ),
    .C1(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__or3_1 _5741_ (.A(_2563_),
    .B(_2565_),
    .C(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__o221a_2 _5742_ (.A1(\gpio_configure[0][1] ),
    .A2(_2526_),
    .B1(_2561_),
    .B2(_2568_),
    .C1(_0819_),
    .X(_2569_));
 sky130_fd_sc_hd__a21o_1 _5743_ (.A1(net407),
    .A2(\serial_data_staging_1[0] ),
    .B1(net353),
    .X(_2570_));
 sky130_fd_sc_hd__o22a_1 _5744_ (.A1(\serial_data_staging_1[1] ),
    .A2(net352),
    .B1(_2569_),
    .B2(_2570_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _5745_ (.A1(\gpio_configure[15][2] ),
    .A2(_2504_),
    .B1(_2531_),
    .B2(\gpio_configure[2][2] ),
    .X(_2571_));
 sky130_fd_sc_hd__a221o_1 _5746_ (.A1(\gpio_configure[31][2] ),
    .A2(_2503_),
    .B1(_2529_),
    .B2(\gpio_configure[12][2] ),
    .C1(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__a22o_1 _5747_ (.A1(\gpio_configure[17][2] ),
    .A2(_2512_),
    .B1(_2520_),
    .B2(\gpio_configure[27][2] ),
    .X(_2573_));
 sky130_fd_sc_hd__a221o_4 _5748_ (.A1(\gpio_configure[20][2] ),
    .A2(_2510_),
    .B1(_2513_),
    .B2(\gpio_configure[29][2] ),
    .C1(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__a22o_1 _5749_ (.A1(\gpio_configure[10][2] ),
    .A2(_2532_),
    .B1(_2534_),
    .B2(\gpio_configure[25][2] ),
    .X(_2575_));
 sky130_fd_sc_hd__a21o_1 _5750_ (.A1(\gpio_configure[5][2] ),
    .A2(_2522_),
    .B1(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__a22o_2 _5751_ (.A1(\gpio_configure[22][2] ),
    .A2(_2516_),
    .B1(_2521_),
    .B2(\gpio_configure[28][2] ),
    .X(_2577_));
 sky130_fd_sc_hd__a221o_1 _5752_ (.A1(\gpio_configure[1][2] ),
    .A2(_2528_),
    .B1(_2533_),
    .B2(\gpio_configure[11][2] ),
    .C1(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__or4_4 _5753_ (.A(_2572_),
    .B(_2574_),
    .C(_2576_),
    .D(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__a22o_1 _5754_ (.A1(\gpio_configure[13][2] ),
    .A2(_2501_),
    .B1(_2519_),
    .B2(\gpio_configure[14][2] ),
    .X(_2580_));
 sky130_fd_sc_hd__a221o_2 _5755_ (.A1(\gpio_configure[3][2] ),
    .A2(_2502_),
    .B1(_2509_),
    .B2(\gpio_configure[8][2] ),
    .C1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__or2_1 _5756_ (.A(\gpio_configure[16][2] ),
    .B(_0830_),
    .X(_2582_));
 sky130_fd_sc_hd__a22o_4 _5757_ (.A1(\gpio_configure[4][2] ),
    .A2(_2530_),
    .B1(_2582_),
    .B2(_2524_),
    .X(_2583_));
 sky130_fd_sc_hd__a221o_4 _5758_ (.A1(\gpio_configure[18][2] ),
    .A2(_2495_),
    .B1(_2511_),
    .B2(\gpio_configure[23][2] ),
    .C1(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__a22o_1 _5759_ (.A1(\gpio_configure[6][2] ),
    .A2(_2517_),
    .B1(_2535_),
    .B2(\gpio_configure[21][2] ),
    .X(_2585_));
 sky130_fd_sc_hd__a221o_1 _5760_ (.A1(\gpio_configure[19][2] ),
    .A2(_2506_),
    .B1(_2527_),
    .B2(\gpio_configure[9][2] ),
    .C1(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__a22o_1 _5761_ (.A1(\gpio_configure[26][2] ),
    .A2(_2497_),
    .B1(_2518_),
    .B2(\gpio_configure[30][2] ),
    .X(_2587_));
 sky130_fd_sc_hd__a221o_1 _5762_ (.A1(\gpio_configure[7][2] ),
    .A2(_2508_),
    .B1(_2515_),
    .B2(\gpio_configure[24][2] ),
    .C1(_2587_),
    .X(_2588_));
 sky130_fd_sc_hd__or4_4 _5763_ (.A(_2581_),
    .B(_2584_),
    .C(_2586_),
    .D(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__o221a_4 _5764_ (.A1(\gpio_configure[0][2] ),
    .A2(_2526_),
    .B1(_2579_),
    .B2(_2589_),
    .C1(net405),
    .X(_2590_));
 sky130_fd_sc_hd__a21o_1 _5765_ (.A1(net407),
    .A2(\serial_data_staging_1[1] ),
    .B1(net353),
    .X(_2591_));
 sky130_fd_sc_hd__o22a_1 _5766_ (.A1(\serial_data_staging_1[2] ),
    .A2(net352),
    .B1(_2590_),
    .B2(_2591_),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _5767_ (.A1(\gpio_configure[5][3] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][3] ),
    .X(_2592_));
 sky130_fd_sc_hd__a22o_1 _5768_ (.A1(\gpio_configure[29][3] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][3] ),
    .X(_2593_));
 sky130_fd_sc_hd__a22o_1 _5769_ (.A1(\gpio_configure[18][3] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][3] ),
    .X(_2594_));
 sky130_fd_sc_hd__a221o_1 _5770_ (.A1(\gpio_configure[23][3] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][3] ),
    .C1(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__a22o_1 _5771_ (.A1(\gpio_configure[14][3] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][3] ),
    .X(_2596_));
 sky130_fd_sc_hd__a221o_1 _5772_ (.A1(\gpio_configure[13][3] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][3] ),
    .C1(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__a22o_1 _5773_ (.A1(\gpio_configure[31][3] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][3] ),
    .X(_2598_));
 sky130_fd_sc_hd__a221o_1 _5774_ (.A1(\gpio_configure[3][3] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][3] ),
    .C1(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__a221o_1 _5775_ (.A1(\gpio_configure[26][3] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(\gpio_configure[16][3] ),
    .C1(_2525_),
    .X(_2600_));
 sky130_fd_sc_hd__a221o_1 _5776_ (.A1(\gpio_configure[15][3] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][3] ),
    .C1(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__or4_4 _5777_ (.A(_2595_),
    .B(_2597_),
    .C(_2599_),
    .D(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__a221o_1 _5778_ (.A1(\gpio_configure[7][3] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][3] ),
    .C1(_2593_),
    .X(_2603_));
 sky130_fd_sc_hd__a211o_2 _5779_ (.A1(\gpio_configure[6][3] ),
    .A2(_2517_),
    .B1(_2592_),
    .C1(_2603_),
    .X(_2604_));
 sky130_fd_sc_hd__a22o_1 _5780_ (.A1(\gpio_configure[20][3] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][3] ),
    .X(_2605_));
 sky130_fd_sc_hd__a221o_1 _5781_ (.A1(\gpio_configure[30][3] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][3] ),
    .C1(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__a22o_1 _5782_ (.A1(\gpio_configure[19][3] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][3] ),
    .X(_2607_));
 sky130_fd_sc_hd__a221o_1 _5783_ (.A1(\gpio_configure[11][3] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][3] ),
    .C1(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__or3_4 _5784_ (.A(_2604_),
    .B(_2606_),
    .C(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__o221a_1 _5785_ (.A1(\gpio_configure[0][3] ),
    .A2(_2526_),
    .B1(_2602_),
    .B2(_2609_),
    .C1(_0819_),
    .X(_2610_));
 sky130_fd_sc_hd__a21o_1 _5786_ (.A1(net407),
    .A2(\serial_data_staging_1[2] ),
    .B1(net353),
    .X(_2611_));
 sky130_fd_sc_hd__o22a_1 _5787_ (.A1(\serial_data_staging_1[3] ),
    .A2(net352),
    .B1(_2610_),
    .B2(_2611_),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _5788_ (.A1(\gpio_configure[19][4] ),
    .A2(_2506_),
    .B1(_2512_),
    .B2(\gpio_configure[17][4] ),
    .X(_2612_));
 sky130_fd_sc_hd__a221o_1 _5789_ (.A1(\gpio_configure[3][4] ),
    .A2(_2502_),
    .B1(_2522_),
    .B2(\gpio_configure[5][4] ),
    .C1(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a22o_1 _5790_ (.A1(\gpio_configure[14][4] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][4] ),
    .X(_2614_));
 sky130_fd_sc_hd__a221o_4 _5791_ (.A1(\gpio_configure[22][4] ),
    .A2(_2516_),
    .B1(_2530_),
    .B2(\gpio_configure[4][4] ),
    .C1(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__a22o_1 _5792_ (.A1(\gpio_configure[6][4] ),
    .A2(_2517_),
    .B1(_2533_),
    .B2(\gpio_configure[11][4] ),
    .X(_2616_));
 sky130_fd_sc_hd__a21o_1 _5793_ (.A1(\gpio_configure[18][4] ),
    .A2(_2495_),
    .B1(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__a22o_1 _5794_ (.A1(\gpio_configure[28][4] ),
    .A2(_2521_),
    .B1(_2531_),
    .B2(\gpio_configure[2][4] ),
    .X(_2618_));
 sky130_fd_sc_hd__a221o_1 _5795_ (.A1(\gpio_configure[9][4] ),
    .A2(_2527_),
    .B1(_2535_),
    .B2(\gpio_configure[21][4] ),
    .C1(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__or4_2 _5796_ (.A(_2613_),
    .B(_2615_),
    .C(_2617_),
    .D(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__a22o_2 _5797_ (.A1(\gpio_configure[13][4] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][4] ),
    .X(_2621_));
 sky130_fd_sc_hd__a221o_1 _5798_ (.A1(\gpio_configure[30][4] ),
    .A2(_2518_),
    .B1(_2520_),
    .B2(\gpio_configure[27][4] ),
    .C1(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__or2_1 _5799_ (.A(\gpio_configure[16][4] ),
    .B(_0830_),
    .X(_2623_));
 sky130_fd_sc_hd__a22o_2 _5800_ (.A1(\gpio_configure[10][4] ),
    .A2(_2532_),
    .B1(_2623_),
    .B2(_2524_),
    .X(_2624_));
 sky130_fd_sc_hd__a221o_1 _5801_ (.A1(\gpio_configure[20][4] ),
    .A2(_2510_),
    .B1(_2534_),
    .B2(\gpio_configure[25][4] ),
    .C1(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__a22o_1 _5802_ (.A1(\gpio_configure[7][4] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][4] ),
    .X(_2626_));
 sky130_fd_sc_hd__a221o_1 _5803_ (.A1(\gpio_configure[31][4] ),
    .A2(_2503_),
    .B1(_2511_),
    .B2(\gpio_configure[23][4] ),
    .C1(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__a22o_1 _5804_ (.A1(\gpio_configure[26][4] ),
    .A2(_2497_),
    .B1(_2515_),
    .B2(\gpio_configure[24][4] ),
    .X(_2628_));
 sky130_fd_sc_hd__a221o_1 _5805_ (.A1(\gpio_configure[15][4] ),
    .A2(_2504_),
    .B1(_2513_),
    .B2(\gpio_configure[29][4] ),
    .C1(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__or4_2 _5806_ (.A(_2622_),
    .B(_2625_),
    .C(_2627_),
    .D(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__o221a_4 _5807_ (.A1(\gpio_configure[0][4] ),
    .A2(_2526_),
    .B1(_2620_),
    .B2(_2630_),
    .C1(net405),
    .X(_2631_));
 sky130_fd_sc_hd__a211o_1 _5808_ (.A1(net407),
    .A2(\serial_data_staging_1[3] ),
    .B1(net353),
    .C1(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__o21a_1 _5809_ (.A1(\serial_data_staging_1[4] ),
    .A2(net352),
    .B1(_2632_),
    .X(_0768_));
 sky130_fd_sc_hd__a22o_1 _5810_ (.A1(\gpio_configure[18][5] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][5] ),
    .X(_2633_));
 sky130_fd_sc_hd__a22o_1 _5811_ (.A1(\gpio_configure[29][5] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][5] ),
    .X(_2634_));
 sky130_fd_sc_hd__a22o_2 _5812_ (.A1(\gpio_configure[5][5] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][5] ),
    .X(_2635_));
 sky130_fd_sc_hd__a221o_1 _5813_ (.A1(\gpio_configure[7][5] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][5] ),
    .C1(_2634_),
    .X(_2636_));
 sky130_fd_sc_hd__a211o_4 _5814_ (.A1(\gpio_configure[6][5] ),
    .A2(_2517_),
    .B1(_2635_),
    .C1(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__a22o_1 _5815_ (.A1(\gpio_configure[20][5] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][5] ),
    .X(_2638_));
 sky130_fd_sc_hd__a221o_2 _5816_ (.A1(\gpio_configure[30][5] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][5] ),
    .C1(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__a22o_1 _5817_ (.A1(\gpio_configure[19][5] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][5] ),
    .X(_2640_));
 sky130_fd_sc_hd__a221o_1 _5818_ (.A1(\gpio_configure[11][5] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][5] ),
    .C1(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__a221o_1 _5819_ (.A1(\gpio_configure[23][5] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][5] ),
    .C1(_2633_),
    .X(_2642_));
 sky130_fd_sc_hd__a22o_1 _5820_ (.A1(\gpio_configure[14][5] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][5] ),
    .X(_2643_));
 sky130_fd_sc_hd__a221o_4 _5821_ (.A1(\gpio_configure[13][5] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][5] ),
    .C1(_2643_),
    .X(_2644_));
 sky130_fd_sc_hd__a22o_1 _5822_ (.A1(\gpio_configure[3][5] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][5] ),
    .X(_2645_));
 sky130_fd_sc_hd__a221o_1 _5823_ (.A1(\gpio_configure[31][5] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][5] ),
    .C1(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__a221o_1 _5824_ (.A1(\gpio_configure[26][5] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(\gpio_configure[16][5] ),
    .C1(_2525_),
    .X(_2647_));
 sky130_fd_sc_hd__a221o_2 _5825_ (.A1(\gpio_configure[15][5] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][5] ),
    .C1(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__or4_2 _5826_ (.A(_2642_),
    .B(_2644_),
    .C(_2646_),
    .D(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__or3_2 _5827_ (.A(_2637_),
    .B(_2639_),
    .C(_2641_),
    .X(_2650_));
 sky130_fd_sc_hd__o221a_4 _5828_ (.A1(\gpio_configure[0][5] ),
    .A2(_2526_),
    .B1(_2649_),
    .B2(_2650_),
    .C1(net405),
    .X(_2651_));
 sky130_fd_sc_hd__a21o_1 _5829_ (.A1(net407),
    .A2(\serial_data_staging_1[4] ),
    .B1(net353),
    .X(_2652_));
 sky130_fd_sc_hd__o22a_1 _5830_ (.A1(\serial_data_staging_1[5] ),
    .A2(net352),
    .B1(_2651_),
    .B2(_2652_),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _5831_ (.A1(\gpio_configure[31][6] ),
    .A2(_2503_),
    .B1(_2515_),
    .B2(\gpio_configure[24][6] ),
    .X(_2653_));
 sky130_fd_sc_hd__a221o_1 _5832_ (.A1(\gpio_configure[28][6] ),
    .A2(_2521_),
    .B1(_2522_),
    .B2(\gpio_configure[5][6] ),
    .C1(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__a22o_1 _5833_ (.A1(\gpio_configure[7][6] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][6] ),
    .X(_2655_));
 sky130_fd_sc_hd__a221o_1 _5834_ (.A1(\gpio_configure[12][6] ),
    .A2(_2529_),
    .B1(_2535_),
    .B2(\gpio_configure[21][6] ),
    .C1(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__a22o_1 _5835_ (.A1(\gpio_configure[29][6] ),
    .A2(_2513_),
    .B1(_2517_),
    .B2(\gpio_configure[6][6] ),
    .X(_2657_));
 sky130_fd_sc_hd__a21o_1 _5836_ (.A1(\gpio_configure[14][6] ),
    .A2(_2519_),
    .B1(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__a22o_1 _5837_ (.A1(\gpio_configure[18][6] ),
    .A2(_2495_),
    .B1(_2509_),
    .B2(\gpio_configure[8][6] ),
    .X(_2659_));
 sky130_fd_sc_hd__a221o_1 _5838_ (.A1(\gpio_configure[13][6] ),
    .A2(_2501_),
    .B1(_2527_),
    .B2(\gpio_configure[9][6] ),
    .C1(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__or4_2 _5839_ (.A(_2654_),
    .B(_2656_),
    .C(_2658_),
    .D(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__a22o_1 _5840_ (.A1(\gpio_configure[3][6] ),
    .A2(_2502_),
    .B1(_2520_),
    .B2(\gpio_configure[27][6] ),
    .X(_2662_));
 sky130_fd_sc_hd__a221o_1 _5841_ (.A1(\gpio_configure[26][6] ),
    .A2(_2497_),
    .B1(_2531_),
    .B2(\gpio_configure[2][6] ),
    .C1(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__or2_1 _5842_ (.A(\gpio_configure[16][6] ),
    .B(net404),
    .X(_2664_));
 sky130_fd_sc_hd__a22o_2 _5843_ (.A1(\gpio_configure[25][6] ),
    .A2(_2534_),
    .B1(_2664_),
    .B2(_2524_),
    .X(_2665_));
 sky130_fd_sc_hd__a221o_1 _5844_ (.A1(\gpio_configure[22][6] ),
    .A2(_2516_),
    .B1(_2518_),
    .B2(\gpio_configure[30][6] ),
    .C1(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__a22o_1 _5845_ (.A1(\gpio_configure[19][6] ),
    .A2(_2506_),
    .B1(_2510_),
    .B2(\gpio_configure[20][6] ),
    .X(_2667_));
 sky130_fd_sc_hd__a221o_1 _5846_ (.A1(\gpio_configure[10][6] ),
    .A2(_2532_),
    .B1(_2533_),
    .B2(\gpio_configure[11][6] ),
    .C1(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__a22o_1 _5847_ (.A1(\gpio_configure[23][6] ),
    .A2(_2511_),
    .B1(_2530_),
    .B2(\gpio_configure[4][6] ),
    .X(_2669_));
 sky130_fd_sc_hd__a221o_1 _5848_ (.A1(\gpio_configure[15][6] ),
    .A2(_2504_),
    .B1(_2512_),
    .B2(\gpio_configure[17][6] ),
    .C1(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__or4_1 _5849_ (.A(_2663_),
    .B(_2666_),
    .C(_2668_),
    .D(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__o221a_2 _5850_ (.A1(\gpio_configure[0][6] ),
    .A2(_2526_),
    .B1(_2661_),
    .B2(_2671_),
    .C1(net405),
    .X(_2672_));
 sky130_fd_sc_hd__a21o_1 _5851_ (.A1(net407),
    .A2(\serial_data_staging_1[5] ),
    .B1(net353),
    .X(_2673_));
 sky130_fd_sc_hd__o22a_1 _5852_ (.A1(\serial_data_staging_1[6] ),
    .A2(net352),
    .B1(_2672_),
    .B2(_2673_),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _5853_ (.A1(\gpio_configure[8][7] ),
    .A2(_2509_),
    .B1(_2535_),
    .B2(\gpio_configure[21][7] ),
    .X(_2674_));
 sky130_fd_sc_hd__a221o_4 _5854_ (.A1(\gpio_configure[13][7] ),
    .A2(_2501_),
    .B1(_2504_),
    .B2(\gpio_configure[15][7] ),
    .C1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__a22o_1 _5855_ (.A1(\gpio_configure[20][7] ),
    .A2(_2510_),
    .B1(_2516_),
    .B2(\gpio_configure[22][7] ),
    .X(_2676_));
 sky130_fd_sc_hd__a221o_1 _5856_ (.A1(\gpio_configure[30][7] ),
    .A2(_2518_),
    .B1(_2532_),
    .B2(\gpio_configure[10][7] ),
    .C1(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__a22o_1 _5857_ (.A1(\gpio_configure[31][7] ),
    .A2(_2503_),
    .B1(_2534_),
    .B2(\gpio_configure[25][7] ),
    .X(_2678_));
 sky130_fd_sc_hd__a21o_1 _5858_ (.A1(\gpio_configure[1][7] ),
    .A2(_2528_),
    .B1(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__a22o_1 _5859_ (.A1(\gpio_configure[7][7] ),
    .A2(_2508_),
    .B1(_2517_),
    .B2(\gpio_configure[6][7] ),
    .X(_2680_));
 sky130_fd_sc_hd__a221o_4 _5860_ (.A1(\gpio_configure[18][7] ),
    .A2(_2495_),
    .B1(_2530_),
    .B2(\gpio_configure[4][7] ),
    .C1(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__or4_2 _5861_ (.A(_2675_),
    .B(_2677_),
    .C(_2679_),
    .D(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__a22o_1 _5862_ (.A1(\gpio_configure[26][7] ),
    .A2(_2497_),
    .B1(_2520_),
    .B2(\gpio_configure[27][7] ),
    .X(_2683_));
 sky130_fd_sc_hd__a221o_1 _5863_ (.A1(\gpio_configure[17][7] ),
    .A2(_2512_),
    .B1(_2531_),
    .B2(\gpio_configure[2][7] ),
    .C1(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__or2_1 _5864_ (.A(\gpio_configure[16][7] ),
    .B(net404),
    .X(_2685_));
 sky130_fd_sc_hd__a22o_1 _5865_ (.A1(\gpio_configure[11][7] ),
    .A2(_2533_),
    .B1(_2685_),
    .B2(_2524_),
    .X(_2686_));
 sky130_fd_sc_hd__a221o_1 _5866_ (.A1(\gpio_configure[19][7] ),
    .A2(_2506_),
    .B1(_2511_),
    .B2(\gpio_configure[23][7] ),
    .C1(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__a22o_1 _5867_ (.A1(\gpio_configure[3][7] ),
    .A2(_2502_),
    .B1(_2515_),
    .B2(\gpio_configure[24][7] ),
    .X(_2688_));
 sky130_fd_sc_hd__a221o_1 _5868_ (.A1(\gpio_configure[28][7] ),
    .A2(_2521_),
    .B1(_2522_),
    .B2(\gpio_configure[5][7] ),
    .C1(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__a22o_1 _5869_ (.A1(\gpio_configure[29][7] ),
    .A2(_2513_),
    .B1(_2529_),
    .B2(\gpio_configure[12][7] ),
    .X(_2690_));
 sky130_fd_sc_hd__a221o_1 _5870_ (.A1(\gpio_configure[14][7] ),
    .A2(_2519_),
    .B1(_2527_),
    .B2(\gpio_configure[9][7] ),
    .C1(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__or4_2 _5871_ (.A(_2684_),
    .B(_2687_),
    .C(_2689_),
    .D(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__o221a_4 _5872_ (.A1(\gpio_configure[0][7] ),
    .A2(_2526_),
    .B1(_2682_),
    .B2(_2692_),
    .C1(net405),
    .X(_2693_));
 sky130_fd_sc_hd__a21o_1 _5873_ (.A1(net407),
    .A2(\serial_data_staging_1[6] ),
    .B1(net353),
    .X(_2694_));
 sky130_fd_sc_hd__o22a_1 _5874_ (.A1(\serial_data_staging_1[7] ),
    .A2(net352),
    .B1(_2693_),
    .B2(_2694_),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _5875_ (.A1(\gpio_configure[15][8] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][8] ),
    .X(_2695_));
 sky130_fd_sc_hd__a221o_1 _5876_ (.A1(\gpio_configure[30][8] ),
    .A2(_2518_),
    .B1(_2533_),
    .B2(\gpio_configure[11][8] ),
    .C1(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__a22o_1 _5877_ (.A1(\gpio_configure[20][8] ),
    .A2(_2510_),
    .B1(_2528_),
    .B2(\gpio_configure[1][8] ),
    .X(_2697_));
 sky130_fd_sc_hd__a221o_1 _5878_ (.A1(\gpio_configure[26][8] ),
    .A2(_2497_),
    .B1(_2506_),
    .B2(\gpio_configure[19][8] ),
    .C1(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__a22o_1 _5879_ (.A1(\gpio_configure[31][8] ),
    .A2(_2503_),
    .B1(_2511_),
    .B2(\gpio_configure[23][8] ),
    .X(_2699_));
 sky130_fd_sc_hd__a21o_1 _5880_ (.A1(\gpio_configure[18][8] ),
    .A2(_2495_),
    .B1(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__a22o_2 _5881_ (.A1(\gpio_configure[17][8] ),
    .A2(_2512_),
    .B1(_2532_),
    .B2(\gpio_configure[10][8] ),
    .X(_2701_));
 sky130_fd_sc_hd__a221o_1 _5882_ (.A1(\gpio_configure[8][8] ),
    .A2(_2509_),
    .B1(_2515_),
    .B2(\gpio_configure[24][8] ),
    .C1(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__or4_1 _5883_ (.A(_2696_),
    .B(_2698_),
    .C(_2700_),
    .D(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a22o_1 _5884_ (.A1(\gpio_configure[7][8] ),
    .A2(_2508_),
    .B1(_2513_),
    .B2(\gpio_configure[29][8] ),
    .X(_2704_));
 sky130_fd_sc_hd__a221o_1 _5885_ (.A1(\gpio_configure[5][8] ),
    .A2(_2522_),
    .B1(_2531_),
    .B2(\gpio_configure[2][8] ),
    .C1(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__or2_1 _5886_ (.A(\gpio_configure[16][8] ),
    .B(_0830_),
    .X(_2706_));
 sky130_fd_sc_hd__a22o_1 _5887_ (.A1(\gpio_configure[6][8] ),
    .A2(_2517_),
    .B1(_2524_),
    .B2(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__a221o_2 _5888_ (.A1(\gpio_configure[9][8] ),
    .A2(_2527_),
    .B1(_2534_),
    .B2(\gpio_configure[25][8] ),
    .C1(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__a22o_1 _5889_ (.A1(\gpio_configure[14][8] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][8] ),
    .X(_2709_));
 sky130_fd_sc_hd__a221o_1 _5890_ (.A1(\gpio_configure[13][8] ),
    .A2(_2501_),
    .B1(_2521_),
    .B2(\gpio_configure[28][8] ),
    .C1(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__a22o_1 _5891_ (.A1(\gpio_configure[3][8] ),
    .A2(_2502_),
    .B1(_2535_),
    .B2(\gpio_configure[21][8] ),
    .X(_2711_));
 sky130_fd_sc_hd__a221o_1 _5892_ (.A1(\gpio_configure[22][8] ),
    .A2(_2516_),
    .B1(_2520_),
    .B2(\gpio_configure[27][8] ),
    .C1(_2711_),
    .X(_2712_));
 sky130_fd_sc_hd__or4_2 _5893_ (.A(_2705_),
    .B(_2708_),
    .C(_2710_),
    .D(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__o221a_4 _5894_ (.A1(\gpio_configure[0][8] ),
    .A2(_2526_),
    .B1(_2703_),
    .B2(_2713_),
    .C1(net405),
    .X(_2714_));
 sky130_fd_sc_hd__a211o_1 _5895_ (.A1(net408),
    .A2(\serial_data_staging_1[7] ),
    .B1(net353),
    .C1(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__o21a_1 _5896_ (.A1(\serial_data_staging_1[8] ),
    .A2(net352),
    .B1(_2715_),
    .X(_0772_));
 sky130_fd_sc_hd__a22o_1 _5897_ (.A1(\gpio_configure[29][9] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][9] ),
    .X(_2716_));
 sky130_fd_sc_hd__a22o_1 _5898_ (.A1(\gpio_configure[11][9] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][9] ),
    .X(_2717_));
 sky130_fd_sc_hd__or2_1 _5899_ (.A(\gpio_configure[16][9] ),
    .B(_0830_),
    .X(_2718_));
 sky130_fd_sc_hd__a221o_1 _5900_ (.A1(\gpio_configure[19][9] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][9] ),
    .C1(_2717_),
    .X(_2719_));
 sky130_fd_sc_hd__a22o_2 _5901_ (.A1(\gpio_configure[5][9] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][9] ),
    .X(_2720_));
 sky130_fd_sc_hd__a22o_1 _5902_ (.A1(\gpio_configure[18][9] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][9] ),
    .X(_2721_));
 sky130_fd_sc_hd__a221o_1 _5903_ (.A1(\gpio_configure[23][9] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][9] ),
    .C1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__a22o_1 _5904_ (.A1(\gpio_configure[14][9] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][9] ),
    .X(_2723_));
 sky130_fd_sc_hd__a221o_2 _5905_ (.A1(\gpio_configure[13][9] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][9] ),
    .C1(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__a22o_1 _5906_ (.A1(\gpio_configure[3][9] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][9] ),
    .X(_2725_));
 sky130_fd_sc_hd__a221o_1 _5907_ (.A1(\gpio_configure[31][9] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][9] ),
    .C1(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__a22o_1 _5908_ (.A1(\gpio_configure[26][9] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(_2718_),
    .X(_2727_));
 sky130_fd_sc_hd__a221o_1 _5909_ (.A1(\gpio_configure[15][9] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][9] ),
    .C1(_2727_),
    .X(_2728_));
 sky130_fd_sc_hd__or4_2 _5910_ (.A(_2722_),
    .B(_2724_),
    .C(_2726_),
    .D(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__a221o_1 _5911_ (.A1(\gpio_configure[7][9] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][9] ),
    .C1(_2716_),
    .X(_2730_));
 sky130_fd_sc_hd__a211o_1 _5912_ (.A1(\gpio_configure[6][9] ),
    .A2(_2517_),
    .B1(_2720_),
    .C1(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__a22o_1 _5913_ (.A1(\gpio_configure[20][9] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][9] ),
    .X(_2732_));
 sky130_fd_sc_hd__a221o_1 _5914_ (.A1(\gpio_configure[30][9] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][9] ),
    .C1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__or4_2 _5915_ (.A(_2719_),
    .B(_2729_),
    .C(_2731_),
    .D(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__o211a_1 _5916_ (.A1(\gpio_configure[0][9] ),
    .A2(_2526_),
    .B1(_2734_),
    .C1(net405),
    .X(_2735_));
 sky130_fd_sc_hd__a211o_1 _5917_ (.A1(net408),
    .A2(\serial_data_staging_1[8] ),
    .B1(net353),
    .C1(_2735_),
    .X(_2736_));
 sky130_fd_sc_hd__o21a_1 _5918_ (.A1(\serial_data_staging_1[9] ),
    .A2(net352),
    .B1(_2736_),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _5919_ (.A1(\gpio_configure[4][10] ),
    .A2(_2530_),
    .B1(_2533_),
    .B2(\gpio_configure[11][10] ),
    .X(_2737_));
 sky130_fd_sc_hd__a221o_1 _5920_ (.A1(\gpio_configure[6][10] ),
    .A2(_2517_),
    .B1(_2522_),
    .B2(\gpio_configure[5][10] ),
    .C1(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__a22o_1 _5921_ (.A1(\gpio_configure[26][10] ),
    .A2(_2497_),
    .B1(_2512_),
    .B2(\gpio_configure[17][10] ),
    .X(_2739_));
 sky130_fd_sc_hd__a221o_1 _5922_ (.A1(\gpio_configure[15][10] ),
    .A2(_2504_),
    .B1(_2510_),
    .B2(\gpio_configure[20][10] ),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__a22o_1 _5923_ (.A1(\gpio_configure[7][10] ),
    .A2(_2508_),
    .B1(_2515_),
    .B2(\gpio_configure[24][10] ),
    .X(_2741_));
 sky130_fd_sc_hd__a21o_1 _5924_ (.A1(\gpio_configure[8][10] ),
    .A2(_2509_),
    .B1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__a22o_1 _5925_ (.A1(\gpio_configure[1][10] ),
    .A2(_2528_),
    .B1(_2529_),
    .B2(\gpio_configure[12][10] ),
    .X(_2743_));
 sky130_fd_sc_hd__a221o_1 _5926_ (.A1(\gpio_configure[30][10] ),
    .A2(_2518_),
    .B1(_2527_),
    .B2(\gpio_configure[9][10] ),
    .C1(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__or4_4 _5927_ (.A(_2738_),
    .B(_2740_),
    .C(_2742_),
    .D(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__a22o_1 _5928_ (.A1(\gpio_configure[31][10] ),
    .A2(_2503_),
    .B1(_2511_),
    .B2(\gpio_configure[23][10] ),
    .X(_2746_));
 sky130_fd_sc_hd__a221o_1 _5929_ (.A1(\gpio_configure[29][10] ),
    .A2(_2513_),
    .B1(_2534_),
    .B2(\gpio_configure[25][10] ),
    .C1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__or2_1 _5930_ (.A(\gpio_configure[16][10] ),
    .B(_0830_),
    .X(_2748_));
 sky130_fd_sc_hd__a22o_4 _5931_ (.A1(\gpio_configure[2][10] ),
    .A2(_2531_),
    .B1(_2748_),
    .B2(_2524_),
    .X(_2749_));
 sky130_fd_sc_hd__a221o_1 _5932_ (.A1(\gpio_configure[28][10] ),
    .A2(_2521_),
    .B1(_2535_),
    .B2(\gpio_configure[21][10] ),
    .C1(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__a22o_1 _5933_ (.A1(\gpio_configure[14][10] ),
    .A2(_2519_),
    .B1(_2532_),
    .B2(\gpio_configure[10][10] ),
    .X(_2751_));
 sky130_fd_sc_hd__a221o_4 _5934_ (.A1(\gpio_configure[13][10] ),
    .A2(_2501_),
    .B1(_2502_),
    .B2(\gpio_configure[3][10] ),
    .C1(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__a22o_1 _5935_ (.A1(\gpio_configure[19][10] ),
    .A2(_2506_),
    .B1(_2516_),
    .B2(\gpio_configure[22][10] ),
    .X(_2753_));
 sky130_fd_sc_hd__a221o_1 _5936_ (.A1(\gpio_configure[18][10] ),
    .A2(_2495_),
    .B1(_2520_),
    .B2(\gpio_configure[27][10] ),
    .C1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__or4_1 _5937_ (.A(_2747_),
    .B(_2750_),
    .C(_2752_),
    .D(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__o221a_4 _5938_ (.A1(\gpio_configure[0][10] ),
    .A2(_2526_),
    .B1(_2745_),
    .B2(_2755_),
    .C1(net405),
    .X(_2756_));
 sky130_fd_sc_hd__a21o_1 _5939_ (.A1(net408),
    .A2(\serial_data_staging_1[9] ),
    .B1(net353),
    .X(_2757_));
 sky130_fd_sc_hd__o22a_1 _5940_ (.A1(\serial_data_staging_1[10] ),
    .A2(net352),
    .B1(_2756_),
    .B2(_2757_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _5941_ (.A1(\gpio_configure[7][11] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][11] ),
    .X(_2758_));
 sky130_fd_sc_hd__or2_1 _5942_ (.A(\gpio_configure[16][11] ),
    .B(_0830_),
    .X(_2759_));
 sky130_fd_sc_hd__a22o_2 _5943_ (.A1(\gpio_configure[5][11] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][11] ),
    .X(_2760_));
 sky130_fd_sc_hd__a22o_1 _5944_ (.A1(\gpio_configure[29][11] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][11] ),
    .X(_2761_));
 sky130_fd_sc_hd__a22o_1 _5945_ (.A1(\gpio_configure[18][11] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][11] ),
    .X(_2762_));
 sky130_fd_sc_hd__a221o_1 _5946_ (.A1(\gpio_configure[23][11] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][11] ),
    .C1(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__a22o_1 _5947_ (.A1(\gpio_configure[14][11] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][11] ),
    .X(_2764_));
 sky130_fd_sc_hd__a221o_2 _5948_ (.A1(\gpio_configure[13][11] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][11] ),
    .C1(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__a22o_1 _5949_ (.A1(\gpio_configure[3][11] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][11] ),
    .X(_2766_));
 sky130_fd_sc_hd__a221o_1 _5950_ (.A1(\gpio_configure[31][11] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][11] ),
    .C1(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__a22o_1 _5951_ (.A1(\gpio_configure[26][11] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(_2759_),
    .X(_2768_));
 sky130_fd_sc_hd__a221o_2 _5952_ (.A1(\gpio_configure[15][11] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][11] ),
    .C1(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__or4_2 _5953_ (.A(_2763_),
    .B(_2765_),
    .C(_2767_),
    .D(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__a211o_2 _5954_ (.A1(\gpio_configure[6][11] ),
    .A2(_2517_),
    .B1(_2758_),
    .C1(_2761_),
    .X(_2771_));
 sky130_fd_sc_hd__a22o_1 _5955_ (.A1(\gpio_configure[20][11] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][11] ),
    .X(_2772_));
 sky130_fd_sc_hd__a221o_1 _5956_ (.A1(\gpio_configure[30][11] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][11] ),
    .C1(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__a22o_1 _5957_ (.A1(\gpio_configure[19][11] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][11] ),
    .X(_2774_));
 sky130_fd_sc_hd__a221o_1 _5958_ (.A1(\gpio_configure[11][11] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][11] ),
    .C1(_2774_),
    .X(_2775_));
 sky130_fd_sc_hd__or4_1 _5959_ (.A(_2760_),
    .B(_2771_),
    .C(_2773_),
    .D(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__o221a_4 _5960_ (.A1(\gpio_configure[0][11] ),
    .A2(_2526_),
    .B1(_2770_),
    .B2(_2776_),
    .C1(net405),
    .X(_2777_));
 sky130_fd_sc_hd__a211o_1 _5961_ (.A1(net408),
    .A2(\serial_data_staging_1[10] ),
    .B1(net353),
    .C1(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__o21a_1 _5962_ (.A1(\serial_data_staging_1[11] ),
    .A2(net352),
    .B1(_2778_),
    .X(_0775_));
 sky130_fd_sc_hd__or2_1 _5963_ (.A(\gpio_configure[16][12] ),
    .B(_0830_),
    .X(_2779_));
 sky130_fd_sc_hd__a22o_1 _5964_ (.A1(\gpio_configure[29][12] ),
    .A2(_2513_),
    .B1(_2527_),
    .B2(\gpio_configure[9][12] ),
    .X(_2780_));
 sky130_fd_sc_hd__a22o_1 _5965_ (.A1(\gpio_configure[19][12] ),
    .A2(_2506_),
    .B1(_2520_),
    .B2(\gpio_configure[27][12] ),
    .X(_2781_));
 sky130_fd_sc_hd__a22o_1 _5966_ (.A1(\gpio_configure[11][12] ),
    .A2(_2533_),
    .B1(_2535_),
    .B2(\gpio_configure[21][12] ),
    .X(_2782_));
 sky130_fd_sc_hd__a22o_1 _5967_ (.A1(\gpio_configure[5][12] ),
    .A2(_2522_),
    .B1(_2534_),
    .B2(\gpio_configure[25][12] ),
    .X(_2783_));
 sky130_fd_sc_hd__a22o_1 _5968_ (.A1(\gpio_configure[18][12] ),
    .A2(_2495_),
    .B1(_2515_),
    .B2(\gpio_configure[24][12] ),
    .X(_2784_));
 sky130_fd_sc_hd__a221o_1 _5969_ (.A1(\gpio_configure[23][12] ),
    .A2(_2511_),
    .B1(_2532_),
    .B2(\gpio_configure[10][12] ),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a22o_1 _5970_ (.A1(\gpio_configure[14][12] ),
    .A2(_2519_),
    .B1(_2529_),
    .B2(\gpio_configure[12][12] ),
    .X(_2786_));
 sky130_fd_sc_hd__a221o_2 _5971_ (.A1(\gpio_configure[13][12] ),
    .A2(_2501_),
    .B1(_2509_),
    .B2(\gpio_configure[8][12] ),
    .C1(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__a22o_1 _5972_ (.A1(\gpio_configure[3][12] ),
    .A2(_2502_),
    .B1(_2516_),
    .B2(\gpio_configure[22][12] ),
    .X(_2788_));
 sky130_fd_sc_hd__a221o_1 _5973_ (.A1(\gpio_configure[31][12] ),
    .A2(_2503_),
    .B1(_2512_),
    .B2(\gpio_configure[17][12] ),
    .C1(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__a22o_1 _5974_ (.A1(\gpio_configure[26][12] ),
    .A2(_2497_),
    .B1(_2524_),
    .B2(_2779_),
    .X(_2790_));
 sky130_fd_sc_hd__a221o_2 _5975_ (.A1(\gpio_configure[15][12] ),
    .A2(_2504_),
    .B1(_2530_),
    .B2(\gpio_configure[4][12] ),
    .C1(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__or4_2 _5976_ (.A(_2785_),
    .B(_2787_),
    .C(_2789_),
    .D(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__a221o_1 _5977_ (.A1(\gpio_configure[7][12] ),
    .A2(_2508_),
    .B1(_2528_),
    .B2(\gpio_configure[1][12] ),
    .C1(_2780_),
    .X(_2793_));
 sky130_fd_sc_hd__a211o_1 _5978_ (.A1(\gpio_configure[6][12] ),
    .A2(_2517_),
    .B1(_2783_),
    .C1(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__a22o_1 _5979_ (.A1(\gpio_configure[20][12] ),
    .A2(_2510_),
    .B1(_2531_),
    .B2(\gpio_configure[2][12] ),
    .X(_2795_));
 sky130_fd_sc_hd__a221o_1 _5980_ (.A1(\gpio_configure[30][12] ),
    .A2(_2518_),
    .B1(_2521_),
    .B2(\gpio_configure[28][12] ),
    .C1(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__or4_1 _5981_ (.A(_2781_),
    .B(_2782_),
    .C(_2794_),
    .D(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__o221a_4 _5982_ (.A1(\gpio_configure[0][12] ),
    .A2(_2526_),
    .B1(_2792_),
    .B2(_2797_),
    .C1(net405),
    .X(_2798_));
 sky130_fd_sc_hd__a21o_1 _5983_ (.A1(net408),
    .A2(\serial_data_staging_1[11] ),
    .B1(net353),
    .X(_2799_));
 sky130_fd_sc_hd__o22a_1 _5984_ (.A1(\serial_data_staging_1[12] ),
    .A2(net352),
    .B1(_2798_),
    .B2(_2799_),
    .X(_0776_));
 sky130_fd_sc_hd__nor2_8 _5985_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .Y(_2800_));
 sky130_fd_sc_hd__nand2_8 _5986_ (.A(_1444_),
    .B(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__nor2_8 _5987_ (.A(_2484_),
    .B(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__nor2_8 _5988_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_2803_));
 sky130_fd_sc_hd__or2_4 _5989_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .X(_2804_));
 sky130_fd_sc_hd__nor2_8 _5990_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .Y(_2805_));
 sky130_fd_sc_hd__nand2_8 _5991_ (.A(_1445_),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__nor2_8 _5992_ (.A(_2804_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__and3b_4 _5993_ (.A_N(_1443_),
    .B(_2800_),
    .C(_2805_),
    .X(_2808_));
 sky130_fd_sc_hd__nor2_8 _5994_ (.A(_1446_),
    .B(_2804_),
    .Y(_2809_));
 sky130_fd_sc_hd__and2b_4 _5995_ (.A_N(\pad_count_2[2] ),
    .B(\pad_count_2[3] ),
    .X(_2810_));
 sky130_fd_sc_hd__and3_4 _5996_ (.A(_1444_),
    .B(_2483_),
    .C(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__and3_4 _5997_ (.A(_1444_),
    .B(_2803_),
    .C(_2810_),
    .X(_2812_));
 sky130_fd_sc_hd__and3b_4 _5998_ (.A_N(_1443_),
    .B(_2474_),
    .C(_2800_),
    .X(_2813_));
 sky130_fd_sc_hd__nor2_8 _5999_ (.A(_1443_),
    .B(_2801_),
    .Y(_2814_));
 sky130_fd_sc_hd__and3_4 _6000_ (.A(_2474_),
    .B(_2478_),
    .C(_2803_),
    .X(_2815_));
 sky130_fd_sc_hd__nand2_8 _6001_ (.A(_1445_),
    .B(_2476_),
    .Y(_2816_));
 sky130_fd_sc_hd__nor2_8 _6002_ (.A(_1443_),
    .B(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__and3_4 _6003_ (.A(_2474_),
    .B(_2800_),
    .C(_2803_),
    .X(_2818_));
 sky130_fd_sc_hd__nor2_8 _6004_ (.A(_2801_),
    .B(_2804_),
    .Y(_2819_));
 sky130_fd_sc_hd__nor2_8 _6005_ (.A(_2804_),
    .B(_2816_),
    .Y(_2820_));
 sky130_fd_sc_hd__and3_4 _6006_ (.A(_2478_),
    .B(_2803_),
    .C(_2805_),
    .X(_2821_));
 sky130_fd_sc_hd__and3_4 _6007_ (.A(_2476_),
    .B(_2803_),
    .C(_2810_),
    .X(_2822_));
 sky130_fd_sc_hd__and3_4 _6008_ (.A(_1445_),
    .B(_2474_),
    .C(_2803_),
    .X(_2823_));
 sky130_fd_sc_hd__and3_4 _6009_ (.A(_2474_),
    .B(_2483_),
    .C(_2810_),
    .X(_2824_));
 sky130_fd_sc_hd__nor2_8 _6010_ (.A(_2484_),
    .B(_2816_),
    .Y(_2825_));
 sky130_fd_sc_hd__and3_4 _6011_ (.A(_1444_),
    .B(_2478_),
    .C(_2483_),
    .X(_2826_));
 sky130_fd_sc_hd__and3_4 _6012_ (.A(_1444_),
    .B(_2478_),
    .C(_2803_),
    .X(_2827_));
 sky130_fd_sc_hd__nand2_8 _6013_ (.A(_2476_),
    .B(_2800_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_8 _6014_ (.A(_2804_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__and3_4 _6015_ (.A(_2474_),
    .B(_2803_),
    .C(_2810_),
    .X(_2830_));
 sky130_fd_sc_hd__and3_4 _6016_ (.A(_2476_),
    .B(_2478_),
    .C(_2803_),
    .X(_2831_));
 sky130_fd_sc_hd__nor2_8 _6017_ (.A(_1443_),
    .B(_2828_),
    .Y(_2832_));
 sky130_fd_sc_hd__and3_4 _6018_ (.A(_2803_),
    .B(_2805_),
    .C(_2810_),
    .X(_2833_));
 sky130_fd_sc_hd__nor2_8 _6019_ (.A(_1443_),
    .B(_2806_),
    .Y(_2834_));
 sky130_fd_sc_hd__or4_1 _6020_ (.A(_2807_),
    .B(_2813_),
    .C(_2823_),
    .D(_2827_),
    .X(_2835_));
 sky130_fd_sc_hd__or4_1 _6021_ (.A(_2809_),
    .B(_2817_),
    .C(_2818_),
    .D(_2834_),
    .X(_2836_));
 sky130_fd_sc_hd__or4_1 _6022_ (.A(_2821_),
    .B(_2830_),
    .C(_2831_),
    .D(_2833_),
    .X(_2837_));
 sky130_fd_sc_hd__or4_1 _6023_ (.A(_2814_),
    .B(_2815_),
    .C(_2819_),
    .D(_2832_),
    .X(_2838_));
 sky130_fd_sc_hd__or4_4 _6024_ (.A(_2835_),
    .B(_2836_),
    .C(_2837_),
    .D(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__or4_4 _6025_ (.A(_2812_),
    .B(_2820_),
    .C(_2822_),
    .D(_2829_),
    .X(_2840_));
 sky130_fd_sc_hd__nor4_4 _6026_ (.A(_2483_),
    .B(_2808_),
    .C(_2839_),
    .D(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__or4_4 _6027_ (.A(_2483_),
    .B(_2808_),
    .C(_2839_),
    .D(_2840_),
    .X(_2842_));
 sky130_fd_sc_hd__and3_4 _6028_ (.A(_2483_),
    .B(_2800_),
    .C(_2805_),
    .X(_2843_));
 sky130_fd_sc_hd__and3_4 _6029_ (.A(_2483_),
    .B(_2805_),
    .C(_2810_),
    .X(_2844_));
 sky130_fd_sc_hd__nor2_8 _6030_ (.A(_1446_),
    .B(_2484_),
    .Y(_2845_));
 sky130_fd_sc_hd__and3_4 _6031_ (.A(_2476_),
    .B(_2478_),
    .C(_2483_),
    .X(_2846_));
 sky130_fd_sc_hd__and3_4 _6032_ (.A(_2476_),
    .B(_2483_),
    .C(_2810_),
    .X(_2847_));
 sky130_fd_sc_hd__and3_4 _6033_ (.A(_2474_),
    .B(_2483_),
    .C(_2800_),
    .X(_2848_));
 sky130_fd_sc_hd__nor2_8 _6034_ (.A(_2484_),
    .B(_2828_),
    .Y(_2849_));
 sky130_fd_sc_hd__and3_4 _6035_ (.A(_2478_),
    .B(_2483_),
    .C(_2805_),
    .X(_2850_));
 sky130_fd_sc_hd__nor2_8 _6036_ (.A(_2484_),
    .B(_2806_),
    .Y(_2851_));
 sky130_fd_sc_hd__and3_4 _6037_ (.A(_1445_),
    .B(_2474_),
    .C(_2483_),
    .X(_2852_));
 sky130_fd_sc_hd__a22o_1 _6038_ (.A1(\gpio_configure[30][0] ),
    .A2(_2826_),
    .B1(_2846_),
    .B2(\gpio_configure[29][0] ),
    .X(_2853_));
 sky130_fd_sc_hd__a22o_1 _6039_ (.A1(\gpio_configure[3][0] ),
    .A2(_2818_),
    .B1(_2831_),
    .B2(\gpio_configure[13][0] ),
    .X(_2854_));
 sky130_fd_sc_hd__a221o_1 _6040_ (.A1(\gpio_configure[5][0] ),
    .A2(_2820_),
    .B1(_2829_),
    .B2(\gpio_configure[1][0] ),
    .C1(_2853_),
    .X(_2855_));
 sky130_fd_sc_hd__a211o_1 _6041_ (.A1(\gpio_configure[32][0] ),
    .A2(_2808_),
    .B1(_2854_),
    .C1(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a22o_1 _6042_ (.A1(\gpio_configure[31][0] ),
    .A2(_2485_),
    .B1(_2843_),
    .B2(\gpio_configure[16][0] ),
    .X(_2857_));
 sky130_fd_sc_hd__a221o_1 _6043_ (.A1(\gpio_configure[18][0] ),
    .A2(_2802_),
    .B1(_2851_),
    .B2(\gpio_configure[20][0] ),
    .C1(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__a22o_1 _6044_ (.A1(\gpio_configure[8][0] ),
    .A2(_2833_),
    .B1(_2847_),
    .B2(\gpio_configure[25][0] ),
    .X(_2859_));
 sky130_fd_sc_hd__a221o_4 _6045_ (.A1(\gpio_configure[33][0] ),
    .A2(_2832_),
    .B1(_2849_),
    .B2(\gpio_configure[17][0] ),
    .C1(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__a22o_1 _6046_ (.A1(\gpio_configure[11][0] ),
    .A2(_2830_),
    .B1(_2848_),
    .B2(\gpio_configure[19][0] ),
    .X(_2861_));
 sky130_fd_sc_hd__a221o_2 _6047_ (.A1(\gpio_configure[28][0] ),
    .A2(_2850_),
    .B1(_2852_),
    .B2(\gpio_configure[23][0] ),
    .C1(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__a221o_1 _6048_ (.A1(\gpio_configure[4][0] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][0] ),
    .C1(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__a22o_2 _6049_ (.A1(\gpio_configure[26][0] ),
    .A2(_2811_),
    .B1(_2844_),
    .B2(\gpio_configure[24][0] ),
    .X(_2864_));
 sky130_fd_sc_hd__a221o_1 _6050_ (.A1(\gpio_configure[35][0] ),
    .A2(_2813_),
    .B1(_2815_),
    .B2(\gpio_configure[15][0] ),
    .C1(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__a22o_1 _6051_ (.A1(\gpio_configure[34][0] ),
    .A2(_2814_),
    .B1(_2827_),
    .B2(\gpio_configure[14][0] ),
    .X(_2866_));
 sky130_fd_sc_hd__a221o_1 _6052_ (.A1(\gpio_configure[6][0] ),
    .A2(_2809_),
    .B1(_2817_),
    .B2(\gpio_configure[37][0] ),
    .C1(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__a22o_1 _6053_ (.A1(\gpio_configure[12][0] ),
    .A2(_2821_),
    .B1(_2824_),
    .B2(\gpio_configure[27][0] ),
    .X(_2868_));
 sky130_fd_sc_hd__a221o_2 _6054_ (.A1(\gpio_configure[9][0] ),
    .A2(_2822_),
    .B1(_2825_),
    .B2(\gpio_configure[21][0] ),
    .C1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__a22o_1 _6055_ (.A1(\gpio_configure[7][0] ),
    .A2(_2823_),
    .B1(_2845_),
    .B2(\gpio_configure[22][0] ),
    .X(_2870_));
 sky130_fd_sc_hd__a221o_1 _6056_ (.A1(\gpio_configure[10][0] ),
    .A2(_2812_),
    .B1(_2819_),
    .B2(\gpio_configure[2][0] ),
    .C1(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__or4_1 _6057_ (.A(_2865_),
    .B(_2867_),
    .C(_2869_),
    .D(_2871_),
    .X(_2872_));
 sky130_fd_sc_hd__or3_1 _6058_ (.A(net351),
    .B(_2863_),
    .C(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__or4_4 _6059_ (.A(_2856_),
    .B(_2858_),
    .C(_2860_),
    .D(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__or2_1 _6060_ (.A(\gpio_configure[0][0] ),
    .B(_2842_),
    .X(_2875_));
 sky130_fd_sc_hd__a32o_1 _6061_ (.A1(_2491_),
    .A2(_2874_),
    .A3(_2875_),
    .B1(net353),
    .B2(\serial_data_staging_2[0] ),
    .X(_0777_));
 sky130_fd_sc_hd__a22o_1 _6062_ (.A1(\gpio_configure[32][1] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][1] ),
    .X(_2876_));
 sky130_fd_sc_hd__and2_1 _6063_ (.A(\gpio_configure[28][1] ),
    .B(_2850_),
    .X(_2877_));
 sky130_fd_sc_hd__a22o_1 _6064_ (.A1(\gpio_configure[35][1] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][1] ),
    .X(_2878_));
 sky130_fd_sc_hd__a221o_1 _6065_ (.A1(\gpio_configure[21][1] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][1] ),
    .C1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a221o_1 _6066_ (.A1(\gpio_configure[20][1] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][1] ),
    .C1(_2877_),
    .X(_2880_));
 sky130_fd_sc_hd__a22o_1 _6067_ (.A1(\gpio_configure[33][1] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][1] ),
    .X(_2881_));
 sky130_fd_sc_hd__a221o_1 _6068_ (.A1(\gpio_configure[18][1] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][1] ),
    .C1(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__a22o_1 _6069_ (.A1(\gpio_configure[27][1] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][1] ),
    .X(_2883_));
 sky130_fd_sc_hd__a221o_2 _6070_ (.A1(\gpio_configure[16][1] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][1] ),
    .C1(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__or4_1 _6071_ (.A(_2879_),
    .B(_2880_),
    .C(_2882_),
    .D(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__a221o_4 _6072_ (.A1(\gpio_configure[4][1] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][1] ),
    .C1(_2876_),
    .X(_2886_));
 sky130_fd_sc_hd__a221o_1 _6073_ (.A1(\gpio_configure[34][1] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][1] ),
    .C1(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__a22o_1 _6074_ (.A1(\gpio_configure[12][1] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][1] ),
    .X(_2888_));
 sky130_fd_sc_hd__a221o_1 _6075_ (.A1(\gpio_configure[6][1] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][1] ),
    .C1(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__a22o_1 _6076_ (.A1(\gpio_configure[13][1] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][1] ),
    .X(_2890_));
 sky130_fd_sc_hd__a221o_1 _6077_ (.A1(\gpio_configure[2][1] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][1] ),
    .C1(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__a22o_2 _6078_ (.A1(\gpio_configure[31][1] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][1] ),
    .X(_2892_));
 sky130_fd_sc_hd__a221o_4 _6079_ (.A1(\gpio_configure[1][1] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][1] ),
    .C1(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a22o_1 _6080_ (.A1(\gpio_configure[15][1] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][1] ),
    .X(_2894_));
 sky130_fd_sc_hd__a221o_1 _6081_ (.A1(\gpio_configure[26][1] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][1] ),
    .C1(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__or4_4 _6082_ (.A(_2889_),
    .B(_2891_),
    .C(_2893_),
    .D(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__or3_1 _6083_ (.A(_2841_),
    .B(_2887_),
    .C(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__o221a_2 _6084_ (.A1(\gpio_configure[0][1] ),
    .A2(_2842_),
    .B1(_2885_),
    .B2(_2897_),
    .C1(_0819_),
    .X(_2898_));
 sky130_fd_sc_hd__a21o_1 _6085_ (.A1(net407),
    .A2(\serial_data_staging_2[0] ),
    .B1(net353),
    .X(_2899_));
 sky130_fd_sc_hd__o22a_1 _6086_ (.A1(\serial_data_staging_2[1] ),
    .A2(net352),
    .B1(_2898_),
    .B2(_2899_),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _6087_ (.A1(\gpio_configure[26][2] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][2] ),
    .X(_2900_));
 sky130_fd_sc_hd__a22o_1 _6088_ (.A1(\gpio_configure[35][2] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][2] ),
    .X(_2901_));
 sky130_fd_sc_hd__a221o_1 _6089_ (.A1(\gpio_configure[15][2] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][2] ),
    .C1(_2900_),
    .X(_2902_));
 sky130_fd_sc_hd__a221o_1 _6090_ (.A1(\gpio_configure[21][2] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][2] ),
    .C1(_2901_),
    .X(_2903_));
 sky130_fd_sc_hd__a22o_1 _6091_ (.A1(\gpio_configure[20][2] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][2] ),
    .X(_2904_));
 sky130_fd_sc_hd__a22o_1 _6092_ (.A1(\gpio_configure[18][2] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][2] ),
    .X(_2905_));
 sky130_fd_sc_hd__a221o_1 _6093_ (.A1(\gpio_configure[33][2] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][2] ),
    .C1(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__a22o_1 _6094_ (.A1(\gpio_configure[27][2] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][2] ),
    .X(_2907_));
 sky130_fd_sc_hd__a221o_1 _6095_ (.A1(\gpio_configure[16][2] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][2] ),
    .C1(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__a2111o_1 _6096_ (.A1(\gpio_configure[28][2] ),
    .A2(_2850_),
    .B1(_2904_),
    .C1(_2906_),
    .D1(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__a22o_1 _6097_ (.A1(\gpio_configure[32][2] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][2] ),
    .X(_2910_));
 sky130_fd_sc_hd__a221o_2 _6098_ (.A1(\gpio_configure[4][2] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][2] ),
    .C1(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__a221o_1 _6099_ (.A1(\gpio_configure[34][2] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][2] ),
    .C1(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__a22o_1 _6100_ (.A1(\gpio_configure[12][2] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][2] ),
    .X(_2913_));
 sky130_fd_sc_hd__a221o_1 _6101_ (.A1(\gpio_configure[6][2] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][2] ),
    .C1(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a22o_1 _6102_ (.A1(\gpio_configure[13][2] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][2] ),
    .X(_2915_));
 sky130_fd_sc_hd__a221o_1 _6103_ (.A1(\gpio_configure[2][2] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][2] ),
    .C1(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__a22o_1 _6104_ (.A1(\gpio_configure[31][2] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][2] ),
    .X(_2917_));
 sky130_fd_sc_hd__a221o_1 _6105_ (.A1(\gpio_configure[1][2] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][2] ),
    .C1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__or4_1 _6106_ (.A(_2902_),
    .B(_2914_),
    .C(_2916_),
    .D(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__or3_4 _6107_ (.A(net351),
    .B(_2912_),
    .C(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__o32a_4 _6108_ (.A1(_2903_),
    .A2(_2909_),
    .A3(_2920_),
    .B1(_2842_),
    .B2(\gpio_configure[0][2] ),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _6109_ (.A0(\serial_data_staging_2[1] ),
    .A1(_2921_),
    .S(net405),
    .X(_2922_));
 sky130_fd_sc_hd__mux2_1 _6110_ (.A0(\serial_data_staging_2[2] ),
    .A1(_2922_),
    .S(net352),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _6111_ (.A(\gpio_configure[28][3] ),
    .B(_2850_),
    .X(_2923_));
 sky130_fd_sc_hd__a22o_1 _6112_ (.A1(\gpio_configure[35][3] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][3] ),
    .X(_2924_));
 sky130_fd_sc_hd__a22o_1 _6113_ (.A1(\gpio_configure[26][3] ),
    .A2(_2811_),
    .B1(_2818_),
    .B2(\gpio_configure[3][3] ),
    .X(_2925_));
 sky130_fd_sc_hd__a22o_1 _6114_ (.A1(\gpio_configure[15][3] ),
    .A2(_2815_),
    .B1(_2823_),
    .B2(\gpio_configure[7][3] ),
    .X(_2926_));
 sky130_fd_sc_hd__a221o_1 _6115_ (.A1(\gpio_configure[21][3] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][3] ),
    .C1(_2924_),
    .X(_2927_));
 sky130_fd_sc_hd__a221o_1 _6116_ (.A1(\gpio_configure[20][3] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][3] ),
    .C1(_2923_),
    .X(_2928_));
 sky130_fd_sc_hd__a22o_1 _6117_ (.A1(\gpio_configure[18][3] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][3] ),
    .X(_2929_));
 sky130_fd_sc_hd__a221o_4 _6118_ (.A1(\gpio_configure[33][3] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][3] ),
    .C1(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__a22o_1 _6119_ (.A1(\gpio_configure[27][3] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][3] ),
    .X(_2931_));
 sky130_fd_sc_hd__a221o_2 _6120_ (.A1(\gpio_configure[16][3] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][3] ),
    .C1(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__or4_4 _6121_ (.A(_2927_),
    .B(_2928_),
    .C(_2930_),
    .D(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__a22o_1 _6122_ (.A1(\gpio_configure[32][3] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][3] ),
    .X(_2934_));
 sky130_fd_sc_hd__a221o_2 _6123_ (.A1(\gpio_configure[4][3] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][3] ),
    .C1(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__a221o_1 _6124_ (.A1(\gpio_configure[34][3] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][3] ),
    .C1(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__a22o_1 _6125_ (.A1(\gpio_configure[12][3] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][3] ),
    .X(_2937_));
 sky130_fd_sc_hd__a221o_1 _6126_ (.A1(\gpio_configure[6][3] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][3] ),
    .C1(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__a22o_1 _6127_ (.A1(\gpio_configure[13][3] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][3] ),
    .X(_2939_));
 sky130_fd_sc_hd__a221o_1 _6128_ (.A1(\gpio_configure[2][3] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][3] ),
    .C1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__a22o_1 _6129_ (.A1(\gpio_configure[31][3] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][3] ),
    .X(_2941_));
 sky130_fd_sc_hd__a221o_1 _6130_ (.A1(\gpio_configure[1][3] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][3] ),
    .C1(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__or4_1 _6131_ (.A(_2925_),
    .B(_2926_),
    .C(_2940_),
    .D(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__or4_4 _6132_ (.A(net351),
    .B(_2936_),
    .C(_2938_),
    .D(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__o221a_1 _6133_ (.A1(\gpio_configure[0][3] ),
    .A2(_2842_),
    .B1(_2933_),
    .B2(_2944_),
    .C1(_0819_),
    .X(_2945_));
 sky130_fd_sc_hd__a211o_1 _6134_ (.A1(net408),
    .A2(\serial_data_staging_2[2] ),
    .B1(net353),
    .C1(_2945_),
    .X(_2946_));
 sky130_fd_sc_hd__o21a_1 _6135_ (.A1(\serial_data_staging_2[3] ),
    .A2(net352),
    .B1(_2946_),
    .X(_0780_));
 sky130_fd_sc_hd__and2_1 _6136_ (.A(\gpio_configure[28][4] ),
    .B(_2850_),
    .X(_2947_));
 sky130_fd_sc_hd__a22o_1 _6137_ (.A1(\gpio_configure[35][4] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][4] ),
    .X(_2948_));
 sky130_fd_sc_hd__a221o_1 _6138_ (.A1(\gpio_configure[21][4] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][4] ),
    .C1(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__a221o_1 _6139_ (.A1(\gpio_configure[20][4] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][4] ),
    .C1(_2947_),
    .X(_2950_));
 sky130_fd_sc_hd__a22o_1 _6140_ (.A1(\gpio_configure[18][4] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][4] ),
    .X(_2951_));
 sky130_fd_sc_hd__a221o_4 _6141_ (.A1(\gpio_configure[33][4] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][4] ),
    .C1(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__a22o_1 _6142_ (.A1(\gpio_configure[27][4] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][4] ),
    .X(_2953_));
 sky130_fd_sc_hd__a221o_1 _6143_ (.A1(\gpio_configure[16][4] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][4] ),
    .C1(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__or4_2 _6144_ (.A(_2949_),
    .B(_2950_),
    .C(_2952_),
    .D(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__a22o_1 _6145_ (.A1(\gpio_configure[32][4] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][4] ),
    .X(_2956_));
 sky130_fd_sc_hd__a221o_4 _6146_ (.A1(\gpio_configure[4][4] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][4] ),
    .C1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__a221o_1 _6147_ (.A1(\gpio_configure[34][4] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][4] ),
    .C1(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__a22o_1 _6148_ (.A1(\gpio_configure[12][4] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][4] ),
    .X(_2959_));
 sky130_fd_sc_hd__a221o_2 _6149_ (.A1(\gpio_configure[6][4] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][4] ),
    .C1(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__a22o_1 _6150_ (.A1(\gpio_configure[13][4] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][4] ),
    .X(_2961_));
 sky130_fd_sc_hd__a221o_1 _6151_ (.A1(\gpio_configure[2][4] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][4] ),
    .C1(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__a22o_1 _6152_ (.A1(\gpio_configure[31][4] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][4] ),
    .X(_2963_));
 sky130_fd_sc_hd__a221o_1 _6153_ (.A1(\gpio_configure[1][4] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][4] ),
    .C1(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__a22o_1 _6154_ (.A1(\gpio_configure[26][4] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][4] ),
    .X(_2965_));
 sky130_fd_sc_hd__a221o_1 _6155_ (.A1(\gpio_configure[15][4] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][4] ),
    .C1(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__or4_2 _6156_ (.A(_2960_),
    .B(_2962_),
    .C(_2964_),
    .D(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__or3_2 _6157_ (.A(net350),
    .B(_2958_),
    .C(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__o221a_4 _6158_ (.A1(\gpio_configure[0][4] ),
    .A2(_2842_),
    .B1(_2955_),
    .B2(_2968_),
    .C1(net405),
    .X(_2969_));
 sky130_fd_sc_hd__a211o_1 _6159_ (.A1(net407),
    .A2(\serial_data_staging_2[3] ),
    .B1(_2492_),
    .C1(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__o21a_1 _6160_ (.A1(\serial_data_staging_2[4] ),
    .A2(_2493_),
    .B1(_2970_),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _6161_ (.A1(\gpio_configure[15][5] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][5] ),
    .X(_2971_));
 sky130_fd_sc_hd__and2_1 _6162_ (.A(\gpio_configure[28][5] ),
    .B(_2850_),
    .X(_2972_));
 sky130_fd_sc_hd__a22o_1 _6163_ (.A1(\gpio_configure[35][5] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][5] ),
    .X(_2973_));
 sky130_fd_sc_hd__a221o_1 _6164_ (.A1(\gpio_configure[21][5] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][5] ),
    .C1(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__a221o_4 _6165_ (.A1(\gpio_configure[20][5] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][5] ),
    .C1(_2972_),
    .X(_2975_));
 sky130_fd_sc_hd__a22o_1 _6166_ (.A1(\gpio_configure[18][5] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][5] ),
    .X(_2976_));
 sky130_fd_sc_hd__a221o_1 _6167_ (.A1(\gpio_configure[33][5] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][5] ),
    .C1(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__a22o_1 _6168_ (.A1(\gpio_configure[27][5] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][5] ),
    .X(_2978_));
 sky130_fd_sc_hd__a221o_1 _6169_ (.A1(\gpio_configure[16][5] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][5] ),
    .C1(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__or4_1 _6170_ (.A(_2974_),
    .B(_2975_),
    .C(_2977_),
    .D(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__a22o_1 _6171_ (.A1(\gpio_configure[32][5] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][5] ),
    .X(_2981_));
 sky130_fd_sc_hd__a221o_2 _6172_ (.A1(\gpio_configure[4][5] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][5] ),
    .C1(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__a221o_1 _6173_ (.A1(\gpio_configure[34][5] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][5] ),
    .C1(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__a22o_1 _6174_ (.A1(\gpio_configure[12][5] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][5] ),
    .X(_2984_));
 sky130_fd_sc_hd__a221o_1 _6175_ (.A1(\gpio_configure[6][5] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][5] ),
    .C1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__a22o_1 _6176_ (.A1(\gpio_configure[13][5] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][5] ),
    .X(_2986_));
 sky130_fd_sc_hd__a221o_1 _6177_ (.A1(\gpio_configure[2][5] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][5] ),
    .C1(_2986_),
    .X(_2987_));
 sky130_fd_sc_hd__a22o_4 _6178_ (.A1(\gpio_configure[31][5] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][5] ),
    .X(_2988_));
 sky130_fd_sc_hd__a221o_1 _6179_ (.A1(\gpio_configure[1][5] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][5] ),
    .C1(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__a221o_1 _6180_ (.A1(\gpio_configure[26][5] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][5] ),
    .C1(_2971_),
    .X(_2990_));
 sky130_fd_sc_hd__or4_1 _6181_ (.A(_2985_),
    .B(_2987_),
    .C(_2989_),
    .D(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__or3_4 _6182_ (.A(net351),
    .B(_2983_),
    .C(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__o221a_4 _6183_ (.A1(\gpio_configure[0][5] ),
    .A2(_2842_),
    .B1(_2980_),
    .B2(_2992_),
    .C1(_0819_),
    .X(_2993_));
 sky130_fd_sc_hd__a21o_1 _6184_ (.A1(net407),
    .A2(\serial_data_staging_2[4] ),
    .B1(_2492_),
    .X(_2994_));
 sky130_fd_sc_hd__o22a_1 _6185_ (.A1(\serial_data_staging_2[5] ),
    .A2(_2493_),
    .B1(_2993_),
    .B2(_2994_),
    .X(_0782_));
 sky130_fd_sc_hd__and2_1 _6186_ (.A(\gpio_configure[23][6] ),
    .B(_2852_),
    .X(_2995_));
 sky130_fd_sc_hd__a22o_1 _6187_ (.A1(\gpio_configure[35][6] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][6] ),
    .X(_2996_));
 sky130_fd_sc_hd__a221o_1 _6188_ (.A1(\gpio_configure[21][6] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][6] ),
    .C1(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__a221o_1 _6189_ (.A1(\gpio_configure[28][6] ),
    .A2(_2850_),
    .B1(_2851_),
    .B2(\gpio_configure[20][6] ),
    .C1(_2995_),
    .X(_2998_));
 sky130_fd_sc_hd__a22o_1 _6190_ (.A1(\gpio_configure[33][6] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][6] ),
    .X(_2999_));
 sky130_fd_sc_hd__a221o_1 _6191_ (.A1(\gpio_configure[18][6] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][6] ),
    .C1(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__a22o_1 _6192_ (.A1(\gpio_configure[27][6] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][6] ),
    .X(_3001_));
 sky130_fd_sc_hd__a221o_2 _6193_ (.A1(\gpio_configure[16][6] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][6] ),
    .C1(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__or4_1 _6194_ (.A(_2997_),
    .B(_2998_),
    .C(_3000_),
    .D(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__a22o_1 _6195_ (.A1(\gpio_configure[32][6] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][6] ),
    .X(_3004_));
 sky130_fd_sc_hd__a221o_4 _6196_ (.A1(\gpio_configure[4][6] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][6] ),
    .C1(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__a221o_1 _6197_ (.A1(\gpio_configure[34][6] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][6] ),
    .C1(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__a22o_1 _6198_ (.A1(\gpio_configure[12][6] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][6] ),
    .X(_3007_));
 sky130_fd_sc_hd__a221o_1 _6199_ (.A1(\gpio_configure[6][6] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][6] ),
    .C1(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__a22o_1 _6200_ (.A1(\gpio_configure[13][6] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][6] ),
    .X(_3009_));
 sky130_fd_sc_hd__a221o_1 _6201_ (.A1(\gpio_configure[2][6] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][6] ),
    .C1(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__a22o_1 _6202_ (.A1(\gpio_configure[31][6] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][6] ),
    .X(_3011_));
 sky130_fd_sc_hd__a221o_1 _6203_ (.A1(\gpio_configure[1][6] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][6] ),
    .C1(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__a22o_1 _6204_ (.A1(\gpio_configure[26][6] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][6] ),
    .X(_3013_));
 sky130_fd_sc_hd__a221o_1 _6205_ (.A1(\gpio_configure[15][6] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][6] ),
    .C1(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__or4_2 _6206_ (.A(_3008_),
    .B(_3010_),
    .C(_3012_),
    .D(_3014_),
    .X(_3015_));
 sky130_fd_sc_hd__or4_4 _6207_ (.A(_2841_),
    .B(_3003_),
    .C(_3006_),
    .D(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__o211a_1 _6208_ (.A1(\gpio_configure[0][6] ),
    .A2(_2842_),
    .B1(_3016_),
    .C1(net405),
    .X(_3017_));
 sky130_fd_sc_hd__a211o_1 _6209_ (.A1(net407),
    .A2(\serial_data_staging_2[5] ),
    .B1(_2492_),
    .C1(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__o21a_1 _6210_ (.A1(\serial_data_staging_2[6] ),
    .A2(_2493_),
    .B1(_3018_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _6211_ (.A(\gpio_configure[28][7] ),
    .B(_2850_),
    .X(_3019_));
 sky130_fd_sc_hd__a22o_1 _6212_ (.A1(\gpio_configure[35][7] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][7] ),
    .X(_3020_));
 sky130_fd_sc_hd__a221o_1 _6213_ (.A1(\gpio_configure[21][7] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][7] ),
    .C1(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__a221o_1 _6214_ (.A1(\gpio_configure[20][7] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][7] ),
    .C1(_3019_),
    .X(_3022_));
 sky130_fd_sc_hd__a22o_4 _6215_ (.A1(\gpio_configure[18][7] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][7] ),
    .X(_3023_));
 sky130_fd_sc_hd__a221o_1 _6216_ (.A1(\gpio_configure[33][7] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][7] ),
    .C1(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__a22o_1 _6217_ (.A1(\gpio_configure[27][7] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][7] ),
    .X(_3025_));
 sky130_fd_sc_hd__a221o_2 _6218_ (.A1(\gpio_configure[16][7] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][7] ),
    .C1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__or4_1 _6219_ (.A(_3021_),
    .B(_3022_),
    .C(_3024_),
    .D(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__a22o_1 _6220_ (.A1(\gpio_configure[32][7] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][7] ),
    .X(_3028_));
 sky130_fd_sc_hd__a221o_4 _6221_ (.A1(\gpio_configure[4][7] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][7] ),
    .C1(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__a221o_1 _6222_ (.A1(\gpio_configure[34][7] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][7] ),
    .C1(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__a22o_1 _6223_ (.A1(\gpio_configure[12][7] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][7] ),
    .X(_3031_));
 sky130_fd_sc_hd__a221o_1 _6224_ (.A1(\gpio_configure[6][7] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][7] ),
    .C1(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__a22o_1 _6225_ (.A1(\gpio_configure[13][7] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][7] ),
    .X(_3033_));
 sky130_fd_sc_hd__a221o_1 _6226_ (.A1(\gpio_configure[2][7] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][7] ),
    .C1(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__a22o_1 _6227_ (.A1(\gpio_configure[31][7] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][7] ),
    .X(_3035_));
 sky130_fd_sc_hd__a221o_4 _6228_ (.A1(\gpio_configure[1][7] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][7] ),
    .C1(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__a22o_1 _6229_ (.A1(\gpio_configure[26][7] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][7] ),
    .X(_3037_));
 sky130_fd_sc_hd__a221o_1 _6230_ (.A1(\gpio_configure[15][7] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][7] ),
    .C1(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__or4_4 _6231_ (.A(_3032_),
    .B(_3034_),
    .C(_3036_),
    .D(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__or3_1 _6232_ (.A(_2841_),
    .B(_3030_),
    .C(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__o221a_2 _6233_ (.A1(\gpio_configure[0][7] ),
    .A2(_2842_),
    .B1(_3027_),
    .B2(_3040_),
    .C1(_0819_),
    .X(_3041_));
 sky130_fd_sc_hd__a21o_1 _6234_ (.A1(net407),
    .A2(\serial_data_staging_2[6] ),
    .B1(_2492_),
    .X(_3042_));
 sky130_fd_sc_hd__o22a_1 _6235_ (.A1(\serial_data_staging_2[7] ),
    .A2(_2493_),
    .B1(_3041_),
    .B2(_3042_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _6236_ (.A1(\gpio_configure[34][8] ),
    .A2(_2814_),
    .B1(_2827_),
    .B2(\gpio_configure[14][8] ),
    .X(_3043_));
 sky130_fd_sc_hd__a22o_1 _6237_ (.A1(\gpio_configure[18][8] ),
    .A2(_2802_),
    .B1(_2830_),
    .B2(\gpio_configure[11][8] ),
    .X(_3044_));
 sky130_fd_sc_hd__a221o_1 _6238_ (.A1(\gpio_configure[5][8] ),
    .A2(_2820_),
    .B1(_2823_),
    .B2(\gpio_configure[7][8] ),
    .C1(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__a22o_1 _6239_ (.A1(\gpio_configure[26][8] ),
    .A2(_2811_),
    .B1(_2815_),
    .B2(\gpio_configure[15][8] ),
    .X(_3046_));
 sky130_fd_sc_hd__a221o_2 _6240_ (.A1(\gpio_configure[1][8] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][8] ),
    .C1(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__a22o_1 _6241_ (.A1(\gpio_configure[31][8] ),
    .A2(_2485_),
    .B1(_2850_),
    .B2(\gpio_configure[28][8] ),
    .X(_3048_));
 sky130_fd_sc_hd__a221o_1 _6242_ (.A1(\gpio_configure[6][8] ),
    .A2(_2809_),
    .B1(_2826_),
    .B2(\gpio_configure[30][8] ),
    .C1(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__a22o_1 _6243_ (.A1(\gpio_configure[10][8] ),
    .A2(_2812_),
    .B1(_2821_),
    .B2(\gpio_configure[12][8] ),
    .X(_3050_));
 sky130_fd_sc_hd__a221o_1 _6244_ (.A1(\gpio_configure[2][8] ),
    .A2(_2819_),
    .B1(_2847_),
    .B2(\gpio_configure[25][8] ),
    .C1(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__a22o_1 _6245_ (.A1(\gpio_configure[32][8] ),
    .A2(_2808_),
    .B1(_2852_),
    .B2(\gpio_configure[23][8] ),
    .X(_3052_));
 sky130_fd_sc_hd__a221o_1 _6246_ (.A1(\gpio_configure[3][8] ),
    .A2(_2818_),
    .B1(_2846_),
    .B2(\gpio_configure[29][8] ),
    .C1(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__or4_1 _6247_ (.A(_3047_),
    .B(_3049_),
    .C(_3051_),
    .D(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__or3_2 _6248_ (.A(_3043_),
    .B(_3045_),
    .C(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__a22o_1 _6249_ (.A1(\gpio_configure[35][8] ),
    .A2(_2813_),
    .B1(_2822_),
    .B2(\gpio_configure[9][8] ),
    .X(_3056_));
 sky130_fd_sc_hd__a221o_1 _6250_ (.A1(\gpio_configure[8][8] ),
    .A2(_2833_),
    .B1(_2851_),
    .B2(\gpio_configure[20][8] ),
    .C1(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__a22o_1 _6251_ (.A1(\gpio_configure[13][8] ),
    .A2(_2831_),
    .B1(_2848_),
    .B2(\gpio_configure[19][8] ),
    .X(_3058_));
 sky130_fd_sc_hd__a221o_1 _6252_ (.A1(\gpio_configure[21][8] ),
    .A2(_2825_),
    .B1(_2832_),
    .B2(\gpio_configure[33][8] ),
    .C1(_3058_),
    .X(_3059_));
 sky130_fd_sc_hd__a22o_1 _6253_ (.A1(\gpio_configure[36][8] ),
    .A2(_2834_),
    .B1(_2845_),
    .B2(\gpio_configure[22][8] ),
    .X(_3060_));
 sky130_fd_sc_hd__a22o_1 _6254_ (.A1(\gpio_configure[37][8] ),
    .A2(_2817_),
    .B1(_2843_),
    .B2(\gpio_configure[16][8] ),
    .X(_3061_));
 sky130_fd_sc_hd__a221o_4 _6255_ (.A1(\gpio_configure[4][8] ),
    .A2(_2807_),
    .B1(_2849_),
    .B2(\gpio_configure[17][8] ),
    .C1(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__a211o_1 _6256_ (.A1(\gpio_configure[27][8] ),
    .A2(_2824_),
    .B1(_3060_),
    .C1(_3062_),
    .X(_3063_));
 sky130_fd_sc_hd__or4_2 _6257_ (.A(net350),
    .B(_3057_),
    .C(_3059_),
    .D(_3063_),
    .X(_3064_));
 sky130_fd_sc_hd__o221a_4 _6258_ (.A1(\gpio_configure[0][8] ),
    .A2(_2842_),
    .B1(_3055_),
    .B2(_3064_),
    .C1(net405),
    .X(_3065_));
 sky130_fd_sc_hd__a21o_2 _6259_ (.A1(net407),
    .A2(\serial_data_staging_2[7] ),
    .B1(net353),
    .X(_3066_));
 sky130_fd_sc_hd__o22a_1 _6260_ (.A1(\serial_data_staging_2[8] ),
    .A2(net352),
    .B1(_3065_),
    .B2(_3066_),
    .X(_0785_));
 sky130_fd_sc_hd__and2_1 _6261_ (.A(\gpio_configure[28][9] ),
    .B(_2850_),
    .X(_3067_));
 sky130_fd_sc_hd__a22o_1 _6262_ (.A1(\gpio_configure[35][9] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][9] ),
    .X(_3068_));
 sky130_fd_sc_hd__a221o_1 _6263_ (.A1(\gpio_configure[21][9] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][9] ),
    .C1(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__a221o_1 _6264_ (.A1(\gpio_configure[20][9] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][9] ),
    .C1(_3067_),
    .X(_3070_));
 sky130_fd_sc_hd__a22o_1 _6265_ (.A1(\gpio_configure[18][9] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][9] ),
    .X(_3071_));
 sky130_fd_sc_hd__a221o_1 _6266_ (.A1(\gpio_configure[33][9] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][9] ),
    .C1(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__a22o_1 _6267_ (.A1(\gpio_configure[27][9] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][9] ),
    .X(_3073_));
 sky130_fd_sc_hd__a221o_2 _6268_ (.A1(\gpio_configure[16][9] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][9] ),
    .C1(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__or4_2 _6269_ (.A(_3069_),
    .B(_3070_),
    .C(_3072_),
    .D(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__a22o_1 _6270_ (.A1(\gpio_configure[4][9] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][9] ),
    .X(_3076_));
 sky130_fd_sc_hd__a221o_1 _6271_ (.A1(\gpio_configure[32][9] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][9] ),
    .C1(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__a221o_2 _6272_ (.A1(\gpio_configure[34][9] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][9] ),
    .C1(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__a22o_2 _6273_ (.A1(\gpio_configure[12][9] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][9] ),
    .X(_3079_));
 sky130_fd_sc_hd__a221o_1 _6274_ (.A1(\gpio_configure[6][9] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][9] ),
    .C1(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__a22o_1 _6275_ (.A1(\gpio_configure[13][9] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][9] ),
    .X(_3081_));
 sky130_fd_sc_hd__a221o_2 _6276_ (.A1(\gpio_configure[2][9] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][9] ),
    .C1(_3081_),
    .X(_3082_));
 sky130_fd_sc_hd__a22o_1 _6277_ (.A1(\gpio_configure[31][9] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][9] ),
    .X(_3083_));
 sky130_fd_sc_hd__a221o_1 _6278_ (.A1(\gpio_configure[1][9] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][9] ),
    .C1(_3083_),
    .X(_3084_));
 sky130_fd_sc_hd__a22o_1 _6279_ (.A1(\gpio_configure[26][9] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][9] ),
    .X(_3085_));
 sky130_fd_sc_hd__a221o_1 _6280_ (.A1(\gpio_configure[15][9] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][9] ),
    .C1(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__or4_1 _6281_ (.A(_3080_),
    .B(_3082_),
    .C(_3084_),
    .D(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__or3_2 _6282_ (.A(net350),
    .B(_3078_),
    .C(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__o221a_2 _6283_ (.A1(\gpio_configure[0][9] ),
    .A2(_2842_),
    .B1(_3075_),
    .B2(_3088_),
    .C1(net405),
    .X(_3089_));
 sky130_fd_sc_hd__a211o_1 _6284_ (.A1(net408),
    .A2(\serial_data_staging_2[8] ),
    .B1(net353),
    .C1(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__o21a_1 _6285_ (.A1(\serial_data_staging_2[9] ),
    .A2(net352),
    .B1(_3090_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _6286_ (.A1(\gpio_configure[12][10] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][10] ),
    .X(_3091_));
 sky130_fd_sc_hd__a22o_1 _6287_ (.A1(\gpio_configure[35][10] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][10] ),
    .X(_3092_));
 sky130_fd_sc_hd__a221o_2 _6288_ (.A1(\gpio_configure[21][10] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][10] ),
    .C1(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__a22o_1 _6289_ (.A1(\gpio_configure[20][10] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][10] ),
    .X(_3094_));
 sky130_fd_sc_hd__a22o_1 _6290_ (.A1(\gpio_configure[18][10] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][10] ),
    .X(_3095_));
 sky130_fd_sc_hd__a221o_1 _6291_ (.A1(\gpio_configure[33][10] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][10] ),
    .C1(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__a22o_2 _6292_ (.A1(\gpio_configure[27][10] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][10] ),
    .X(_3097_));
 sky130_fd_sc_hd__a221o_4 _6293_ (.A1(\gpio_configure[16][10] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][10] ),
    .C1(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__a2111o_1 _6294_ (.A1(\gpio_configure[28][10] ),
    .A2(_2850_),
    .B1(_3094_),
    .C1(_3096_),
    .D1(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__a22o_1 _6295_ (.A1(\gpio_configure[32][10] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][10] ),
    .X(_3100_));
 sky130_fd_sc_hd__a221o_1 _6296_ (.A1(\gpio_configure[4][10] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][10] ),
    .C1(_3100_),
    .X(_3101_));
 sky130_fd_sc_hd__a221o_2 _6297_ (.A1(\gpio_configure[34][10] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][10] ),
    .C1(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__a221o_1 _6298_ (.A1(\gpio_configure[6][10] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][10] ),
    .C1(_3091_),
    .X(_3103_));
 sky130_fd_sc_hd__a22o_1 _6299_ (.A1(\gpio_configure[13][10] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][10] ),
    .X(_3104_));
 sky130_fd_sc_hd__a221o_1 _6300_ (.A1(\gpio_configure[2][10] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][10] ),
    .C1(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__a22o_1 _6301_ (.A1(\gpio_configure[31][10] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][10] ),
    .X(_3106_));
 sky130_fd_sc_hd__a221o_1 _6302_ (.A1(\gpio_configure[1][10] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][10] ),
    .C1(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__a22o_1 _6303_ (.A1(\gpio_configure[26][10] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][10] ),
    .X(_3108_));
 sky130_fd_sc_hd__a221o_1 _6304_ (.A1(\gpio_configure[15][10] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][10] ),
    .C1(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__or4_1 _6305_ (.A(_3103_),
    .B(_3105_),
    .C(_3107_),
    .D(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__or3_4 _6306_ (.A(net351),
    .B(_3102_),
    .C(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__o32a_4 _6307_ (.A1(_3093_),
    .A2(_3099_),
    .A3(_3111_),
    .B1(_2842_),
    .B2(\gpio_configure[0][10] ),
    .X(_3112_));
 sky130_fd_sc_hd__mux2_1 _6308_ (.A0(\serial_data_staging_2[9] ),
    .A1(_3112_),
    .S(net405),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _6309_ (.A0(\serial_data_staging_2[10] ),
    .A1(_3113_),
    .S(net352),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _6310_ (.A1(\gpio_configure[13][11] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][11] ),
    .X(_3114_));
 sky130_fd_sc_hd__and2_1 _6311_ (.A(\gpio_configure[28][11] ),
    .B(_2850_),
    .X(_3115_));
 sky130_fd_sc_hd__a22o_1 _6312_ (.A1(\gpio_configure[35][11] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][11] ),
    .X(_3116_));
 sky130_fd_sc_hd__a22o_1 _6313_ (.A1(\gpio_configure[26][11] ),
    .A2(_2811_),
    .B1(_2818_),
    .B2(\gpio_configure[3][11] ),
    .X(_3117_));
 sky130_fd_sc_hd__a22o_1 _6314_ (.A1(\gpio_configure[15][11] ),
    .A2(_2815_),
    .B1(_2823_),
    .B2(\gpio_configure[7][11] ),
    .X(_3118_));
 sky130_fd_sc_hd__a221o_1 _6315_ (.A1(\gpio_configure[21][11] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][11] ),
    .C1(_3116_),
    .X(_3119_));
 sky130_fd_sc_hd__a221o_1 _6316_ (.A1(\gpio_configure[20][11] ),
    .A2(_2851_),
    .B1(_2852_),
    .B2(\gpio_configure[23][11] ),
    .C1(_3115_),
    .X(_3120_));
 sky130_fd_sc_hd__a22o_1 _6317_ (.A1(\gpio_configure[33][11] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][11] ),
    .X(_3121_));
 sky130_fd_sc_hd__a221o_1 _6318_ (.A1(\gpio_configure[18][11] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][11] ),
    .C1(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__a22o_1 _6319_ (.A1(\gpio_configure[27][11] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][11] ),
    .X(_3123_));
 sky130_fd_sc_hd__a221o_2 _6320_ (.A1(\gpio_configure[16][11] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][11] ),
    .C1(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__or4_1 _6321_ (.A(_3119_),
    .B(_3120_),
    .C(_3122_),
    .D(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__a22o_1 _6322_ (.A1(\gpio_configure[4][11] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][11] ),
    .X(_3126_));
 sky130_fd_sc_hd__a221o_1 _6323_ (.A1(\gpio_configure[32][11] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][11] ),
    .C1(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__a221o_2 _6324_ (.A1(\gpio_configure[34][11] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][11] ),
    .C1(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__a22o_1 _6325_ (.A1(\gpio_configure[12][11] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][11] ),
    .X(_3129_));
 sky130_fd_sc_hd__a221o_1 _6326_ (.A1(\gpio_configure[6][11] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][11] ),
    .C1(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__a221o_1 _6327_ (.A1(\gpio_configure[2][11] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][11] ),
    .C1(_3114_),
    .X(_3131_));
 sky130_fd_sc_hd__a22o_1 _6328_ (.A1(\gpio_configure[31][11] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][11] ),
    .X(_3132_));
 sky130_fd_sc_hd__a221o_2 _6329_ (.A1(\gpio_configure[1][11] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][11] ),
    .C1(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__or4_1 _6330_ (.A(_3117_),
    .B(_3118_),
    .C(_3131_),
    .D(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__or4_4 _6331_ (.A(net350),
    .B(_3128_),
    .C(_3130_),
    .D(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__o221a_2 _6332_ (.A1(\gpio_configure[0][11] ),
    .A2(_2842_),
    .B1(_3125_),
    .B2(_3135_),
    .C1(net405),
    .X(_3136_));
 sky130_fd_sc_hd__a211o_1 _6333_ (.A1(net408),
    .A2(\serial_data_staging_2[10] ),
    .B1(net353),
    .C1(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__o21a_1 _6334_ (.A1(\serial_data_staging_2[11] ),
    .A2(net352),
    .B1(_3137_),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _6335_ (.A(\gpio_configure[23][12] ),
    .B(_2852_),
    .X(_3138_));
 sky130_fd_sc_hd__a22o_1 _6336_ (.A1(\gpio_configure[35][12] ),
    .A2(_2813_),
    .B1(_2826_),
    .B2(\gpio_configure[30][12] ),
    .X(_3139_));
 sky130_fd_sc_hd__a221o_1 _6337_ (.A1(\gpio_configure[21][12] ),
    .A2(_2825_),
    .B1(_2846_),
    .B2(\gpio_configure[29][12] ),
    .C1(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__a221o_1 _6338_ (.A1(\gpio_configure[28][12] ),
    .A2(_2850_),
    .B1(_2851_),
    .B2(\gpio_configure[20][12] ),
    .C1(_3138_),
    .X(_3141_));
 sky130_fd_sc_hd__a22o_1 _6339_ (.A1(\gpio_configure[33][12] ),
    .A2(_2832_),
    .B1(_2845_),
    .B2(\gpio_configure[22][12] ),
    .X(_3142_));
 sky130_fd_sc_hd__a221o_1 _6340_ (.A1(\gpio_configure[18][12] ),
    .A2(_2802_),
    .B1(_2833_),
    .B2(\gpio_configure[8][12] ),
    .C1(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__a22o_1 _6341_ (.A1(\gpio_configure[27][12] ),
    .A2(_2824_),
    .B1(_2827_),
    .B2(\gpio_configure[14][12] ),
    .X(_3144_));
 sky130_fd_sc_hd__a221o_2 _6342_ (.A1(\gpio_configure[16][12] ),
    .A2(_2843_),
    .B1(_2849_),
    .B2(\gpio_configure[17][12] ),
    .C1(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__or4_1 _6343_ (.A(_3140_),
    .B(_3141_),
    .C(_3143_),
    .D(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__a22o_1 _6344_ (.A1(\gpio_configure[32][12] ),
    .A2(_2808_),
    .B1(_2817_),
    .B2(\gpio_configure[37][12] ),
    .X(_3147_));
 sky130_fd_sc_hd__a221o_2 _6345_ (.A1(\gpio_configure[4][12] ),
    .A2(_2807_),
    .B1(_2834_),
    .B2(\gpio_configure[36][12] ),
    .C1(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__a221o_2 _6346_ (.A1(\gpio_configure[34][12] ),
    .A2(_2814_),
    .B1(_2848_),
    .B2(\gpio_configure[19][12] ),
    .C1(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__a22o_1 _6347_ (.A1(\gpio_configure[12][12] ),
    .A2(_2821_),
    .B1(_2822_),
    .B2(\gpio_configure[9][12] ),
    .X(_3150_));
 sky130_fd_sc_hd__a221o_1 _6348_ (.A1(\gpio_configure[6][12] ),
    .A2(_2809_),
    .B1(_2812_),
    .B2(\gpio_configure[10][12] ),
    .C1(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__a22o_1 _6349_ (.A1(\gpio_configure[13][12] ),
    .A2(_2831_),
    .B1(_2847_),
    .B2(\gpio_configure[25][12] ),
    .X(_3152_));
 sky130_fd_sc_hd__a221o_1 _6350_ (.A1(\gpio_configure[2][12] ),
    .A2(_2819_),
    .B1(_2820_),
    .B2(\gpio_configure[5][12] ),
    .C1(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__a22o_1 _6351_ (.A1(\gpio_configure[31][12] ),
    .A2(_2485_),
    .B1(_2830_),
    .B2(\gpio_configure[11][12] ),
    .X(_3154_));
 sky130_fd_sc_hd__a221o_1 _6352_ (.A1(\gpio_configure[1][12] ),
    .A2(_2829_),
    .B1(_2844_),
    .B2(\gpio_configure[24][12] ),
    .C1(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__a22o_1 _6353_ (.A1(\gpio_configure[26][12] ),
    .A2(_2811_),
    .B1(_2823_),
    .B2(\gpio_configure[7][12] ),
    .X(_3156_));
 sky130_fd_sc_hd__a221o_1 _6354_ (.A1(\gpio_configure[15][12] ),
    .A2(_2815_),
    .B1(_2818_),
    .B2(\gpio_configure[3][12] ),
    .C1(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__or4_2 _6355_ (.A(_3151_),
    .B(_3153_),
    .C(_3155_),
    .D(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__or4_2 _6356_ (.A(net350),
    .B(_3146_),
    .C(_3149_),
    .D(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__o211a_4 _6357_ (.A1(\gpio_configure[0][12] ),
    .A2(_2842_),
    .B1(_3159_),
    .C1(net405),
    .X(_3160_));
 sky130_fd_sc_hd__a21o_1 _6358_ (.A1(net408),
    .A2(\serial_data_staging_2[11] ),
    .B1(net353),
    .X(_3161_));
 sky130_fd_sc_hd__o22a_1 _6359_ (.A1(\serial_data_staging_2[12] ),
    .A2(net352),
    .B1(_3160_),
    .B2(_3161_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(_0816_),
    .B(\wbbd_state[6] ),
    .Y(_3162_));
 sky130_fd_sc_hd__a32o_1 _6361_ (.A1(net317),
    .A2(_1441_),
    .A3(_3162_),
    .B1(_1453_),
    .B2(\wbbd_state[1] ),
    .X(_0790_));
 sky130_fd_sc_hd__and2_4 _6362_ (.A(\wbbd_state[1] ),
    .B(net457),
    .X(_3163_));
 sky130_fd_sc_hd__mux2_1 _6363_ (.A0(net334),
    .A1(_1373_),
    .S(_3163_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _6364_ (.A0(net335),
    .A1(_1308_),
    .S(_3163_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _6365_ (.A0(net336),
    .A1(_1247_),
    .S(_3163_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _6366_ (.A0(net337),
    .A1(_1189_),
    .S(_3163_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _6367_ (.A0(net338),
    .A1(clknet_1_1__leaf__1132_),
    .S(_3163_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _6368_ (.A0(net339),
    .A1(_1037_),
    .S(_3163_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _6369_ (.A0(net341),
    .A1(_1002_),
    .S(_3163_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _6370_ (.A0(net342),
    .A1(_0968_),
    .S(_3163_),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _6371_ (.A(net170),
    .B(net166),
    .Y(_3164_));
 sky130_fd_sc_hd__nand2_1 _6372_ (.A(net170),
    .B(net167),
    .Y(_3165_));
 sky130_fd_sc_hd__a22o_1 _6373_ (.A1(\wbbd_state[8] ),
    .A2(_3164_),
    .B1(_3165_),
    .B2(\wbbd_state[7] ),
    .X(_3166_));
 sky130_fd_sc_hd__a21bo_1 _6374_ (.A1(net170),
    .A2(net165),
    .B1_N(\wbbd_state[5] ),
    .X(_3167_));
 sky130_fd_sc_hd__a21boi_1 _6375_ (.A1(net168),
    .A2(net170),
    .B1_N(\wbbd_state[9] ),
    .Y(_3168_));
 sky130_fd_sc_hd__or4b_4 _6376_ (.A(_1534_),
    .B(_3168_),
    .C(_3166_),
    .D_N(_3167_),
    .X(_3169_));
 sky130_fd_sc_hd__a22o_1 _6377_ (.A1(\wbbd_state[7] ),
    .A2(net139),
    .B1(net162),
    .B2(\wbbd_state[8] ),
    .X(_3170_));
 sky130_fd_sc_hd__a221o_1 _6378_ (.A1(\wbbd_state[9] ),
    .A2(net148),
    .B1(net132),
    .B2(_1532_),
    .C1(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__mux2_1 _6379_ (.A0(_3171_),
    .A1(\wbbd_data[0] ),
    .S(_3169_),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _6380_ (.A1(\wbbd_state[9] ),
    .A2(net149),
    .B1(net163),
    .B2(\wbbd_state[8] ),
    .X(_3172_));
 sky130_fd_sc_hd__a221o_1 _6381_ (.A1(\wbbd_state[7] ),
    .A2(net140),
    .B1(net143),
    .B2(_1532_),
    .C1(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__mux2_1 _6382_ (.A0(_3173_),
    .A1(\wbbd_data[1] ),
    .S(_3169_),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _6383_ (.A1(\wbbd_state[7] ),
    .A2(net141),
    .B1(net154),
    .B2(_1532_),
    .X(_3174_));
 sky130_fd_sc_hd__a221o_1 _6384_ (.A1(\wbbd_state[9] ),
    .A2(net150),
    .B1(net133),
    .B2(\wbbd_state[8] ),
    .C1(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(_3175_),
    .A1(\wbbd_data[2] ),
    .S(_3169_),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_1 _6386_ (.A1(\wbbd_state[9] ),
    .A2(net151),
    .B1(net134),
    .B2(\wbbd_state[8] ),
    .X(_3176_));
 sky130_fd_sc_hd__a221o_1 _6387_ (.A1(\wbbd_state[7] ),
    .A2(net142),
    .B1(net157),
    .B2(_1532_),
    .C1(_3176_),
    .X(_3177_));
 sky130_fd_sc_hd__mux2_1 _6388_ (.A0(_3177_),
    .A1(\wbbd_data[3] ),
    .S(_3169_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _6389_ (.A1(\wbbd_state[7] ),
    .A2(net144),
    .B1(net158),
    .B2(_1532_),
    .X(_3178_));
 sky130_fd_sc_hd__a221o_1 _6390_ (.A1(\wbbd_state[9] ),
    .A2(net152),
    .B1(net135),
    .B2(\wbbd_state[8] ),
    .C1(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__mux2_1 _6391_ (.A0(_3179_),
    .A1(\wbbd_data[4] ),
    .S(_3169_),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(\wbbd_state[7] ),
    .A2(net145),
    .B1(net136),
    .B2(\wbbd_state[8] ),
    .X(_3180_));
 sky130_fd_sc_hd__a221o_1 _6393_ (.A1(\wbbd_state[9] ),
    .A2(net153),
    .B1(net159),
    .B2(_1532_),
    .C1(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(_3181_),
    .A1(\wbbd_data[5] ),
    .S(_3169_),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _6395_ (.A1(\wbbd_state[7] ),
    .A2(net146),
    .B1(net137),
    .B2(\wbbd_state[8] ),
    .X(_3182_));
 sky130_fd_sc_hd__a221o_1 _6396_ (.A1(\wbbd_state[9] ),
    .A2(net155),
    .B1(net160),
    .B2(_1532_),
    .C1(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__mux2_1 _6397_ (.A0(_3183_),
    .A1(\wbbd_data[6] ),
    .S(_3169_),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _6398_ (.A1(\wbbd_state[9] ),
    .A2(net156),
    .B1(net138),
    .B2(\wbbd_state[8] ),
    .X(_3184_));
 sky130_fd_sc_hd__a221o_1 _6399_ (.A1(\wbbd_state[7] ),
    .A2(net147),
    .B1(net161),
    .B2(_1532_),
    .C1(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__mux2_1 _6400_ (.A0(_3185_),
    .A1(\wbbd_data[7] ),
    .S(_3169_),
    .X(_0806_));
 sky130_fd_sc_hd__o211a_2 _6401_ (.A1(clknet_1_1__leaf_wbbd_sck),
    .A2(_1533_),
    .B1(_1534_),
    .C1(_0817_),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _6402_ (.A1(\wbbd_state[9] ),
    .A2(net168),
    .B1(net167),
    .B2(\wbbd_state[7] ),
    .X(_3186_));
 sky130_fd_sc_hd__a21o_1 _6403_ (.A1(\wbbd_state[8] ),
    .A2(net166),
    .B1(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__a32o_4 _6404_ (.A1(_0817_),
    .A2(_1532_),
    .A3(_3167_),
    .B1(_3187_),
    .B2(net170),
    .X(_3188_));
 sky130_fd_sc_hd__o31a_1 _6405_ (.A1(wbbd_write),
    .A2(\wbbd_state[6] ),
    .A3(_1535_),
    .B1(_3188_),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_4 _6406_ (.A(_1081_),
    .B(net362),
    .Y(_3189_));
 sky130_fd_sc_hd__mux2_1 _6407_ (.A0(net400),
    .A1(net1620),
    .S(_3189_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _6408_ (.A0(net395),
    .A1(net979),
    .S(_3189_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _6409_ (.A0(net388),
    .A1(net1457),
    .S(_3189_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(net383),
    .A1(net1439),
    .S(_3189_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _6411_ (.A0(net379),
    .A1(net1212),
    .S(_3189_),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(net416),
    .B(net411),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _6413_ (.A(net415),
    .B(net410),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _6414_ (.A(net415),
    .B(net410),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _6415_ (.A(net441),
    .B(net413),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _6416_ (.A(net441),
    .B(net413),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _6417_ (.A(net441),
    .B(net413),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _6418_ (.A(net441),
    .B(net413),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _6419_ (.A(net441),
    .B(net413),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(net441),
    .B(net413),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _6421_ (.A(net441),
    .B(net413),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _6422_ (.A(net416),
    .B(net411),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _6423_ (.A(net416),
    .B(net411),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _6424_ (.A(net416),
    .B(net411),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net416),
    .B(net410),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(net416),
    .B(net411),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _6427_ (.A(net416),
    .B(net411),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(net416),
    .B(net410),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _6429_ (.A(net415),
    .B(net410),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(net416),
    .B(net411),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net415),
    .B(net410),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net415),
    .B(net410),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net415),
    .B(net410),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(net415),
    .B(net410),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(net414),
    .B(net410),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(net414),
    .B(net410),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(net415),
    .B(net410),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _6438_ (.A(net414),
    .B(net410),
    .X(_0047_));
 sky130_fd_sc_hd__and2_1 _6439_ (.A(net414),
    .B(net410),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(net415),
    .B(net410),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(net415),
    .B(net410),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _6442_ (.A(net415),
    .B(net410),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(net416),
    .B(net410),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _6444_ (.A(net415),
    .B(net410),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _6445_ (.A(net416),
    .B(net411),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _6446_ (.A(net415),
    .B(net410),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _6447_ (.A(net416),
    .B(net411),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _6448_ (.A(net416),
    .B(net411),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(net416),
    .B(net411),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _6450_ (.A(net425),
    .B(net411),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _6451_ (.A(net425),
    .B(net412),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _6452_ (.A(net425),
    .B(net412),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _6453_ (.A(net425),
    .B(net412),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _6454_ (.A(net425),
    .B(net412),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(net416),
    .B(net411),
    .X(_0064_));
 sky130_fd_sc_hd__dfrtn_1 _6456_ (.CLK_N(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0065_),
    .RESET_B(_0019_),
    .Q(\hkspi.wrstb ));
 sky130_fd_sc_hd__dfrtp_2 _6457_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0066_),
    .RESET_B(_0020_),
    .Q(\hkspi.pre_pass_thru_user ));
 sky130_fd_sc_hd__dfstp_4 _6458_ (.CLK(net461),
    .D(_0018_),
    .SET_B(_0021_),
    .Q(\hkspi.sdoenb ));
 sky130_fd_sc_hd__dfrtp_2 _6459_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0067_),
    .RESET_B(_0023_),
    .Q(\hkspi.pre_pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_2 _6460_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0068_),
    .RESET_B(_0024_),
    .Q(\hkspi.odata[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6461_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0069_),
    .RESET_B(_0025_),
    .Q(\hkspi.odata[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6462_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0070_),
    .RESET_B(_0026_),
    .Q(\hkspi.odata[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6463_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0071_),
    .RESET_B(_0027_),
    .Q(\hkspi.odata[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6464_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0072_),
    .RESET_B(_0028_),
    .Q(\hkspi.odata[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6465_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0073_),
    .RESET_B(_0029_),
    .Q(\hkspi.odata[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6466_ (.CLK(clknet_2_3_0_mgmt_gpio_in[4]),
    .D(_0074_),
    .RESET_B(_0030_),
    .Q(\hkspi.odata[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6467_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0075_),
    .RESET_B(_0031_),
    .Q(\hkspi.fixed[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6468_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0076_),
    .RESET_B(_0032_),
    .Q(\hkspi.fixed[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6469_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0077_),
    .RESET_B(_0033_),
    .Q(\hkspi.fixed[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6470_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0078_),
    .RESET_B(_0034_),
    .Q(\hkspi.readmode ));
 sky130_fd_sc_hd__dfrtp_4 _6471_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0079_),
    .RESET_B(_0035_),
    .Q(\hkspi.writemode ));
 sky130_fd_sc_hd__dfrtp_2 _6472_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0080_),
    .RESET_B(_0036_),
    .Q(\hkspi.rdstb ));
 sky130_fd_sc_hd__dfrtp_2 _6473_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0081_),
    .RESET_B(_0037_),
    .Q(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_2 _6474_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0082_),
    .RESET_B(_0038_),
    .Q(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__dfrtp_2 _6475_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0083_),
    .RESET_B(_0039_),
    .Q(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__dfrtp_2 _6476_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0084_),
    .RESET_B(_0040_),
    .Q(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__dfrtp_2 _6477_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0085_),
    .RESET_B(_0041_),
    .Q(\hkspi.addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6478_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0086_),
    .RESET_B(_0042_),
    .Q(\hkspi.addr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6479_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0087_),
    .RESET_B(_0043_),
    .Q(\hkspi.addr[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6480_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0088_),
    .RESET_B(_0044_),
    .Q(\hkspi.addr[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6481_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0089_),
    .RESET_B(_0045_),
    .Q(\hkspi.addr[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6482_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0090_),
    .RESET_B(_0046_),
    .Q(\hkspi.addr[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6483_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0091_),
    .RESET_B(_0047_),
    .Q(\hkspi.addr[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6484_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0092_),
    .RESET_B(_0048_),
    .Q(\hkspi.addr[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6485_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0093_),
    .RESET_B(_0049_),
    .Q(\hkspi.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6486_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0094_),
    .RESET_B(_0050_),
    .Q(\hkspi.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6487_ (.CLK(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0095_),
    .RESET_B(_0051_),
    .Q(\hkspi.count[2] ));
 sky130_fd_sc_hd__dfstp_2 _6488_ (.CLK(clknet_leaf_72_csclk),
    .D(net1666),
    .SET_B(net421),
    .Q(net299));
 sky130_fd_sc_hd__dfstp_4 _6489_ (.CLK(clknet_leaf_72_csclk),
    .D(_0097_),
    .SET_B(net421),
    .Q(net300));
 sky130_fd_sc_hd__dfstp_4 _6490_ (.CLK(clknet_leaf_72_csclk),
    .D(_0098_),
    .SET_B(net421),
    .Q(net276));
 sky130_fd_sc_hd__dfstp_2 _6491_ (.CLK(clknet_leaf_72_csclk),
    .D(_0099_),
    .SET_B(net421),
    .Q(net277));
 sky130_fd_sc_hd__dfrtp_2 _6492_ (.CLK(clknet_leaf_71_csclk),
    .D(net933),
    .RESET_B(net421),
    .Q(net278));
 sky130_fd_sc_hd__dfstp_4 _6493_ (.CLK(clknet_leaf_58_csclk),
    .D(_0101_),
    .SET_B(net428),
    .Q(net279));
 sky130_fd_sc_hd__dfstp_4 _6494_ (.CLK(clknet_leaf_58_csclk),
    .D(_0102_),
    .SET_B(net428),
    .Q(net280));
 sky130_fd_sc_hd__dfstp_4 _6495_ (.CLK(clknet_leaf_58_csclk),
    .D(_0103_),
    .SET_B(net429),
    .Q(net281));
 sky130_fd_sc_hd__dfstp_4 _6496_ (.CLK(clknet_leaf_75_csclk),
    .D(_0104_),
    .SET_B(net419),
    .Q(net275));
 sky130_fd_sc_hd__dfstp_4 _6497_ (.CLK(clknet_leaf_72_csclk),
    .D(_0105_),
    .SET_B(net419),
    .Q(net286));
 sky130_fd_sc_hd__dfstp_4 _6498_ (.CLK(clknet_leaf_75_csclk),
    .D(_0106_),
    .SET_B(net419),
    .Q(net293));
 sky130_fd_sc_hd__dfstp_4 _6499_ (.CLK(clknet_leaf_75_csclk),
    .D(_0107_),
    .SET_B(net419),
    .Q(net294));
 sky130_fd_sc_hd__dfstp_4 _6500_ (.CLK(clknet_leaf_72_csclk),
    .D(_0108_),
    .SET_B(net419),
    .Q(net295));
 sky130_fd_sc_hd__dfstp_4 _6501_ (.CLK(clknet_leaf_72_csclk),
    .D(_0109_),
    .SET_B(net419),
    .Q(net296));
 sky130_fd_sc_hd__dfstp_4 _6502_ (.CLK(clknet_leaf_72_csclk),
    .D(net689),
    .SET_B(net421),
    .Q(net297));
 sky130_fd_sc_hd__dfstp_4 _6503_ (.CLK(clknet_leaf_72_csclk),
    .D(_0111_),
    .SET_B(net421),
    .Q(net298));
 sky130_fd_sc_hd__dfstp_4 _6504_ (.CLK(clknet_leaf_71_csclk),
    .D(_0112_),
    .SET_B(net429),
    .Q(net291));
 sky130_fd_sc_hd__dfstp_4 _6505_ (.CLK(clknet_leaf_71_csclk),
    .D(net624),
    .SET_B(net429),
    .Q(net292));
 sky130_fd_sc_hd__dfrtp_2 _6506_ (.CLK(clknet_leaf_37_csclk),
    .D(net1411),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6507_ (.CLK(clknet_leaf_36_csclk),
    .D(net1182),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6508_ (.CLK(clknet_leaf_37_csclk),
    .D(net1339),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data[10] ));
 sky130_fd_sc_hd__dfrtp_2 _6509_ (.CLK(clknet_leaf_36_csclk),
    .D(net1406),
    .RESET_B(net453),
    .Q(net215));
 sky130_fd_sc_hd__dfrtp_2 _6510_ (.CLK(clknet_leaf_38_csclk),
    .D(net1233),
    .RESET_B(net450),
    .Q(net216));
 sky130_fd_sc_hd__dfrtp_2 _6511_ (.CLK(clknet_leaf_30_csclk),
    .D(net1265),
    .RESET_B(net447),
    .Q(\mgmt_gpio_data[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6512_ (.CLK(clknet_leaf_37_csclk),
    .D(net1352),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6513_ (.CLK(clknet_leaf_32_csclk),
    .D(net744),
    .RESET_B(net447),
    .Q(\mgmt_gpio_data[15] ));
 sky130_fd_sc_hd__dfrtp_2 _6514_ (.CLK(clknet_leaf_30_csclk),
    .D(net1445),
    .RESET_B(net447),
    .Q(net229));
 sky130_fd_sc_hd__dfrtp_2 _6515_ (.CLK(clknet_leaf_30_csclk),
    .D(net772),
    .RESET_B(net447),
    .Q(net230));
 sky130_fd_sc_hd__dfrtp_2 _6516_ (.CLK(clknet_leaf_31_csclk),
    .D(net972),
    .RESET_B(net447),
    .Q(net231));
 sky130_fd_sc_hd__dfrtp_2 _6517_ (.CLK(clknet_leaf_31_csclk),
    .D(net628),
    .RESET_B(net452),
    .Q(net232));
 sky130_fd_sc_hd__dfrtp_2 _6518_ (.CLK(clknet_leaf_31_csclk),
    .D(net715),
    .RESET_B(net452),
    .Q(net233));
 sky130_fd_sc_hd__dfrtp_2 _6519_ (.CLK(clknet_leaf_34_csclk),
    .D(net847),
    .RESET_B(net452),
    .Q(net234));
 sky130_fd_sc_hd__dfrtp_2 _6520_ (.CLK(clknet_leaf_34_csclk),
    .D(net1000),
    .RESET_B(net452),
    .Q(net236));
 sky130_fd_sc_hd__dfrtp_2 _6521_ (.CLK(clknet_leaf_34_csclk),
    .D(net782),
    .RESET_B(net452),
    .Q(net237));
 sky130_fd_sc_hd__dfrtp_1 _6522_ (.CLK(clknet_leaf_37_csclk),
    .D(net1222),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data_buf[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6523_ (.CLK(clknet_leaf_36_csclk),
    .D(net784),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6524_ (.CLK(clknet_leaf_37_csclk),
    .D(net988),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data_buf[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6525_ (.CLK(clknet_leaf_36_csclk),
    .D(net1178),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6526_ (.CLK(clknet_leaf_37_csclk),
    .D(net730),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data_buf[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6527_ (.CLK(clknet_leaf_30_csclk),
    .D(net874),
    .RESET_B(net447),
    .Q(\mgmt_gpio_data_buf[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6528_ (.CLK(clknet_leaf_37_csclk),
    .D(net593),
    .RESET_B(net450),
    .Q(\mgmt_gpio_data_buf[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6529_ (.CLK(clknet_leaf_30_csclk),
    .D(net818),
    .RESET_B(net447),
    .Q(\mgmt_gpio_data_buf[15] ));
 sky130_fd_sc_hd__dfrtp_2 _6530_ (.CLK(clknet_leaf_1_csclk),
    .D(net1693),
    .RESET_B(net417),
    .Q(\gpio_configure[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6531_ (.CLK(clknet_leaf_1_csclk),
    .D(net1362),
    .RESET_B(net417),
    .Q(\gpio_configure[0][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6532_ (.CLK(clknet_leaf_1_csclk),
    .D(net1461),
    .RESET_B(net422),
    .Q(\gpio_configure[0][10] ));
 sky130_fd_sc_hd__dfstp_4 _6533_ (.CLK(clknet_leaf_2_csclk),
    .D(_0141_),
    .SET_B(net424),
    .Q(\gpio_configure[0][11] ));
 sky130_fd_sc_hd__dfstp_4 _6534_ (.CLK(clknet_leaf_2_csclk),
    .D(_0142_),
    .SET_B(net424),
    .Q(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6535_ (.CLK(clknet_leaf_2_csclk),
    .D(net1676),
    .RESET_B(net424),
    .Q(\gpio_configure[1][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6536_ (.CLK(clknet_leaf_1_csclk),
    .D(net1354),
    .RESET_B(net417),
    .Q(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6537_ (.CLK(clknet_leaf_3_csclk),
    .D(net1137),
    .RESET_B(net424),
    .Q(\gpio_configure[1][10] ));
 sky130_fd_sc_hd__dfstp_4 _6538_ (.CLK(clknet_leaf_1_csclk),
    .D(_0146_),
    .SET_B(net417),
    .Q(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__dfstp_4 _6539_ (.CLK(clknet_leaf_2_csclk),
    .D(_0147_),
    .SET_B(net424),
    .Q(\gpio_configure[1][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6540_ (.CLK(clknet_leaf_15_csclk),
    .D(net1562),
    .RESET_B(net440),
    .Q(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6541_ (.CLK(clknet_leaf_1_csclk),
    .D(net1356),
    .RESET_B(net417),
    .Q(\gpio_configure[2][9] ));
 sky130_fd_sc_hd__dfstp_4 _6542_ (.CLK(clknet_leaf_13_csclk),
    .D(_0150_),
    .SET_B(net440),
    .Q(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6543_ (.CLK(clknet_leaf_2_csclk),
    .D(net1469),
    .RESET_B(net418),
    .Q(\gpio_configure[2][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6544_ (.CLK(clknet_leaf_2_csclk),
    .D(net1511),
    .RESET_B(net424),
    .Q(\gpio_configure[2][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6545_ (.CLK(clknet_leaf_11_csclk),
    .D(net1590),
    .RESET_B(net439),
    .Q(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6546_ (.CLK(clknet_leaf_12_csclk),
    .D(net786),
    .RESET_B(net439),
    .Q(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6547_ (.CLK(clknet_leaf_11_csclk),
    .D(net1421),
    .RESET_B(net439),
    .Q(\gpio_configure[3][10] ));
 sky130_fd_sc_hd__dfstp_4 _6548_ (.CLK(clknet_leaf_3_csclk),
    .D(_0156_),
    .SET_B(net424),
    .Q(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6549_ (.CLK(clknet_leaf_3_csclk),
    .D(net1506),
    .RESET_B(net424),
    .Q(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6550_ (.CLK(clknet_leaf_16_csclk),
    .D(net1584),
    .RESET_B(net441),
    .Q(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6551_ (.CLK(clknet_leaf_14_csclk),
    .D(net1120),
    .RESET_B(net441),
    .Q(\gpio_configure[4][9] ));
 sky130_fd_sc_hd__dfstp_4 _6552_ (.CLK(clknet_leaf_15_csclk),
    .D(_0160_),
    .SET_B(net440),
    .Q(\gpio_configure[4][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6553_ (.CLK(clknet_leaf_16_csclk),
    .D(net768),
    .RESET_B(net440),
    .Q(\gpio_configure[4][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6554_ (.CLK(clknet_leaf_16_csclk),
    .D(net1341),
    .RESET_B(net441),
    .Q(\gpio_configure[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _6555_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0163_),
    .Q(net325));
 sky130_fd_sc_hd__dfxtp_4 _6556_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0164_),
    .Q(net326));
 sky130_fd_sc_hd__dfxtp_2 _6557_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0165_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_2 _6558_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0166_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_4 _6559_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0167_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_4 _6560_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0168_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_4 _6561_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0169_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_4 _6562_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0170_),
    .Q(net333));
 sky130_fd_sc_hd__dfrtp_2 _6563_ (.CLK(clknet_leaf_10_csclk),
    .D(net1642),
    .RESET_B(net439),
    .Q(\gpio_configure[5][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6564_ (.CLK(clknet_leaf_12_csclk),
    .D(net807),
    .RESET_B(net439),
    .Q(\gpio_configure[5][9] ));
 sky130_fd_sc_hd__dfstp_2 _6565_ (.CLK(clknet_leaf_13_csclk),
    .D(net1449),
    .SET_B(net439),
    .Q(\gpio_configure[5][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6566_ (.CLK(clknet_leaf_12_csclk),
    .D(net534),
    .RESET_B(net439),
    .Q(\gpio_configure[5][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6567_ (.CLK(clknet_leaf_12_csclk),
    .D(net674),
    .RESET_B(net439),
    .Q(\gpio_configure[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6568_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0176_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_2 _6569_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0177_),
    .Q(net349));
 sky130_fd_sc_hd__dfxtp_2 _6570_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0178_),
    .Q(net319));
 sky130_fd_sc_hd__dfxtp_2 _6571_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0179_),
    .Q(net320));
 sky130_fd_sc_hd__dfxtp_2 _6572_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0180_),
    .Q(net321));
 sky130_fd_sc_hd__dfxtp_2 _6573_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0181_),
    .Q(net322));
 sky130_fd_sc_hd__dfxtp_2 _6574_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0182_),
    .Q(net323));
 sky130_fd_sc_hd__dfxtp_4 _6575_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0183_),
    .Q(net324));
 sky130_fd_sc_hd__dfrtp_2 _6576_ (.CLK(clknet_leaf_4_csclk),
    .D(net1588),
    .RESET_B(net426),
    .Q(\gpio_configure[6][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6577_ (.CLK(clknet_leaf_3_csclk),
    .D(net958),
    .RESET_B(net424),
    .Q(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__dfstp_4 _6578_ (.CLK(clknet_leaf_4_csclk),
    .D(_0186_),
    .SET_B(net426),
    .Q(\gpio_configure[6][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6579_ (.CLK(clknet_leaf_4_csclk),
    .D(net1243),
    .RESET_B(net426),
    .Q(\gpio_configure[6][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6580_ (.CLK(clknet_leaf_4_csclk),
    .D(net1502),
    .RESET_B(net426),
    .Q(\gpio_configure[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6581_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0189_),
    .Q(net318));
 sky130_fd_sc_hd__dfxtp_2 _6582_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0190_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_1 _6583_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0191_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_2 _6584_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0192_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_2 _6585_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0193_),
    .Q(net344));
 sky130_fd_sc_hd__dfxtp_2 _6586_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0194_),
    .Q(net345));
 sky130_fd_sc_hd__dfxtp_2 _6587_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0195_),
    .Q(net346));
 sky130_fd_sc_hd__dfxtp_2 _6588_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0196_),
    .Q(net347));
 sky130_fd_sc_hd__dfrtp_2 _6589_ (.CLK(clknet_leaf_11_csclk),
    .D(net1601),
    .RESET_B(net439),
    .Q(\gpio_configure[7][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6590_ (.CLK(clknet_leaf_5_csclk),
    .D(net1020),
    .RESET_B(net426),
    .Q(\gpio_configure[7][9] ));
 sky130_fd_sc_hd__dfstp_2 _6591_ (.CLK(clknet_leaf_11_csclk),
    .D(_0199_),
    .SET_B(net439),
    .Q(\gpio_configure[7][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6592_ (.CLK(clknet_leaf_5_csclk),
    .D(net1292),
    .RESET_B(net426),
    .Q(\gpio_configure[7][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6593_ (.CLK(clknet_leaf_5_csclk),
    .D(net1528),
    .RESET_B(net426),
    .Q(\gpio_configure[7][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6594_ (.CLK(clknet_leaf_3_csclk),
    .D(net1668),
    .RESET_B(net424),
    .Q(\gpio_configure[8][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6595_ (.CLK(clknet_leaf_3_csclk),
    .D(net976),
    .RESET_B(net424),
    .Q(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__dfstp_4 _6596_ (.CLK(clknet_leaf_3_csclk),
    .D(_0204_),
    .SET_B(net424),
    .Q(\gpio_configure[8][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6597_ (.CLK(clknet_leaf_3_csclk),
    .D(net1224),
    .RESET_B(net424),
    .Q(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6598_ (.CLK(clknet_leaf_3_csclk),
    .D(net1493),
    .RESET_B(net424),
    .Q(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6599_ (.CLK(clknet_leaf_21_csclk),
    .D(net1592),
    .RESET_B(net440),
    .Q(\gpio_configure[9][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6600_ (.CLK(clknet_leaf_15_csclk),
    .D(net994),
    .RESET_B(net440),
    .Q(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__dfstp_4 _6601_ (.CLK(clknet_leaf_15_csclk),
    .D(_0209_),
    .SET_B(net440),
    .Q(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6602_ (.CLK(clknet_leaf_15_csclk),
    .D(net695),
    .RESET_B(net440),
    .Q(\gpio_configure[9][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6603_ (.CLK(clknet_leaf_15_csclk),
    .D(net1269),
    .RESET_B(net440),
    .Q(\gpio_configure[9][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6604_ (.CLK(clknet_leaf_11_csclk),
    .D(net1603),
    .RESET_B(net439),
    .Q(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6605_ (.CLK(clknet_leaf_2_csclk),
    .D(net966),
    .RESET_B(net425),
    .Q(\gpio_configure[10][9] ));
 sky130_fd_sc_hd__dfstp_2 _6606_ (.CLK(clknet_leaf_11_csclk),
    .D(_0214_),
    .SET_B(net439),
    .Q(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6607_ (.CLK(clknet_3_1_0_csclk),
    .D(net1513),
    .RESET_B(net425),
    .Q(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6608_ (.CLK(clknet_leaf_2_csclk),
    .D(net1515),
    .RESET_B(net425),
    .Q(\gpio_configure[10][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6609_ (.CLK(clknet_leaf_15_csclk),
    .D(net1572),
    .RESET_B(net440),
    .Q(\gpio_configure[11][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6610_ (.CLK(clknet_leaf_14_csclk),
    .D(net1144),
    .RESET_B(net440),
    .Q(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__dfstp_4 _6611_ (.CLK(clknet_leaf_15_csclk),
    .D(_0219_),
    .SET_B(net440),
    .Q(\gpio_configure[11][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6612_ (.CLK(clknet_leaf_15_csclk),
    .D(net705),
    .RESET_B(net440),
    .Q(\gpio_configure[11][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6613_ (.CLK(clknet_leaf_15_csclk),
    .D(net1257),
    .RESET_B(net440),
    .Q(\gpio_configure[11][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6614_ (.CLK(clknet_leaf_13_csclk),
    .D(net1630),
    .RESET_B(net439),
    .Q(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6615_ (.CLK(clknet_leaf_12_csclk),
    .D(net793),
    .RESET_B(net439),
    .Q(\gpio_configure[12][9] ));
 sky130_fd_sc_hd__dfstp_2 _6616_ (.CLK(clknet_leaf_13_csclk),
    .D(_0224_),
    .SET_B(net439),
    .Q(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6617_ (.CLK(clknet_leaf_5_csclk),
    .D(net1271),
    .RESET_B(net427),
    .Q(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6618_ (.CLK(clknet_leaf_5_csclk),
    .D(net1526),
    .RESET_B(net427),
    .Q(\gpio_configure[12][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6619_ (.CLK(clknet_leaf_11_csclk),
    .D(net1607),
    .RESET_B(net439),
    .Q(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6620_ (.CLK(clknet_leaf_11_csclk),
    .D(net1100),
    .RESET_B(net439),
    .Q(\gpio_configure[13][9] ));
 sky130_fd_sc_hd__dfstp_2 _6621_ (.CLK(clknet_leaf_11_csclk),
    .D(net1413),
    .SET_B(net456),
    .Q(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6622_ (.CLK(clknet_leaf_5_csclk),
    .D(net1280),
    .RESET_B(net426),
    .Q(\gpio_configure[13][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6623_ (.CLK(clknet_leaf_12_csclk),
    .D(net665),
    .RESET_B(net439),
    .Q(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6624_ (.CLK(clknet_leaf_15_csclk),
    .D(net1556),
    .RESET_B(net440),
    .Q(\gpio_configure[16][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6625_ (.CLK(clknet_leaf_15_csclk),
    .D(net998),
    .RESET_B(net440),
    .Q(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__dfstp_2 _6626_ (.CLK(clknet_leaf_15_csclk),
    .D(_0234_),
    .SET_B(net440),
    .Q(\gpio_configure[16][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6627_ (.CLK(clknet_leaf_21_csclk),
    .D(net775),
    .RESET_B(net440),
    .Q(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6628_ (.CLK(clknet_leaf_15_csclk),
    .D(net1278),
    .RESET_B(net440),
    .Q(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6629_ (.CLK(clknet_leaf_10_csclk),
    .D(net1636),
    .RESET_B(net456),
    .Q(\gpio_configure[36][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6630_ (.CLK(clknet_leaf_8_csclk),
    .D(net1058),
    .RESET_B(net427),
    .Q(\gpio_configure[36][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6631_ (.CLK(clknet_leaf_22_csclk),
    .D(net1431),
    .RESET_B(net456),
    .Q(\gpio_configure[36][10] ));
 sky130_fd_sc_hd__dfstp_4 _6632_ (.CLK(clknet_leaf_22_csclk),
    .D(_0240_),
    .SET_B(net456),
    .Q(\gpio_configure[36][11] ));
 sky130_fd_sc_hd__dfstp_1 _6633_ (.CLK(clknet_leaf_8_csclk),
    .D(_0241_),
    .SET_B(net427),
    .Q(\gpio_configure[36][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6634_ (.CLK(clknet_leaf_1_csclk),
    .D(net1617),
    .RESET_B(net417),
    .Q(\gpio_configure[31][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6635_ (.CLK(clknet_leaf_1_csclk),
    .D(net1358),
    .RESET_B(net418),
    .Q(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__dfstp_4 _6636_ (.CLK(clknet_leaf_1_csclk),
    .D(_0244_),
    .SET_B(net418),
    .Q(\gpio_configure[31][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6637_ (.CLK(clknet_leaf_1_csclk),
    .D(net1429),
    .RESET_B(net418),
    .Q(\gpio_configure[31][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6638_ (.CLK(clknet_leaf_1_csclk),
    .D(net1217),
    .RESET_B(net417),
    .Q(\gpio_configure[31][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6639_ (.CLK(clknet_leaf_1_csclk),
    .D(net1691),
    .RESET_B(net417),
    .Q(\gpio_configure[24][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6640_ (.CLK(clknet_leaf_1_csclk),
    .D(net1373),
    .RESET_B(net417),
    .Q(\gpio_configure[24][9] ));
 sky130_fd_sc_hd__dfstp_4 _6641_ (.CLK(clknet_leaf_74_csclk),
    .D(_0249_),
    .SET_B(net417),
    .Q(\gpio_configure[24][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6642_ (.CLK(clknet_leaf_78_csclk),
    .D(net1482),
    .RESET_B(net417),
    .Q(\gpio_configure[24][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6643_ (.CLK(clknet_leaf_1_csclk),
    .D(net1207),
    .RESET_B(net417),
    .Q(\gpio_configure[24][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6644_ (.CLK(clknet_leaf_67_csclk),
    .D(net1685),
    .RESET_B(net427),
    .Q(\gpio_configure[29][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6645_ (.CLK(clknet_leaf_68_csclk),
    .D(net1070),
    .RESET_B(net427),
    .Q(\gpio_configure[29][9] ));
 sky130_fd_sc_hd__dfstp_4 _6646_ (.CLK(clknet_leaf_67_csclk),
    .D(_0254_),
    .SET_B(net436),
    .Q(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6647_ (.CLK(clknet_leaf_69_csclk),
    .D(net1324),
    .RESET_B(net427),
    .Q(\gpio_configure[29][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6648_ (.CLK(clknet_leaf_68_csclk),
    .D(net1564),
    .RESET_B(net427),
    .Q(\gpio_configure[29][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6649_ (.CLK(clknet_leaf_11_csclk),
    .D(net1605),
    .RESET_B(net456),
    .Q(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6650_ (.CLK(clknet_leaf_12_csclk),
    .D(net805),
    .RESET_B(net439),
    .Q(\gpio_configure[25][9] ));
 sky130_fd_sc_hd__dfstp_4 _6651_ (.CLK(clknet_leaf_2_csclk),
    .D(_0259_),
    .SET_B(net424),
    .Q(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6652_ (.CLK(clknet_leaf_2_csclk),
    .D(net1267),
    .RESET_B(net424),
    .Q(\gpio_configure[25][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6653_ (.CLK(clknet_leaf_2_csclk),
    .D(net1521),
    .RESET_B(net424),
    .Q(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6654_ (.CLK(clknet_leaf_74_csclk),
    .D(net1628),
    .RESET_B(net422),
    .Q(\gpio_configure[28][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6655_ (.CLK(clknet_leaf_74_csclk),
    .D(net1360),
    .RESET_B(net422),
    .Q(\gpio_configure[28][9] ));
 sky130_fd_sc_hd__dfstp_4 _6656_ (.CLK(clknet_leaf_74_csclk),
    .D(_0264_),
    .SET_B(net422),
    .Q(\gpio_configure[28][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6657_ (.CLK(clknet_leaf_74_csclk),
    .D(net1435),
    .RESET_B(net422),
    .Q(\gpio_configure[28][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6658_ (.CLK(clknet_leaf_74_csclk),
    .D(net1194),
    .RESET_B(net422),
    .Q(\gpio_configure[28][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6659_ (.CLK(clknet_leaf_78_csclk),
    .D(net1640),
    .RESET_B(net417),
    .Q(\gpio_configure[26][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6660_ (.CLK(clknet_leaf_78_csclk),
    .D(net1403),
    .RESET_B(net417),
    .Q(\gpio_configure[26][9] ));
 sky130_fd_sc_hd__dfstp_4 _6661_ (.CLK(clknet_leaf_78_csclk),
    .D(_0269_),
    .SET_B(net417),
    .Q(\gpio_configure[26][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6662_ (.CLK(clknet_leaf_78_csclk),
    .D(net1496),
    .RESET_B(net417),
    .Q(\gpio_configure[26][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6663_ (.CLK(clknet_leaf_78_csclk),
    .D(net1284),
    .RESET_B(net414),
    .Q(\gpio_configure[26][12] ));
 sky130_fd_sc_hd__dfstp_4 _6664_ (.CLK(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0004_),
    .SET_B(_0052_),
    .Q(\hkspi.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6665_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0005_),
    .RESET_B(_0053_),
    .Q(\hkspi.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6666_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0006_),
    .RESET_B(_0054_),
    .Q(\hkspi.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6667_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0007_),
    .RESET_B(_0055_),
    .Q(\hkspi.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6668_ (.CLK(clknet_2_1_0_mgmt_gpio_in[4]),
    .D(_0008_),
    .RESET_B(_0056_),
    .Q(\hkspi.state[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6669_ (.CLK(clknet_leaf_36_csclk),
    .D(net1416),
    .RESET_B(net453),
    .Q(net220));
 sky130_fd_sc_hd__dfrtp_2 _6670_ (.CLK(clknet_leaf_36_csclk),
    .D(net1190),
    .RESET_B(net453),
    .Q(net221));
 sky130_fd_sc_hd__dfrtp_2 _6671_ (.CLK(clknet_leaf_36_csclk),
    .D(net1350),
    .RESET_B(net453),
    .Q(net222));
 sky130_fd_sc_hd__dfrtp_2 _6672_ (.CLK(clknet_leaf_36_csclk),
    .D(net1379),
    .RESET_B(net453),
    .Q(net223));
 sky130_fd_sc_hd__dfrtp_2 _6673_ (.CLK(clknet_leaf_29_csclk),
    .D(net922),
    .RESET_B(net446),
    .Q(net225));
 sky130_fd_sc_hd__dfrtp_2 _6674_ (.CLK(clknet_leaf_29_csclk),
    .D(net736),
    .RESET_B(net446),
    .Q(net226));
 sky130_fd_sc_hd__dfrtp_2 _6675_ (.CLK(clknet_leaf_29_csclk),
    .D(net1337),
    .RESET_B(net447),
    .Q(net227));
 sky130_fd_sc_hd__dfrtp_2 _6676_ (.CLK(clknet_leaf_29_csclk),
    .D(net717),
    .RESET_B(net448),
    .Q(net228));
 sky130_fd_sc_hd__dfstp_4 _6677_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0014_),
    .SET_B(net433),
    .Q(\xfer_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6678_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0015_),
    .RESET_B(net433),
    .Q(\xfer_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6679_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0016_),
    .RESET_B(net433),
    .Q(\xfer_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6680_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0017_),
    .RESET_B(net433),
    .Q(\xfer_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6681_ (.CLK(clknet_leaf_78_csclk),
    .D(net1689),
    .RESET_B(net416),
    .Q(\mgmt_gpio_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6682_ (.CLK(clknet_leaf_0_csclk),
    .D(net1544),
    .RESET_B(net416),
    .Q(\mgmt_gpio_data[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6683_ (.CLK(clknet_leaf_51_csclk),
    .D(net1384),
    .RESET_B(net434),
    .Q(net235));
 sky130_fd_sc_hd__dfrtp_2 _6684_ (.CLK(clknet_leaf_51_csclk),
    .D(net909),
    .RESET_B(net434),
    .Q(net244));
 sky130_fd_sc_hd__dfrtp_2 _6685_ (.CLK(clknet_leaf_47_csclk),
    .D(net1011),
    .RESET_B(net438),
    .Q(net245));
 sky130_fd_sc_hd__dfrtp_2 _6686_ (.CLK(clknet_leaf_47_csclk),
    .D(net1393),
    .RESET_B(net438),
    .Q(net246));
 sky130_fd_sc_hd__dfrtp_2 _6687_ (.CLK(clknet_leaf_0_csclk),
    .D(net986),
    .RESET_B(net416),
    .Q(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6688_ (.CLK(clknet_leaf_51_csclk),
    .D(net1310),
    .RESET_B(net434),
    .Q(net248));
 sky130_fd_sc_hd__dfrtp_2 _6689_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0288_),
    .RESET_B(net457),
    .Q(wbbd_busy));
 sky130_fd_sc_hd__dfrtp_1 _6690_ (.CLK(clknet_leaf_35_csclk),
    .D(net1419),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6691_ (.CLK(clknet_leaf_35_csclk),
    .D(net780),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6692_ (.CLK(clknet_leaf_35_csclk),
    .D(net1017),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6693_ (.CLK(clknet_leaf_35_csclk),
    .D(net1104),
    .RESET_B(net453),
    .Q(\mgmt_gpio_data_buf[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6694_ (.CLK(clknet_leaf_18_csclk),
    .D(net1276),
    .RESET_B(net446),
    .Q(\mgmt_gpio_data_buf[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6695_ (.CLK(clknet_leaf_29_csclk),
    .D(net470),
    .RESET_B(net446),
    .Q(\mgmt_gpio_data_buf[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6696_ (.CLK(clknet_leaf_29_csclk),
    .D(net984),
    .RESET_B(net448),
    .Q(\mgmt_gpio_data_buf[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6697_ (.CLK(clknet_leaf_29_csclk),
    .D(net466),
    .RESET_B(net448),
    .Q(\mgmt_gpio_data_buf[23] ));
 sky130_fd_sc_hd__dfstp_1 _6698_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0009_),
    .SET_B(net457),
    .Q(\wbbd_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6699_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0000_),
    .RESET_B(net457),
    .Q(\wbbd_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6700_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0001_),
    .RESET_B(net457),
    .Q(\wbbd_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6701_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0002_),
    .RESET_B(net457),
    .Q(\wbbd_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6702_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0003_),
    .RESET_B(net457),
    .Q(\wbbd_state[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6703_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0010_),
    .RESET_B(net457),
    .Q(\wbbd_state[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6704_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(\wbbd_state[1] ),
    .RESET_B(net457),
    .Q(\wbbd_state[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6705_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0011_),
    .RESET_B(net457),
    .Q(\wbbd_state[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6706_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0012_),
    .RESET_B(net457),
    .Q(\wbbd_state[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6707_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0013_),
    .RESET_B(net457),
    .Q(\wbbd_state[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6708_ (.CLK(clknet_leaf_4_csclk),
    .D(net1626),
    .RESET_B(net426),
    .Q(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6709_ (.CLK(clknet_leaf_4_csclk),
    .D(net952),
    .RESET_B(net426),
    .Q(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__dfstp_4 _6710_ (.CLK(clknet_leaf_4_csclk),
    .D(_0299_),
    .SET_B(net426),
    .Q(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6711_ (.CLK(clknet_leaf_4_csclk),
    .D(net1235),
    .RESET_B(net426),
    .Q(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6712_ (.CLK(clknet_leaf_4_csclk),
    .D(net1509),
    .RESET_B(net426),
    .Q(\gpio_configure[14][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6713_ (.CLK(clknet_leaf_5_csclk),
    .D(net1680),
    .RESET_B(net426),
    .Q(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6714_ (.CLK(clknet_leaf_4_csclk),
    .D(net990),
    .RESET_B(net426),
    .Q(\gpio_configure[15][9] ));
 sky130_fd_sc_hd__dfstp_4 _6715_ (.CLK(clknet_leaf_12_csclk),
    .D(_0304_),
    .SET_B(net439),
    .Q(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6716_ (.CLK(clknet_leaf_4_csclk),
    .D(net1205),
    .RESET_B(net426),
    .Q(\gpio_configure[15][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6717_ (.CLK(clknet_leaf_4_csclk),
    .D(net1499),
    .RESET_B(net426),
    .Q(\gpio_configure[15][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6718_ (.CLK(clknet_leaf_21_csclk),
    .D(net1613),
    .RESET_B(net442),
    .Q(\gpio_configure[37][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6719_ (.CLK(clknet_leaf_7_csclk),
    .D(net1074),
    .RESET_B(net427),
    .Q(\gpio_configure[37][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6720_ (.CLK(clknet_leaf_21_csclk),
    .D(net1632),
    .RESET_B(net442),
    .Q(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__dfstp_2 _6721_ (.CLK(clknet_leaf_8_csclk),
    .D(net1304),
    .SET_B(net427),
    .Q(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__dfstp_1 _6722_ (.CLK(clknet_3_1_0_csclk),
    .D(_0311_),
    .SET_B(net427),
    .Q(\gpio_configure[37][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6723_ (.CLK(clknet_leaf_15_csclk),
    .D(net1532),
    .RESET_B(net442),
    .Q(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6724_ (.CLK(clknet_leaf_7_csclk),
    .D(net1072),
    .RESET_B(net427),
    .Q(\gpio_configure[17][9] ));
 sky130_fd_sc_hd__dfstp_4 _6725_ (.CLK(clknet_leaf_15_csclk),
    .D(_0314_),
    .SET_B(net440),
    .Q(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6726_ (.CLK(clknet_leaf_7_csclk),
    .D(net1333),
    .RESET_B(net427),
    .Q(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6727_ (.CLK(clknet_leaf_8_csclk),
    .D(net1335),
    .RESET_B(net427),
    .Q(\gpio_configure[17][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6728_ (.CLK(clknet_leaf_76_csclk),
    .D(net1638),
    .RESET_B(net414),
    .Q(\gpio_configure[18][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6729_ (.CLK(clknet_leaf_76_csclk),
    .D(net1397),
    .RESET_B(net414),
    .Q(\gpio_configure[18][9] ));
 sky130_fd_sc_hd__dfstp_4 _6730_ (.CLK(clknet_leaf_76_csclk),
    .D(_0319_),
    .SET_B(net414),
    .Q(\gpio_configure[18][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6731_ (.CLK(clknet_leaf_76_csclk),
    .D(net1480),
    .RESET_B(net414),
    .Q(\gpio_configure[18][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6732_ (.CLK(clknet_leaf_76_csclk),
    .D(net1251),
    .RESET_B(net414),
    .Q(\gpio_configure[18][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6733_ (.CLK(clknet_leaf_17_csclk),
    .D(net1368),
    .RESET_B(net441),
    .Q(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6734_ (.CLK(clknet_leaf_69_csclk),
    .D(net1029),
    .RESET_B(net427),
    .Q(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__dfstp_4 _6735_ (.CLK(clknet_leaf_16_csclk),
    .D(_0324_),
    .SET_B(net441),
    .Q(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6736_ (.CLK(clknet_leaf_69_csclk),
    .D(net1328),
    .RESET_B(net427),
    .Q(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6737_ (.CLK(clknet_leaf_69_csclk),
    .D(net1388),
    .RESET_B(net427),
    .Q(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6738_ (.CLK(clknet_leaf_75_csclk),
    .D(net1657),
    .RESET_B(net419),
    .Q(\gpio_configure[19][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6739_ (.CLK(clknet_leaf_72_csclk),
    .D(net876),
    .RESET_B(net421),
    .Q(\gpio_configure[19][9] ));
 sky130_fd_sc_hd__dfstp_4 _6740_ (.CLK(clknet_leaf_72_csclk),
    .D(_0329_),
    .SET_B(net421),
    .Q(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6741_ (.CLK(clknet_leaf_72_csclk),
    .D(net1453),
    .RESET_B(net419),
    .Q(\gpio_configure[19][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6742_ (.CLK(clknet_leaf_72_csclk),
    .D(net1202),
    .RESET_B(net419),
    .Q(\gpio_configure[19][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6743_ (.CLK(clknet_leaf_16_csclk),
    .D(net1582),
    .RESET_B(net442),
    .Q(\gpio_configure[34][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6744_ (.CLK(clknet_leaf_69_csclk),
    .D(net1031),
    .RESET_B(net427),
    .Q(\gpio_configure[34][9] ));
 sky130_fd_sc_hd__dfstp_4 _6745_ (.CLK(clknet_leaf_16_csclk),
    .D(_0334_),
    .SET_B(net442),
    .Q(\gpio_configure[34][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6746_ (.CLK(clknet_leaf_8_csclk),
    .D(net1298),
    .RESET_B(net427),
    .Q(\gpio_configure[34][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6747_ (.CLK(clknet_leaf_7_csclk),
    .D(net1567),
    .RESET_B(net456),
    .Q(\gpio_configure[34][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6748_ (.CLK(clknet_leaf_75_csclk),
    .D(net1655),
    .RESET_B(net419),
    .Q(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6749_ (.CLK(clknet_leaf_75_csclk),
    .D(net1370),
    .RESET_B(net419),
    .Q(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__dfstp_4 _6750_ (.CLK(clknet_leaf_74_csclk),
    .D(_0339_),
    .SET_B(net419),
    .Q(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6751_ (.CLK(clknet_leaf_75_csclk),
    .D(net1456),
    .RESET_B(net419),
    .Q(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6752_ (.CLK(clknet_leaf_74_csclk),
    .D(net1211),
    .RESET_B(net420),
    .Q(\gpio_configure[20][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6753_ (.CLK(clknet_leaf_70_csclk),
    .D(net1683),
    .RESET_B(net422),
    .Q(\gpio_configure[33][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6754_ (.CLK(clknet_leaf_73_csclk),
    .D(net960),
    .RESET_B(net422),
    .Q(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__dfstp_2 _6755_ (.CLK(clknet_leaf_70_csclk),
    .D(net1553),
    .SET_B(net423),
    .Q(\gpio_configure[33][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6756_ (.CLK(clknet_leaf_70_csclk),
    .D(net1551),
    .RESET_B(net423),
    .Q(\gpio_configure[33][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6757_ (.CLK(clknet_leaf_73_csclk),
    .D(net1294),
    .RESET_B(net423),
    .Q(\gpio_configure[33][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6758_ (.CLK(clknet_leaf_73_csclk),
    .D(net1674),
    .RESET_B(net420),
    .Q(\gpio_configure[21][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6759_ (.CLK(clknet_leaf_72_csclk),
    .D(net916),
    .RESET_B(net420),
    .Q(\gpio_configure[21][9] ));
 sky130_fd_sc_hd__dfstp_4 _6760_ (.CLK(clknet_leaf_73_csclk),
    .D(_0349_),
    .SET_B(net420),
    .Q(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6761_ (.CLK(clknet_leaf_73_csclk),
    .D(net1261),
    .RESET_B(net420),
    .Q(\gpio_configure[21][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6762_ (.CLK(clknet_leaf_74_csclk),
    .D(net1226),
    .RESET_B(net420),
    .Q(\gpio_configure[21][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6763_ (.CLK(clknet_leaf_0_csclk),
    .D(net1695),
    .RESET_B(net417),
    .Q(\gpio_configure[32][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6764_ (.CLK(clknet_leaf_0_csclk),
    .D(net1377),
    .RESET_B(net418),
    .Q(\gpio_configure[32][9] ));
 sky130_fd_sc_hd__dfstp_4 _6765_ (.CLK(clknet_leaf_0_csclk),
    .D(_0354_),
    .SET_B(net418),
    .Q(\gpio_configure[32][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6766_ (.CLK(clknet_leaf_0_csclk),
    .D(net1475),
    .RESET_B(net418),
    .Q(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6767_ (.CLK(clknet_leaf_3_csclk),
    .D(net1485),
    .RESET_B(net424),
    .Q(\gpio_configure[32][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6768_ (.CLK(clknet_leaf_73_csclk),
    .D(net1678),
    .RESET_B(net422),
    .Q(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6769_ (.CLK(clknet_leaf_73_csclk),
    .D(net964),
    .RESET_B(net422),
    .Q(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__dfstp_4 _6770_ (.CLK(clknet_leaf_70_csclk),
    .D(_0359_),
    .SET_B(net423),
    .Q(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6771_ (.CLK(clknet_leaf_73_csclk),
    .D(net1263),
    .RESET_B(net422),
    .Q(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6772_ (.CLK(clknet_leaf_73_csclk),
    .D(net1253),
    .RESET_B(net422),
    .Q(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6773_ (.CLK(clknet_leaf_0_csclk),
    .D(net1577),
    .RESET_B(net418),
    .Q(\gpio_configure[23][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6774_ (.CLK(clknet_leaf_0_csclk),
    .D(net1391),
    .RESET_B(net418),
    .Q(\gpio_configure[23][9] ));
 sky130_fd_sc_hd__dfstp_4 _6775_ (.CLK(clknet_leaf_3_csclk),
    .D(_0364_),
    .SET_B(net424),
    .Q(\gpio_configure[23][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6776_ (.CLK(clknet_leaf_0_csclk),
    .D(net1463),
    .RESET_B(net418),
    .Q(\gpio_configure[23][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6777_ (.CLK(clknet_leaf_2_csclk),
    .D(net1517),
    .RESET_B(net424),
    .Q(\gpio_configure[23][12] ));
 sky130_fd_sc_hd__dfrtp_2 _6778_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0367_),
    .RESET_B(net457),
    .Q(\wbbd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6779_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0368_),
    .RESET_B(net457),
    .Q(\wbbd_addr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6780_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0369_),
    .RESET_B(net458),
    .Q(\wbbd_addr[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6781_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0370_),
    .RESET_B(net458),
    .Q(\wbbd_addr[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6782_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0371_),
    .RESET_B(net458),
    .Q(\wbbd_addr[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6783_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0372_),
    .RESET_B(net458),
    .Q(\wbbd_addr[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6784_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0373_),
    .RESET_B(net458),
    .Q(\wbbd_addr[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6785_ (.CLK(clknet_leaf_74_csclk),
    .D(net1648),
    .RESET_B(net422),
    .Q(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6786_ (.CLK(clknet_leaf_1_csclk),
    .D(net1364),
    .RESET_B(net422),
    .Q(\gpio_configure[30][9] ));
 sky130_fd_sc_hd__dfstp_4 _6787_ (.CLK(clknet_leaf_74_csclk),
    .D(_0376_),
    .SET_B(net422),
    .Q(\gpio_configure[30][10] ));
 sky130_fd_sc_hd__dfrtp_2 _6788_ (.CLK(clknet_leaf_74_csclk),
    .D(net1433),
    .RESET_B(net422),
    .Q(\gpio_configure[30][11] ));
 sky130_fd_sc_hd__dfrtp_2 _6789_ (.CLK(clknet_leaf_74_csclk),
    .D(net1196),
    .RESET_B(net422),
    .Q(\gpio_configure[30][12] ));
 sky130_fd_sc_hd__dfrtn_1 _6790_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0379_),
    .RESET_B(_0057_),
    .Q(\hkspi.ldata[0] ));
 sky130_fd_sc_hd__dfrtn_1 _6791_ (.CLK_N(clknet_2_0_0_mgmt_gpio_in[4]),
    .D(_0380_),
    .RESET_B(_0058_),
    .Q(\hkspi.ldata[1] ));
 sky130_fd_sc_hd__dfrtn_1 _6792_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0381_),
    .RESET_B(_0059_),
    .Q(\hkspi.ldata[2] ));
 sky130_fd_sc_hd__dfrtn_1 _6793_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0382_),
    .RESET_B(_0060_),
    .Q(\hkspi.ldata[3] ));
 sky130_fd_sc_hd__dfrtn_1 _6794_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0383_),
    .RESET_B(_0061_),
    .Q(\hkspi.ldata[4] ));
 sky130_fd_sc_hd__dfrtn_1 _6795_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0384_),
    .RESET_B(_0062_),
    .Q(\hkspi.ldata[5] ));
 sky130_fd_sc_hd__dfrtn_1 _6796_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0385_),
    .RESET_B(_0063_),
    .Q(\hkspi.ldata[6] ));
 sky130_fd_sc_hd__dfrtn_1 _6797_ (.CLK_N(clknet_2_2_0_mgmt_gpio_in[4]),
    .D(_0386_),
    .RESET_B(_0064_),
    .Q(\hkspi.SDO ));
 sky130_fd_sc_hd__dfrtp_2 _6798_ (.CLK(clknet_leaf_77_csclk),
    .D(net1670),
    .RESET_B(net414),
    .Q(net271));
 sky130_fd_sc_hd__dfstp_4 _6799_ (.CLK(clknet_leaf_76_csclk),
    .D(_0388_),
    .SET_B(net414),
    .Q(net265));
 sky130_fd_sc_hd__dfrtp_2 _6800_ (.CLK(clknet_leaf_76_csclk),
    .D(net1659),
    .RESET_B(net414),
    .Q(net266));
 sky130_fd_sc_hd__dfrtp_2 _6801_ (.CLK(clknet_leaf_76_csclk),
    .D(net1395),
    .RESET_B(net414),
    .Q(net267));
 sky130_fd_sc_hd__dfstp_4 _6802_ (.CLK(clknet_leaf_76_csclk),
    .D(_0391_),
    .SET_B(net414),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_2 _6803_ (.CLK(clknet_leaf_76_csclk),
    .D(net1477),
    .RESET_B(net414),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_2 _6804_ (.CLK(clknet_leaf_76_csclk),
    .D(net1286),
    .RESET_B(net414),
    .Q(net270));
 sky130_fd_sc_hd__dfrtp_2 _6805_ (.CLK(clknet_leaf_75_csclk),
    .D(net1652),
    .RESET_B(net414),
    .Q(net272));
 sky130_fd_sc_hd__dfstp_4 _6806_ (.CLK(clknet_leaf_75_csclk),
    .D(_0395_),
    .SET_B(net414),
    .Q(net273));
 sky130_fd_sc_hd__dfrtp_2 _6807_ (.CLK(clknet_leaf_75_csclk),
    .D(net1489),
    .RESET_B(net419),
    .Q(net274));
 sky130_fd_sc_hd__dfrtp_2 _6808_ (.CLK(clknet_leaf_75_csclk),
    .D(net1443),
    .RESET_B(net419),
    .Q(net261));
 sky130_fd_sc_hd__dfstp_4 _6809_ (.CLK(clknet_leaf_75_csclk),
    .D(_0398_),
    .SET_B(net419),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_2 _6810_ (.CLK(clknet_leaf_75_csclk),
    .D(net1068),
    .RESET_B(net419),
    .Q(net263));
 sky130_fd_sc_hd__dfstp_2 _6811_ (.CLK(clknet_leaf_71_csclk),
    .D(net1634),
    .SET_B(net421),
    .Q(net282));
 sky130_fd_sc_hd__dfstp_4 _6812_ (.CLK(clknet_leaf_59_csclk),
    .D(_0401_),
    .SET_B(net429),
    .Q(net283));
 sky130_fd_sc_hd__dfstp_4 _6813_ (.CLK(clknet_leaf_59_csclk),
    .D(_0402_),
    .SET_B(net429),
    .Q(net284));
 sky130_fd_sc_hd__dfstp_2 _6814_ (.CLK(clknet_leaf_71_csclk),
    .D(net1366),
    .SET_B(net421),
    .Q(net285));
 sky130_fd_sc_hd__dfstp_2 _6815_ (.CLK(clknet_leaf_71_csclk),
    .D(net929),
    .SET_B(net429),
    .Q(net287));
 sky130_fd_sc_hd__dfstp_4 _6816_ (.CLK(clknet_leaf_57_csclk),
    .D(_0405_),
    .SET_B(net432),
    .Q(net288));
 sky130_fd_sc_hd__dfstp_4 _6817_ (.CLK(clknet_leaf_57_csclk),
    .D(_0406_),
    .SET_B(net432),
    .Q(net289));
 sky130_fd_sc_hd__dfstp_4 _6818_ (.CLK(clknet_leaf_57_csclk),
    .D(_0407_),
    .SET_B(net428),
    .Q(net290));
 sky130_fd_sc_hd__dfstp_2 _6819_ (.CLK(clknet_leaf_59_csclk),
    .D(_0408_),
    .SET_B(net429),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_2 _6820_ (.CLK(clknet_leaf_52_csclk),
    .D(net1536),
    .RESET_B(net433),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_2 _6821_ (.CLK(clknet_leaf_52_csclk),
    .D(net816),
    .RESET_B(net433),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_2 _6822_ (.CLK(clknet_leaf_52_csclk),
    .D(_0411_),
    .RESET_B(net433),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_2 _6823_ (.CLK(clknet_leaf_52_csclk),
    .D(net641),
    .RESET_B(net433),
    .Q(net304));
 sky130_fd_sc_hd__dfrtp_4 _6824_ (.CLK(clknet_leaf_77_csclk),
    .D(net1663),
    .RESET_B(net415),
    .Q(reset_reg));
 sky130_fd_sc_hd__dfrtp_2 _6825_ (.CLK(clknet_leaf_71_csclk),
    .D(net1596),
    .RESET_B(net429),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_2 _6826_ (.CLK(clknet_leaf_52_csclk),
    .D(net632),
    .RESET_B(net433),
    .Q(serial_bb_clock));
 sky130_fd_sc_hd__dfrtp_2 _6827_ (.CLK(clknet_leaf_52_csclk),
    .D(net599),
    .RESET_B(net433),
    .Q(serial_bb_load));
 sky130_fd_sc_hd__dfrtp_2 _6828_ (.CLK(clknet_leaf_52_csclk),
    .D(net1167),
    .RESET_B(net432),
    .Q(serial_bb_resetn));
 sky130_fd_sc_hd__dfrtp_2 _6829_ (.CLK(clknet_leaf_52_csclk),
    .D(net1038),
    .RESET_B(net432),
    .Q(serial_bb_data_1));
 sky130_fd_sc_hd__dfrtp_2 _6830_ (.CLK(clknet_leaf_52_csclk),
    .D(net1135),
    .RESET_B(net432),
    .Q(serial_bb_data_2));
 sky130_fd_sc_hd__dfrtp_2 _6831_ (.CLK(clknet_leaf_52_csclk),
    .D(net821),
    .RESET_B(net433),
    .Q(serial_bb_enable));
 sky130_fd_sc_hd__dfrtp_2 _6832_ (.CLK(clknet_leaf_54_csclk),
    .D(net1661),
    .RESET_B(net433),
    .Q(serial_xfer));
 sky130_fd_sc_hd__dfrtp_2 _6833_ (.CLK(clknet_leaf_22_csclk),
    .D(net1646),
    .RESET_B(net456),
    .Q(hkspi_disable));
 sky130_fd_sc_hd__dfrtp_2 _6834_ (.CLK(clknet_leaf_25_csclk),
    .D(net1188),
    .RESET_B(net444),
    .Q(clk1_output_dest));
 sky130_fd_sc_hd__dfrtp_2 _6835_ (.CLK(clknet_leaf_25_csclk),
    .D(net888),
    .RESET_B(net444),
    .Q(clk2_output_dest));
 sky130_fd_sc_hd__dfrtp_2 _6836_ (.CLK(clknet_leaf_25_csclk),
    .D(net1530),
    .RESET_B(net444),
    .Q(trap_output_dest));
 sky130_fd_sc_hd__dfrtp_2 _6837_ (.CLK(clknet_leaf_78_csclk),
    .D(net1687),
    .RESET_B(net417),
    .Q(irq_1_inputsrc));
 sky130_fd_sc_hd__dfrtp_2 _6838_ (.CLK(clknet_leaf_78_csclk),
    .D(net1399),
    .RESET_B(net417),
    .Q(irq_2_inputsrc));
 sky130_fd_sc_hd__dfrtp_2 _6839_ (.CLK(clknet_leaf_3_csclk),
    .D(net1672),
    .RESET_B(net425),
    .Q(\mgmt_gpio_data[32] ));
 sky130_fd_sc_hd__dfrtp_2 _6840_ (.CLK(clknet_leaf_3_csclk),
    .D(net954),
    .RESET_B(net425),
    .Q(\mgmt_gpio_data[33] ));
 sky130_fd_sc_hd__dfrtp_2 _6841_ (.CLK(clknet_leaf_35_csclk),
    .D(net1004),
    .RESET_B(net453),
    .Q(net240));
 sky130_fd_sc_hd__dfrtp_2 _6842_ (.CLK(clknet_leaf_0_csclk),
    .D(net1473),
    .RESET_B(net425),
    .Q(\mgmt_gpio_data[35] ));
 sky130_fd_sc_hd__dfrtp_2 _6843_ (.CLK(clknet_leaf_14_csclk),
    .D(net1343),
    .RESET_B(net441),
    .Q(\mgmt_gpio_data[36] ));
 sky130_fd_sc_hd__dfrtp_2 _6844_ (.CLK(clknet_leaf_17_csclk),
    .D(net558),
    .RESET_B(net441),
    .Q(\mgmt_gpio_data[37] ));
 sky130_fd_sc_hd__dfrtp_1 _6845_ (.CLK(clknet_leaf_78_csclk),
    .D(net1426),
    .RESET_B(net416),
    .Q(\mgmt_gpio_data_buf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6846_ (.CLK(clknet_leaf_0_csclk),
    .D(net1375),
    .RESET_B(net423),
    .Q(\mgmt_gpio_data_buf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6847_ (.CLK(clknet_leaf_51_csclk),
    .D(net1150),
    .RESET_B(net434),
    .Q(\mgmt_gpio_data_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6848_ (.CLK(clknet_leaf_51_csclk),
    .D(net679),
    .RESET_B(net434),
    .Q(\mgmt_gpio_data_buf[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6849_ (.CLK(clknet_leaf_48_csclk),
    .D(net756),
    .RESET_B(net438),
    .Q(\mgmt_gpio_data_buf[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6850_ (.CLK(clknet_leaf_47_csclk),
    .D(net1163),
    .RESET_B(net438),
    .Q(\mgmt_gpio_data_buf[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6851_ (.CLK(clknet_leaf_0_csclk),
    .D(net709),
    .RESET_B(net417),
    .Q(\mgmt_gpio_data_buf[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6852_ (.CLK(clknet_leaf_51_csclk),
    .D(net892),
    .RESET_B(net434),
    .Q(\mgmt_gpio_data_buf[7] ));
 sky130_fd_sc_hd__dfstp_4 _6853_ (.CLK(clknet_leaf_56_csclk),
    .D(_0442_),
    .SET_B(net430),
    .Q(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__dfstp_2 _6854_ (.CLK(clknet_leaf_62_csclk),
    .D(net858),
    .SET_B(net430),
    .Q(\gpio_configure[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6855_ (.CLK(clknet_leaf_43_csclk),
    .D(net1219),
    .RESET_B(net437),
    .Q(\gpio_configure[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6856_ (.CLK(clknet_leaf_56_csclk),
    .D(net661),
    .RESET_B(net428),
    .Q(\gpio_configure[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6857_ (.CLK(clknet_leaf_43_csclk),
    .D(net740),
    .RESET_B(net437),
    .Q(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6858_ (.CLK(clknet_leaf_46_csclk),
    .D(net1112),
    .RESET_B(net438),
    .Q(\gpio_configure[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6859_ (.CLK(clknet_leaf_53_csclk),
    .D(net1169),
    .RESET_B(net432),
    .Q(\gpio_configure[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6860_ (.CLK(clknet_leaf_45_csclk),
    .D(net571),
    .RESET_B(net438),
    .Q(\gpio_configure[0][7] ));
 sky130_fd_sc_hd__dfstp_4 _6861_ (.CLK(clknet_leaf_30_csclk),
    .D(_0450_),
    .SET_B(net448),
    .Q(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__dfstp_4 _6862_ (.CLK(clknet_leaf_29_csclk),
    .D(_0451_),
    .SET_B(net446),
    .Q(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6863_ (.CLK(clknet_leaf_29_csclk),
    .D(net1548),
    .RESET_B(net449),
    .Q(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6864_ (.CLK(clknet_leaf_31_csclk),
    .D(net634),
    .RESET_B(net452),
    .Q(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6865_ (.CLK(clknet_leaf_29_csclk),
    .D(net1083),
    .RESET_B(net449),
    .Q(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6866_ (.CLK(clknet_leaf_33_csclk),
    .D(net541),
    .RESET_B(net452),
    .Q(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6867_ (.CLK(clknet_leaf_46_csclk),
    .D(net719),
    .RESET_B(net438),
    .Q(\gpio_configure[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6868_ (.CLK(clknet_leaf_44_csclk),
    .D(net492),
    .RESET_B(net437),
    .Q(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__dfstp_4 _6869_ (.CLK(clknet_leaf_28_csclk),
    .D(_0458_),
    .SET_B(net447),
    .Q(\gpio_configure[2][0] ));
 sky130_fd_sc_hd__dfstp_4 _6870_ (.CLK(clknet_leaf_17_csclk),
    .D(_0459_),
    .SET_B(net441),
    .Q(\gpio_configure[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6871_ (.CLK(clknet_leaf_19_csclk),
    .D(net1623),
    .RESET_B(net444),
    .Q(\gpio_configure[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6872_ (.CLK(clknet_leaf_40_csclk),
    .D(_0461_),
    .RESET_B(net443),
    .Q(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6873_ (.CLK(clknet_leaf_19_csclk),
    .D(net1318),
    .RESET_B(net441),
    .Q(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6874_ (.CLK(clknet_leaf_40_csclk),
    .D(net727),
    .RESET_B(net443),
    .Q(\gpio_configure[2][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6875_ (.CLK(clknet_leaf_39_csclk),
    .D(net1230),
    .RESET_B(net450),
    .Q(\gpio_configure[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6876_ (.CLK(clknet_leaf_42_csclk),
    .D(net982),
    .RESET_B(net443),
    .Q(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__dfstp_4 _6877_ (.CLK(clknet_leaf_18_csclk),
    .D(_0466_),
    .SET_B(net449),
    .Q(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6878_ (.CLK(clknet_leaf_17_csclk),
    .D(net1050),
    .RESET_B(net441),
    .Q(\gpio_configure[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6879_ (.CLK(clknet_leaf_18_csclk),
    .D(net1611),
    .RESET_B(net449),
    .Q(\gpio_configure[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6880_ (.CLK(clknet_leaf_35_csclk),
    .D(_0469_),
    .RESET_B(net453),
    .Q(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6881_ (.CLK(clknet_leaf_17_csclk),
    .D(net1306),
    .RESET_B(net441),
    .Q(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6882_ (.CLK(clknet_leaf_34_csclk),
    .D(net856),
    .RESET_B(net453),
    .Q(\gpio_configure[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6883_ (.CLK(clknet_leaf_35_csclk),
    .D(net1062),
    .RESET_B(net453),
    .Q(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6884_ (.CLK(clknet_leaf_32_csclk),
    .D(net840),
    .RESET_B(net447),
    .Q(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__dfstp_4 _6885_ (.CLK(clknet_leaf_26_csclk),
    .D(_0474_),
    .SET_B(net444),
    .Q(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__dfstp_4 _6886_ (.CLK(clknet_leaf_27_csclk),
    .D(_0475_),
    .SET_B(net444),
    .Q(\gpio_configure[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6887_ (.CLK(clknet_leaf_19_csclk),
    .D(net1408),
    .RESET_B(net444),
    .Q(\gpio_configure[4][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6888_ (.CLK(clknet_leaf_37_csclk),
    .D(_0477_),
    .RESET_B(net450),
    .Q(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6889_ (.CLK(clknet_leaf_19_csclk),
    .D(net1314),
    .RESET_B(net444),
    .Q(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6890_ (.CLK(clknet_leaf_33_csclk),
    .D(net931),
    .RESET_B(net451),
    .Q(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6891_ (.CLK(clknet_leaf_37_csclk),
    .D(net1002),
    .RESET_B(net450),
    .Q(\gpio_configure[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6892_ (.CLK(clknet_leaf_32_csclk),
    .D(net829),
    .RESET_B(net444),
    .Q(\gpio_configure[4][7] ));
 sky130_fd_sc_hd__dfstp_4 _6893_ (.CLK(clknet_leaf_30_csclk),
    .D(_0482_),
    .SET_B(net448),
    .Q(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__dfstp_4 _6894_ (.CLK(clknet_leaf_19_csclk),
    .D(_0483_),
    .SET_B(net441),
    .Q(\gpio_configure[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6895_ (.CLK(clknet_leaf_18_csclk),
    .D(net1599),
    .RESET_B(net449),
    .Q(\gpio_configure[5][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6896_ (.CLK(clknet_leaf_37_csclk),
    .D(_0485_),
    .RESET_B(net450),
    .Q(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6897_ (.CLK(clknet_leaf_17_csclk),
    .D(net1290),
    .RESET_B(net441),
    .Q(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6898_ (.CLK(clknet_leaf_38_csclk),
    .D(net1015),
    .RESET_B(net451),
    .Q(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6899_ (.CLK(clknet_leaf_35_csclk),
    .D(net1122),
    .RESET_B(net453),
    .Q(\gpio_configure[5][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6900_ (.CLK(clknet_leaf_32_csclk),
    .D(net849),
    .RESET_B(net444),
    .Q(\gpio_configure[5][7] ));
 sky130_fd_sc_hd__dfstp_4 _6901_ (.CLK(clknet_leaf_25_csclk),
    .D(_0490_),
    .SET_B(net445),
    .Q(\gpio_configure[6][0] ));
 sky130_fd_sc_hd__dfstp_4 _6902_ (.CLK(clknet_leaf_20_csclk),
    .D(_0491_),
    .SET_B(net444),
    .Q(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6903_ (.CLK(clknet_leaf_19_csclk),
    .D(net1619),
    .RESET_B(net444),
    .Q(\gpio_configure[6][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6904_ (.CLK(clknet_leaf_38_csclk),
    .D(net1241),
    .RESET_B(net450),
    .Q(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6905_ (.CLK(clknet_leaf_20_csclk),
    .D(net907),
    .RESET_B(net442),
    .Q(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6906_ (.CLK(clknet_leaf_39_csclk),
    .D(net1044),
    .RESET_B(net451),
    .Q(\gpio_configure[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6907_ (.CLK(clknet_leaf_38_csclk),
    .D(net1200),
    .RESET_B(net450),
    .Q(\gpio_configure[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6908_ (.CLK(clknet_leaf_25_csclk),
    .D(net992),
    .RESET_B(net445),
    .Q(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__dfstp_4 _6909_ (.CLK(clknet_leaf_26_csclk),
    .D(_0498_),
    .SET_B(net445),
    .Q(\gpio_configure[7][0] ));
 sky130_fd_sc_hd__dfstp_4 _6910_ (.CLK(clknet_leaf_28_csclk),
    .D(net778),
    .SET_B(net446),
    .Q(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6911_ (.CLK(clknet_leaf_28_csclk),
    .D(net974),
    .RESET_B(net446),
    .Q(\gpio_configure[7][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6912_ (.CLK(clknet_leaf_37_csclk),
    .D(net1036),
    .RESET_B(net450),
    .Q(\gpio_configure[7][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6913_ (.CLK(clknet_leaf_28_csclk),
    .D(net1198),
    .RESET_B(net446),
    .Q(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6914_ (.CLK(clknet_leaf_33_csclk),
    .D(net912),
    .RESET_B(net451),
    .Q(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6915_ (.CLK(clknet_leaf_33_csclk),
    .D(net1048),
    .RESET_B(net450),
    .Q(\gpio_configure[7][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6916_ (.CLK(clknet_leaf_32_csclk),
    .D(net810),
    .RESET_B(net447),
    .Q(\gpio_configure[7][7] ));
 sky130_fd_sc_hd__dfstp_4 _6917_ (.CLK(clknet_leaf_29_csclk),
    .D(_0506_),
    .SET_B(net447),
    .Q(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__dfstp_4 _6918_ (.CLK(clknet_leaf_17_csclk),
    .D(_0507_),
    .SET_B(net442),
    .Q(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6919_ (.CLK(clknet_leaf_17_csclk),
    .D(net1615),
    .RESET_B(net442),
    .Q(\gpio_configure[8][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6920_ (.CLK(clknet_leaf_33_csclk),
    .D(net1126),
    .RESET_B(net452),
    .Q(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6921_ (.CLK(clknet_leaf_17_csclk),
    .D(net1300),
    .RESET_B(net442),
    .Q(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6922_ (.CLK(clknet_leaf_34_csclk),
    .D(net867),
    .RESET_B(net452),
    .Q(\gpio_configure[8][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6923_ (.CLK(clknet_leaf_33_csclk),
    .D(net1052),
    .RESET_B(net452),
    .Q(\gpio_configure[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6924_ (.CLK(clknet_leaf_31_csclk),
    .D(net800),
    .RESET_B(net452),
    .Q(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__dfstp_4 _6925_ (.CLK(clknet_leaf_29_csclk),
    .D(_0514_),
    .SET_B(net448),
    .Q(\gpio_configure[9][0] ));
 sky130_fd_sc_hd__dfstp_4 _6926_ (.CLK(clknet_leaf_28_csclk),
    .D(_0515_),
    .SET_B(net446),
    .Q(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6927_ (.CLK(clknet_leaf_18_csclk),
    .D(net1586),
    .RESET_B(net446),
    .Q(\gpio_configure[9][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6928_ (.CLK(clknet_leaf_34_csclk),
    .D(net1054),
    .RESET_B(net453),
    .Q(\gpio_configure[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6929_ (.CLK(clknet_leaf_18_csclk),
    .D(net764),
    .RESET_B(net449),
    .Q(\gpio_configure[9][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6930_ (.CLK(clknet_leaf_34_csclk),
    .D(net837),
    .RESET_B(net452),
    .Q(\gpio_configure[9][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6931_ (.CLK(clknet_leaf_34_csclk),
    .D(net1008),
    .RESET_B(net453),
    .Q(\gpio_configure[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6932_ (.CLK(clknet_leaf_30_csclk),
    .D(net798),
    .RESET_B(net448),
    .Q(\gpio_configure[9][7] ));
 sky130_fd_sc_hd__dfstp_4 _6933_ (.CLK(clknet_leaf_26_csclk),
    .D(_0522_),
    .SET_B(net445),
    .Q(\gpio_configure[10][0] ));
 sky130_fd_sc_hd__dfstp_4 _6934_ (.CLK(clknet_leaf_28_csclk),
    .D(_0523_),
    .SET_B(net447),
    .Q(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6935_ (.CLK(clknet_leaf_17_csclk),
    .D(net1609),
    .RESET_B(net442),
    .Q(\gpio_configure[10][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6936_ (.CLK(clknet_leaf_38_csclk),
    .D(_0525_),
    .RESET_B(net450),
    .Q(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6937_ (.CLK(clknet_leaf_17_csclk),
    .D(net1308),
    .RESET_B(net442),
    .Q(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6938_ (.CLK(clknet_leaf_33_csclk),
    .D(net905),
    .RESET_B(net451),
    .Q(\gpio_configure[10][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6939_ (.CLK(clknet_leaf_35_csclk),
    .D(net1087),
    .RESET_B(net454),
    .Q(\gpio_configure[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6940_ (.CLK(clknet_leaf_24_csclk),
    .D(net1056),
    .RESET_B(net443),
    .Q(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__dfstp_4 _6941_ (.CLK(clknet_leaf_57_csclk),
    .D(_0530_),
    .SET_B(net428),
    .Q(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__dfstp_4 _6942_ (.CLK(clknet_leaf_57_csclk),
    .D(_0531_),
    .SET_B(net428),
    .Q(\gpio_configure[11][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6943_ (.CLK(clknet_leaf_59_csclk),
    .D(net506),
    .RESET_B(net429),
    .Q(\gpio_configure[11][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6944_ (.CLK(clknet_leaf_47_csclk),
    .D(net725),
    .RESET_B(net438),
    .Q(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6945_ (.CLK(clknet_leaf_59_csclk),
    .D(net700),
    .RESET_B(net429),
    .Q(\gpio_configure[11][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6946_ (.CLK(clknet_leaf_48_csclk),
    .D(net1173),
    .RESET_B(net438),
    .Q(\gpio_configure[11][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6947_ (.CLK(clknet_leaf_51_csclk),
    .D(net1085),
    .RESET_B(net434),
    .Q(\gpio_configure[11][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6948_ (.CLK(clknet_leaf_56_csclk),
    .D(net861),
    .RESET_B(net430),
    .Q(\gpio_configure[11][7] ));
 sky130_fd_sc_hd__dfstp_4 _6949_ (.CLK(clknet_leaf_27_csclk),
    .D(_0538_),
    .SET_B(net445),
    .Q(\gpio_configure[12][0] ));
 sky130_fd_sc_hd__dfstp_4 _6950_ (.CLK(clknet_leaf_21_csclk),
    .D(_0539_),
    .SET_B(net442),
    .Q(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6951_ (.CLK(clknet_leaf_21_csclk),
    .D(net1644),
    .RESET_B(net442),
    .Q(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6952_ (.CLK(clknet_leaf_38_csclk),
    .D(net1259),
    .RESET_B(net450),
    .Q(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6953_ (.CLK(clknet_leaf_19_csclk),
    .D(net1312),
    .RESET_B(net442),
    .Q(\gpio_configure[12][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6954_ (.CLK(clknet_leaf_39_csclk),
    .D(net1025),
    .RESET_B(net451),
    .Q(\gpio_configure[12][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6955_ (.CLK(clknet_leaf_38_csclk),
    .D(net1215),
    .RESET_B(net450),
    .Q(\gpio_configure[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6956_ (.CLK(clknet_leaf_25_csclk),
    .D(net962),
    .RESET_B(net443),
    .Q(\gpio_configure[12][7] ));
 sky130_fd_sc_hd__dfstp_2 _6957_ (.CLK(clknet_leaf_42_csclk),
    .D(net1348),
    .SET_B(net443),
    .Q(\gpio_configure[13][0] ));
 sky130_fd_sc_hd__dfstp_4 _6958_ (.CLK(clknet_leaf_26_csclk),
    .D(_0547_),
    .SET_B(net445),
    .Q(\gpio_configure[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6959_ (.CLK(clknet_leaf_20_csclk),
    .D(net1650),
    .RESET_B(net444),
    .Q(\gpio_configure[13][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6960_ (.CLK(clknet_leaf_39_csclk),
    .D(net758),
    .RESET_B(net443),
    .Q(\gpio_configure[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6961_ (.CLK(clknet_leaf_23_csclk),
    .D(net896),
    .RESET_B(net443),
    .Q(\gpio_configure[13][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6962_ (.CLK(clknet_leaf_39_csclk),
    .D(net1042),
    .RESET_B(net451),
    .Q(\gpio_configure[13][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6963_ (.CLK(clknet_leaf_42_csclk),
    .D(net754),
    .RESET_B(net443),
    .Q(\gpio_configure[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6964_ (.CLK(clknet_leaf_25_csclk),
    .D(net564),
    .RESET_B(net451),
    .Q(\gpio_configure[13][7] ));
 sky130_fd_sc_hd__dfstp_4 _6965_ (.CLK(clknet_leaf_26_csclk),
    .D(_0554_),
    .SET_B(net445),
    .Q(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__dfstp_4 _6966_ (.CLK(clknet_leaf_27_csclk),
    .D(net796),
    .SET_B(net444),
    .Q(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6967_ (.CLK(clknet_leaf_27_csclk),
    .D(net1013),
    .RESET_B(net444),
    .Q(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6968_ (.CLK(clknet_leaf_33_csclk),
    .D(net1093),
    .RESET_B(net451),
    .Q(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6969_ (.CLK(clknet_leaf_27_csclk),
    .D(net746),
    .RESET_B(net444),
    .Q(\gpio_configure[14][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6970_ (.CLK(clknet_leaf_33_csclk),
    .D(net939),
    .RESET_B(net451),
    .Q(\gpio_configure[14][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6971_ (.CLK(clknet_leaf_39_csclk),
    .D(net1209),
    .RESET_B(net451),
    .Q(\gpio_configure[14][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6972_ (.CLK(clknet_leaf_32_csclk),
    .D(net831),
    .RESET_B(net451),
    .Q(\gpio_configure[14][7] ));
 sky130_fd_sc_hd__dfstp_4 _6973_ (.CLK(clknet_leaf_23_csclk),
    .D(_0562_),
    .SET_B(net443),
    .Q(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__dfstp_4 _6974_ (.CLK(clknet_leaf_27_csclk),
    .D(_0563_),
    .SET_B(net444),
    .Q(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6975_ (.CLK(clknet_leaf_24_csclk),
    .D(net1247),
    .RESET_B(net443),
    .Q(\gpio_configure[15][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6976_ (.CLK(clknet_leaf_38_csclk),
    .D(net1245),
    .RESET_B(net450),
    .Q(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6977_ (.CLK(clknet_leaf_23_csclk),
    .D(net941),
    .RESET_B(net443),
    .Q(\gpio_configure[15][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6978_ (.CLK(clknet_leaf_42_csclk),
    .D(net650),
    .RESET_B(net443),
    .Q(\gpio_configure[15][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6979_ (.CLK(clknet_leaf_47_csclk),
    .D(net723),
    .RESET_B(net438),
    .Q(\gpio_configure[15][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6980_ (.CLK(clknet_leaf_42_csclk),
    .D(net956),
    .RESET_B(net443),
    .Q(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__dfstp_4 _6981_ (.CLK(clknet_leaf_30_csclk),
    .D(_0570_),
    .SET_B(net447),
    .Q(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__dfstp_4 _6982_ (.CLK(clknet_leaf_28_csclk),
    .D(_0571_),
    .SET_B(net447),
    .Q(\gpio_configure[16][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6983_ (.CLK(clknet_leaf_28_csclk),
    .D(net978),
    .RESET_B(net446),
    .Q(\gpio_configure[16][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6984_ (.CLK(clknet_leaf_37_csclk),
    .D(net1080),
    .RESET_B(net451),
    .Q(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6985_ (.CLK(clknet_leaf_27_csclk),
    .D(net742),
    .RESET_B(net446),
    .Q(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6986_ (.CLK(clknet_leaf_34_csclk),
    .D(net872),
    .RESET_B(net452),
    .Q(\gpio_configure[16][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6987_ (.CLK(clknet_leaf_37_csclk),
    .D(net1023),
    .RESET_B(net453),
    .Q(\gpio_configure[16][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6988_ (.CLK(clknet_leaf_32_csclk),
    .D(net833),
    .RESET_B(net452),
    .Q(\gpio_configure[16][7] ));
 sky130_fd_sc_hd__dfstp_4 _6989_ (.CLK(clknet_leaf_62_csclk),
    .D(_0578_),
    .SET_B(net430),
    .Q(\gpio_configure[17][0] ));
 sky130_fd_sc_hd__dfstp_2 _6990_ (.CLK(clknet_leaf_63_csclk),
    .D(_0579_),
    .SET_B(net436),
    .Q(\gpio_configure[17][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6991_ (.CLK(clknet_leaf_60_csclk),
    .D(net1139),
    .RESET_B(net431),
    .Q(\gpio_configure[17][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6992_ (.CLK(clknet_leaf_51_csclk),
    .D(_0581_),
    .RESET_B(net434),
    .Q(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6993_ (.CLK(clknet_leaf_60_csclk),
    .D(net693),
    .RESET_B(net431),
    .Q(\gpio_configure[17][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6994_ (.CLK(clknet_leaf_48_csclk),
    .D(net580),
    .RESET_B(net438),
    .Q(\gpio_configure[17][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6995_ (.CLK(clknet_leaf_48_csclk),
    .D(net1237),
    .RESET_B(net434),
    .Q(\gpio_configure[17][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6996_ (.CLK(clknet_leaf_55_csclk),
    .D(net945),
    .RESET_B(net434),
    .Q(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__dfstp_4 _6997_ (.CLK(clknet_leaf_58_csclk),
    .D(_0586_),
    .SET_B(net428),
    .Q(\gpio_configure[18][0] ));
 sky130_fd_sc_hd__dfstp_4 _6998_ (.CLK(clknet_leaf_59_csclk),
    .D(net814),
    .SET_B(net429),
    .Q(\gpio_configure[18][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6999_ (.CLK(clknet_leaf_59_csclk),
    .D(net511),
    .RESET_B(net429),
    .Q(\gpio_configure[18][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7000_ (.CLK(clknet_leaf_31_csclk),
    .D(_0589_),
    .RESET_B(net452),
    .Q(\gpio_configure[18][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7001_ (.CLK(clknet_leaf_18_csclk),
    .D(net766),
    .RESET_B(net446),
    .Q(\gpio_configure[18][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7002_ (.CLK(clknet_leaf_53_csclk),
    .D(net1033),
    .RESET_B(net432),
    .Q(\gpio_configure[18][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7003_ (.CLK(clknet_leaf_33_csclk),
    .D(_0592_),
    .RESET_B(net452),
    .Q(\gpio_configure[18][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7004_ (.CLK(clknet_leaf_32_csclk),
    .D(net843),
    .RESET_B(net445),
    .Q(\gpio_configure[18][7] ));
 sky130_fd_sc_hd__dfstp_4 _7005_ (.CLK(clknet_leaf_56_csclk),
    .D(_0594_),
    .SET_B(net430),
    .Q(\gpio_configure[19][0] ));
 sky130_fd_sc_hd__dfstp_2 _7006_ (.CLK(clknet_leaf_61_csclk),
    .D(_0595_),
    .SET_B(net430),
    .Q(\gpio_configure[19][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7007_ (.CLK(clknet_leaf_60_csclk),
    .D(net1180),
    .RESET_B(net431),
    .Q(\gpio_configure[19][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7008_ (.CLK(clknet_leaf_50_csclk),
    .D(net721),
    .RESET_B(net434),
    .Q(\gpio_configure[19][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7009_ (.CLK(clknet_leaf_64_csclk),
    .D(net738),
    .RESET_B(net436),
    .Q(\gpio_configure[19][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7010_ (.CLK(clknet_leaf_45_csclk),
    .D(net601),
    .RESET_B(net438),
    .Q(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7011_ (.CLK(clknet_leaf_54_csclk),
    .D(net1159),
    .RESET_B(net434),
    .Q(\gpio_configure[19][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7012_ (.CLK(clknet_leaf_63_csclk),
    .D(net937),
    .RESET_B(net436),
    .Q(\gpio_configure[19][7] ));
 sky130_fd_sc_hd__dfstp_4 _7013_ (.CLK(clknet_leaf_60_csclk),
    .D(_0602_),
    .SET_B(net428),
    .Q(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__dfstp_2 _7014_ (.CLK(clknet_leaf_60_csclk),
    .D(_0603_),
    .SET_B(net430),
    .Q(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7015_ (.CLK(clknet_leaf_60_csclk),
    .D(net1128),
    .RESET_B(net431),
    .Q(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7016_ (.CLK(clknet_leaf_56_csclk),
    .D(net612),
    .RESET_B(net430),
    .Q(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7017_ (.CLK(clknet_leaf_60_csclk),
    .D(net652),
    .RESET_B(net429),
    .Q(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7018_ (.CLK(clknet_leaf_54_csclk),
    .D(net1095),
    .RESET_B(net434),
    .Q(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7019_ (.CLK(clknet_leaf_54_csclk),
    .D(net1148),
    .RESET_B(net434),
    .Q(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7020_ (.CLK(clknet_leaf_56_csclk),
    .D(net884),
    .RESET_B(net430),
    .Q(\gpio_configure[20][7] ));
 sky130_fd_sc_hd__dfstp_4 _7021_ (.CLK(clknet_leaf_58_csclk),
    .D(_0610_),
    .SET_B(net428),
    .Q(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__dfstp_2 _7022_ (.CLK(clknet_leaf_61_csclk),
    .D(_0611_),
    .SET_B(net430),
    .Q(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7023_ (.CLK(clknet_leaf_56_csclk),
    .D(net496),
    .RESET_B(net430),
    .Q(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7024_ (.CLK(clknet_leaf_62_csclk),
    .D(net691),
    .RESET_B(net430),
    .Q(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7025_ (.CLK(clknet_leaf_65_csclk),
    .D(net760),
    .RESET_B(net437),
    .Q(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7026_ (.CLK(clknet_leaf_46_csclk),
    .D(net1154),
    .RESET_B(net438),
    .Q(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7027_ (.CLK(clknet_leaf_54_csclk),
    .D(net1192),
    .RESET_B(net435),
    .Q(\gpio_configure[21][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7028_ (.CLK(clknet_leaf_55_csclk),
    .D(net935),
    .RESET_B(net434),
    .Q(\gpio_configure[21][7] ));
 sky130_fd_sc_hd__dfstp_4 _7029_ (.CLK(clknet_leaf_44_csclk),
    .D(_0618_),
    .SET_B(net436),
    .Q(\gpio_configure[22][0] ));
 sky130_fd_sc_hd__dfstp_4 _7030_ (.CLK(clknet_leaf_59_csclk),
    .D(_0619_),
    .SET_B(net429),
    .Q(\gpio_configure[22][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7031_ (.CLK(clknet_leaf_64_csclk),
    .D(net1239),
    .RESET_B(net436),
    .Q(\gpio_configure[22][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7032_ (.CLK(clknet_leaf_63_csclk),
    .D(net703),
    .RESET_B(net436),
    .Q(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7033_ (.CLK(clknet_leaf_64_csclk),
    .D(net1320),
    .RESET_B(net436),
    .Q(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7034_ (.CLK(clknet_leaf_53_csclk),
    .D(net1078),
    .RESET_B(net432),
    .Q(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7035_ (.CLK(clknet_leaf_52_csclk),
    .D(net1116),
    .RESET_B(net432),
    .Q(\gpio_configure[22][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7036_ (.CLK(clknet_leaf_57_csclk),
    .D(net869),
    .RESET_B(net428),
    .Q(\gpio_configure[22][7] ));
 sky130_fd_sc_hd__dfstp_4 _7037_ (.CLK(clknet_leaf_57_csclk),
    .D(_0626_),
    .SET_B(net428),
    .Q(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__dfstp_4 _7038_ (.CLK(clknet_leaf_58_csclk),
    .D(_0627_),
    .SET_B(net428),
    .Q(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7039_ (.CLK(clknet_leaf_59_csclk),
    .D(net1146),
    .RESET_B(net429),
    .Q(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7040_ (.CLK(clknet_leaf_56_csclk),
    .D(net659),
    .RESET_B(net432),
    .Q(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7041_ (.CLK(clknet_leaf_58_csclk),
    .D(net648),
    .RESET_B(net429),
    .Q(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7042_ (.CLK(clknet_leaf_53_csclk),
    .D(net1040),
    .RESET_B(net432),
    .Q(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7043_ (.CLK(clknet_leaf_53_csclk),
    .D(net1106),
    .RESET_B(net432),
    .Q(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7044_ (.CLK(clknet_leaf_57_csclk),
    .D(net886),
    .RESET_B(net428),
    .Q(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__dfstp_4 _7045_ (.CLK(clknet_leaf_62_csclk),
    .D(_0634_),
    .SET_B(net430),
    .Q(\gpio_configure[24][0] ));
 sky130_fd_sc_hd__dfstp_4 _7046_ (.CLK(clknet_leaf_61_csclk),
    .D(_0635_),
    .SET_B(net431),
    .Q(\gpio_configure[24][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7047_ (.CLK(clknet_leaf_60_csclk),
    .D(net1165),
    .RESET_B(net429),
    .Q(\gpio_configure[24][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7048_ (.CLK(clknet_leaf_55_csclk),
    .D(_0637_),
    .RESET_B(net434),
    .Q(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7049_ (.CLK(clknet_leaf_61_csclk),
    .D(net734),
    .RESET_B(net431),
    .Q(\gpio_configure[24][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7050_ (.CLK(clknet_leaf_46_csclk),
    .D(net1118),
    .RESET_B(net438),
    .Q(\gpio_configure[24][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7051_ (.CLK(clknet_leaf_55_csclk),
    .D(net1184),
    .RESET_B(net434),
    .Q(\gpio_configure[24][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7052_ (.CLK(clknet_leaf_44_csclk),
    .D(net968),
    .RESET_B(net436),
    .Q(\gpio_configure[24][7] ));
 sky130_fd_sc_hd__dfstp_4 _7053_ (.CLK(clknet_leaf_27_csclk),
    .D(_0642_),
    .SET_B(net445),
    .Q(\gpio_configure[25][0] ));
 sky130_fd_sc_hd__dfstp_4 _7054_ (.CLK(clknet_leaf_26_csclk),
    .D(_0643_),
    .SET_B(net445),
    .Q(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7055_ (.CLK(clknet_leaf_18_csclk),
    .D(net1401),
    .RESET_B(net446),
    .Q(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7056_ (.CLK(clknet_leaf_31_csclk),
    .D(net618),
    .RESET_B(net448),
    .Q(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7057_ (.CLK(clknet_leaf_19_csclk),
    .D(net1316),
    .RESET_B(net442),
    .Q(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7058_ (.CLK(clknet_leaf_33_csclk),
    .D(net919),
    .RESET_B(net454),
    .Q(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7059_ (.CLK(clknet_leaf_33_csclk),
    .D(net1060),
    .RESET_B(net451),
    .Q(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7060_ (.CLK(clknet_leaf_31_csclk),
    .D(net826),
    .RESET_B(net454),
    .Q(\gpio_configure[25][7] ));
 sky130_fd_sc_hd__dfstp_4 _7061_ (.CLK(clknet_leaf_58_csclk),
    .D(_0650_),
    .SET_B(net428),
    .Q(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__dfstp_4 _7062_ (.CLK(clknet_leaf_29_csclk),
    .D(net751),
    .SET_B(net446),
    .Q(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7063_ (.CLK(clknet_leaf_29_csclk),
    .D(net894),
    .RESET_B(net449),
    .Q(\gpio_configure[26][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7064_ (.CLK(clknet_leaf_31_csclk),
    .D(net626),
    .RESET_B(net454),
    .Q(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7065_ (.CLK(clknet_leaf_23_csclk),
    .D(net925),
    .RESET_B(net443),
    .Q(\gpio_configure[26][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7066_ (.CLK(clknet_leaf_34_csclk),
    .D(net865),
    .RESET_B(net454),
    .Q(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7067_ (.CLK(clknet_leaf_53_csclk),
    .D(net1156),
    .RESET_B(net432),
    .Q(\gpio_configure[26][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7068_ (.CLK(clknet_leaf_42_csclk),
    .D(net947),
    .RESET_B(net443),
    .Q(\gpio_configure[26][7] ));
 sky130_fd_sc_hd__dfstp_4 _7069_ (.CLK(clknet_leaf_63_csclk),
    .D(_0658_),
    .SET_B(net436),
    .Q(\gpio_configure[27][0] ));
 sky130_fd_sc_hd__dfstp_2 _7070_ (.CLK(clknet_leaf_63_csclk),
    .D(_0659_),
    .SET_B(net436),
    .Q(\gpio_configure[27][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7071_ (.CLK(clknet_leaf_63_csclk),
    .D(net556),
    .RESET_B(net436),
    .Q(\gpio_configure[27][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7072_ (.CLK(clknet_leaf_63_csclk),
    .D(_0661_),
    .RESET_B(net436),
    .Q(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7073_ (.CLK(clknet_leaf_63_csclk),
    .D(net711),
    .RESET_B(net436),
    .Q(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7074_ (.CLK(clknet_leaf_49_csclk),
    .D(net1228),
    .RESET_B(net438),
    .Q(\gpio_configure[27][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7075_ (.CLK(clknet_leaf_49_csclk),
    .D(net770),
    .RESET_B(net438),
    .Q(\gpio_configure[27][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7076_ (.CLK(clknet_leaf_44_csclk),
    .D(net949),
    .RESET_B(net438),
    .Q(\gpio_configure[27][7] ));
 sky130_fd_sc_hd__dfstp_4 _7077_ (.CLK(clknet_leaf_44_csclk),
    .D(_0666_),
    .SET_B(net436),
    .Q(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__dfstp_2 _7078_ (.CLK(clknet_leaf_61_csclk),
    .D(net878),
    .SET_B(net430),
    .Q(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7079_ (.CLK(clknet_leaf_65_csclk),
    .D(net620),
    .RESET_B(net437),
    .Q(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7080_ (.CLK(clknet_leaf_43_csclk),
    .D(net698),
    .RESET_B(net437),
    .Q(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7081_ (.CLK(clknet_leaf_65_csclk),
    .D(net762),
    .RESET_B(net437),
    .Q(\gpio_configure[28][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7082_ (.CLK(clknet_leaf_50_csclk),
    .D(net1133),
    .RESET_B(net435),
    .Q(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7083_ (.CLK(clknet_leaf_50_csclk),
    .D(net1176),
    .RESET_B(net435),
    .Q(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7084_ (.CLK(clknet_leaf_56_csclk),
    .D(net863),
    .RESET_B(net430),
    .Q(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__dfstp_4 _7085_ (.CLK(clknet_leaf_57_csclk),
    .D(_0674_),
    .SET_B(net428),
    .Q(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__dfstp_4 _7086_ (.CLK(clknet_leaf_58_csclk),
    .D(_0675_),
    .SET_B(net428),
    .Q(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7087_ (.CLK(clknet_leaf_60_csclk),
    .D(net518),
    .RESET_B(net428),
    .Q(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7088_ (.CLK(clknet_leaf_45_csclk),
    .D(_0677_),
    .RESET_B(net438),
    .Q(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7089_ (.CLK(clknet_leaf_43_csclk),
    .D(net713),
    .RESET_B(net437),
    .Q(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7090_ (.CLK(clknet_leaf_46_csclk),
    .D(net1130),
    .RESET_B(net438),
    .Q(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7091_ (.CLK(clknet_leaf_53_csclk),
    .D(net1110),
    .RESET_B(net432),
    .Q(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7092_ (.CLK(clknet_leaf_62_csclk),
    .D(net898),
    .RESET_B(net430),
    .Q(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__dfstp_4 _7093_ (.CLK(clknet_leaf_62_csclk),
    .D(_0682_),
    .SET_B(net430),
    .Q(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__dfstp_2 _7094_ (.CLK(clknet_leaf_60_csclk),
    .D(_0683_),
    .SET_B(net430),
    .Q(\gpio_configure[30][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7095_ (.CLK(clknet_leaf_43_csclk),
    .D(net589),
    .RESET_B(net437),
    .Q(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7096_ (.CLK(clknet_leaf_54_csclk),
    .D(_0685_),
    .RESET_B(net434),
    .Q(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7097_ (.CLK(clknet_leaf_43_csclk),
    .D(net732),
    .RESET_B(net437),
    .Q(\gpio_configure[30][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7098_ (.CLK(clknet_leaf_50_csclk),
    .D(net1097),
    .RESET_B(net435),
    .Q(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7099_ (.CLK(clknet_leaf_50_csclk),
    .D(net1171),
    .RESET_B(net435),
    .Q(\gpio_configure[30][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7100_ (.CLK(clknet_leaf_62_csclk),
    .D(net881),
    .RESET_B(net431),
    .Q(\gpio_configure[30][7] ));
 sky130_fd_sc_hd__dfstp_4 _7101_ (.CLK(clknet_leaf_62_csclk),
    .D(_0690_),
    .SET_B(net430),
    .Q(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__dfstp_2 _7102_ (.CLK(clknet_leaf_64_csclk),
    .D(net530),
    .SET_B(net436),
    .Q(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7103_ (.CLK(clknet_leaf_67_csclk),
    .D(net1322),
    .RESET_B(net436),
    .Q(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7104_ (.CLK(clknet_leaf_54_csclk),
    .D(_0693_),
    .RESET_B(net434),
    .Q(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7105_ (.CLK(clknet_leaf_68_csclk),
    .D(net1570),
    .RESET_B(net436),
    .Q(\gpio_configure[31][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7106_ (.CLK(clknet_leaf_48_csclk),
    .D(net582),
    .RESET_B(net438),
    .Q(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7107_ (.CLK(clknet_leaf_51_csclk),
    .D(net1102),
    .RESET_B(net435),
    .Q(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7108_ (.CLK(clknet_leaf_63_csclk),
    .D(net485),
    .RESET_B(net436),
    .Q(\gpio_configure[31][7] ));
 sky130_fd_sc_hd__dfstp_4 _7109_ (.CLK(clknet_leaf_30_csclk),
    .D(_0698_),
    .SET_B(net447),
    .Q(\gpio_configure[32][0] ));
 sky130_fd_sc_hd__dfstp_4 _7110_ (.CLK(clknet_leaf_18_csclk),
    .D(_0699_),
    .SET_B(net446),
    .Q(\gpio_configure[32][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7111_ (.CLK(clknet_leaf_27_csclk),
    .D(net1006),
    .RESET_B(net444),
    .Q(\gpio_configure[32][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7112_ (.CLK(clknet_leaf_34_csclk),
    .D(_0701_),
    .RESET_B(net454),
    .Q(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7113_ (.CLK(clknet_leaf_18_csclk),
    .D(net1282),
    .RESET_B(net446),
    .Q(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7114_ (.CLK(clknet_leaf_33_csclk),
    .D(net549),
    .RESET_B(net452),
    .Q(\gpio_configure[32][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7115_ (.CLK(clknet_leaf_33_csclk),
    .D(net1108),
    .RESET_B(net451),
    .Q(\gpio_configure[32][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7116_ (.CLK(clknet_leaf_31_csclk),
    .D(net477),
    .RESET_B(net447),
    .Q(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__dfstp_4 _7117_ (.CLK(clknet_leaf_30_csclk),
    .D(_0706_),
    .SET_B(net447),
    .Q(\gpio_configure[33][0] ));
 sky130_fd_sc_hd__dfstp_1 _7118_ (.CLK(clknet_leaf_64_csclk),
    .D(net499),
    .SET_B(net436),
    .Q(\gpio_configure[33][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7119_ (.CLK(clknet_opt_3_0_csclk),
    .D(net1288),
    .RESET_B(net437),
    .Q(\gpio_configure[33][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7120_ (.CLK(clknet_leaf_34_csclk),
    .D(net1027),
    .RESET_B(net454),
    .Q(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7121_ (.CLK(clknet_leaf_17_csclk),
    .D(net1296),
    .RESET_B(net442),
    .Q(\gpio_configure[33][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7122_ (.CLK(clknet_leaf_42_csclk),
    .D(net605),
    .RESET_B(net443),
    .Q(\gpio_configure[33][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7123_ (.CLK(clknet_leaf_55_csclk),
    .D(net1161),
    .RESET_B(net434),
    .Q(\gpio_configure[33][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7124_ (.CLK(clknet_leaf_44_csclk),
    .D(net943),
    .RESET_B(net437),
    .Q(\gpio_configure[33][7] ));
 sky130_fd_sc_hd__dfstp_4 _7125_ (.CLK(clknet_leaf_29_csclk),
    .D(_0714_),
    .SET_B(net448),
    .Q(\gpio_configure[34][0] ));
 sky130_fd_sc_hd__dfstp_4 _7126_ (.CLK(clknet_leaf_58_csclk),
    .D(_0715_),
    .SET_B(net428),
    .Q(\gpio_configure[34][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7127_ (.CLK(clknet_leaf_29_csclk),
    .D(net900),
    .RESET_B(net449),
    .Q(\gpio_configure[34][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7128_ (.CLK(clknet_leaf_34_csclk),
    .D(net1064),
    .RESET_B(net454),
    .Q(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7129_ (.CLK(clknet_leaf_58_csclk),
    .D(net681),
    .RESET_B(net429),
    .Q(\gpio_configure[34][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7130_ (.CLK(clknet_leaf_34_csclk),
    .D(net851),
    .RESET_B(net454),
    .Q(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7131_ (.CLK(clknet_leaf_53_csclk),
    .D(net1114),
    .RESET_B(net432),
    .Q(\gpio_configure[34][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7132_ (.CLK(clknet_leaf_57_csclk),
    .D(net902),
    .RESET_B(net432),
    .Q(\gpio_configure[34][7] ));
 sky130_fd_sc_hd__dfstp_1 _7133_ (.CLK(clknet_leaf_23_csclk),
    .D(_0722_),
    .SET_B(net443),
    .Q(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__dfstp_2 _7134_ (.CLK(clknet_leaf_59_csclk),
    .D(_0723_),
    .SET_B(net428),
    .Q(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7135_ (.CLK(clknet_leaf_60_csclk),
    .D(net525),
    .RESET_B(net430),
    .Q(\gpio_configure[35][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7136_ (.CLK(clknet_leaf_63_csclk),
    .D(net707),
    .RESET_B(net437),
    .Q(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7137_ (.CLK(clknet_3_6_0_csclk),
    .D(net1331),
    .RESET_B(net443),
    .Q(\gpio_configure[35][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7138_ (.CLK(clknet_leaf_47_csclk),
    .D(net1124),
    .RESET_B(net456),
    .Q(\gpio_configure[35][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7139_ (.CLK(clknet_leaf_50_csclk),
    .D(net1186),
    .RESET_B(net435),
    .Q(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7140_ (.CLK(clknet_leaf_56_csclk),
    .D(net890),
    .RESET_B(net428),
    .Q(\gpio_configure[35][7] ));
 sky130_fd_sc_hd__dfstp_4 _7141_ (.CLK(clknet_leaf_30_csclk),
    .D(_0730_),
    .SET_B(net448),
    .Q(\gpio_configure[36][0] ));
 sky130_fd_sc_hd__dfstp_4 _7142_ (.CLK(clknet_leaf_28_csclk),
    .D(_0731_),
    .SET_B(net446),
    .Q(\gpio_configure[36][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7143_ (.CLK(clknet_leaf_18_csclk),
    .D(net1594),
    .RESET_B(net449),
    .Q(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7144_ (.CLK(clknet_leaf_31_csclk),
    .D(net615),
    .RESET_B(net454),
    .Q(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7145_ (.CLK(clknet_leaf_18_csclk),
    .D(net1302),
    .RESET_B(net446),
    .Q(\gpio_configure[36][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7146_ (.CLK(clknet_leaf_33_csclk),
    .D(net914),
    .RESET_B(net452),
    .Q(\gpio_configure[36][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7147_ (.CLK(clknet_leaf_33_csclk),
    .D(net672),
    .RESET_B(net451),
    .Q(\gpio_configure[36][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7148_ (.CLK(clknet_leaf_32_csclk),
    .D(net812),
    .RESET_B(net447),
    .Q(\gpio_configure[36][7] ));
 sky130_fd_sc_hd__dfstp_4 _7149_ (.CLK(clknet_leaf_28_csclk),
    .D(_0738_),
    .SET_B(net445),
    .Q(\gpio_configure[37][0] ));
 sky130_fd_sc_hd__dfstp_2 _7150_ (.CLK(clknet_leaf_18_csclk),
    .D(_0739_),
    .SET_B(net444),
    .Q(\gpio_configure[37][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7151_ (.CLK(clknet_leaf_28_csclk),
    .D(net996),
    .RESET_B(net446),
    .Q(\gpio_configure[37][2] ));
 sky130_fd_sc_hd__dfrtp_2 _7152_ (.CLK(clknet_leaf_31_csclk),
    .D(net603),
    .RESET_B(net452),
    .Q(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7153_ (.CLK(clknet_leaf_19_csclk),
    .D(net1326),
    .RESET_B(net444),
    .Q(\gpio_configure[37][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7154_ (.CLK(clknet_leaf_33_csclk),
    .D(net927),
    .RESET_B(net451),
    .Q(\gpio_configure[37][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7155_ (.CLK(clknet_leaf_32_csclk),
    .D(net1066),
    .RESET_B(net452),
    .Q(\gpio_configure[37][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7156_ (.CLK(clknet_leaf_32_csclk),
    .D(net853),
    .RESET_B(net447),
    .Q(\gpio_configure[37][7] ));
 sky130_fd_sc_hd__dfrtp_2 _7157_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0746_),
    .RESET_B(net433),
    .Q(\xfer_count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7158_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0747_),
    .RESET_B(net433),
    .Q(\xfer_count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7159_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0748_),
    .RESET_B(net433),
    .Q(\xfer_count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7160_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0749_),
    .RESET_B(net433),
    .Q(\xfer_count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7161_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0750_),
    .RESET_B(net435),
    .Q(\pad_count_1[0] ));
 sky130_fd_sc_hd__dfstp_4 _7162_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0751_),
    .SET_B(net443),
    .Q(\pad_count_1[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7163_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0752_),
    .RESET_B(net455),
    .Q(\pad_count_1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7164_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0753_),
    .RESET_B(net455),
    .Q(\pad_count_1[3] ));
 sky130_fd_sc_hd__dfstp_4 _7165_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0754_),
    .SET_B(net455),
    .Q(\pad_count_1[4] ));
 sky130_fd_sc_hd__dfstp_4 _7166_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0755_),
    .SET_B(net455),
    .Q(\pad_count_2[0] ));
 sky130_fd_sc_hd__dfstp_4 _7167_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0756_),
    .SET_B(net455),
    .Q(\pad_count_2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7168_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0757_),
    .RESET_B(net455),
    .Q(\pad_count_2[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7169_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0758_),
    .RESET_B(net455),
    .Q(\pad_count_2[3] ));
 sky130_fd_sc_hd__dfstp_4 _7170_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0759_),
    .SET_B(net455),
    .Q(\pad_count_2[4] ));
 sky130_fd_sc_hd__dfrtp_2 _7171_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0760_),
    .RESET_B(net456),
    .Q(\pad_count_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7172_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(net460),
    .RESET_B(net433),
    .Q(serial_resetn_pre));
 sky130_fd_sc_hd__dfrtp_2 _7173_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0761_),
    .RESET_B(net433),
    .Q(serial_clock_pre));
 sky130_fd_sc_hd__dfrtp_1 _7174_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0762_),
    .RESET_B(net433),
    .Q(serial_load_pre));
 sky130_fd_sc_hd__dfrtp_2 _7175_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0763_),
    .RESET_B(net435),
    .Q(serial_busy));
 sky130_fd_sc_hd__dfrtp_4 _7176_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0764_),
    .RESET_B(net431),
    .Q(\serial_data_staging_1[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7177_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0765_),
    .RESET_B(net431),
    .Q(\serial_data_staging_1[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7178_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0766_),
    .RESET_B(net431),
    .Q(\serial_data_staging_1[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7179_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0767_),
    .RESET_B(net432),
    .Q(\serial_data_staging_1[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7180_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0768_),
    .RESET_B(net433),
    .Q(\serial_data_staging_1[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7181_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0769_),
    .RESET_B(net435),
    .Q(\serial_data_staging_1[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7182_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0770_),
    .RESET_B(net435),
    .Q(\serial_data_staging_1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _7183_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0771_),
    .RESET_B(net432),
    .Q(\serial_data_staging_1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7184_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0772_),
    .RESET_B(net420),
    .Q(\serial_data_staging_1[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7185_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0773_),
    .RESET_B(net415),
    .Q(\serial_data_staging_1[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7186_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0774_),
    .RESET_B(net420),
    .Q(\serial_data_staging_1[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7187_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0775_),
    .RESET_B(net419),
    .Q(\serial_data_staging_1[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7188_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0776_),
    .RESET_B(net419),
    .Q(\serial_data_staging_1[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7189_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0777_),
    .RESET_B(net431),
    .Q(\serial_data_staging_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7190_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0778_),
    .RESET_B(net429),
    .Q(\serial_data_staging_2[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7191_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0779_),
    .RESET_B(net432),
    .Q(\serial_data_staging_2[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7192_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0780_),
    .RESET_B(net432),
    .Q(\serial_data_staging_2[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7193_ (.CLK(clknet_3_3_0_wb_clk_i),
    .D(_0781_),
    .RESET_B(net435),
    .Q(\serial_data_staging_2[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7194_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0782_),
    .RESET_B(net435),
    .Q(\serial_data_staging_2[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7195_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0783_),
    .RESET_B(net435),
    .Q(\serial_data_staging_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7196_ (.CLK(clknet_3_2_0_wb_clk_i),
    .D(_0784_),
    .RESET_B(net435),
    .Q(\serial_data_staging_2[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7197_ (.CLK(clknet_3_1_0_wb_clk_i),
    .D(_0785_),
    .RESET_B(net421),
    .Q(\serial_data_staging_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7198_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0786_),
    .RESET_B(net415),
    .Q(\serial_data_staging_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7199_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0787_),
    .RESET_B(net415),
    .Q(\serial_data_staging_2[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7200_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0788_),
    .RESET_B(net414),
    .Q(\serial_data_staging_2[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7201_ (.CLK(clknet_3_0_0_wb_clk_i),
    .D(_0789_),
    .RESET_B(net419),
    .Q(\serial_data_staging_2[12] ));
 sky130_fd_sc_hd__dfrtp_2 _7202_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0790_),
    .RESET_B(net457),
    .Q(net317));
 sky130_fd_sc_hd__dfxtp_4 _7203_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0791_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_4 _7204_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0792_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_4 _7205_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0793_),
    .Q(net336));
 sky130_fd_sc_hd__dfxtp_4 _7206_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0794_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_4 _7207_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0795_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_4 _7208_ (.CLK(clknet_3_6_0_wb_clk_i),
    .D(_0796_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_4 _7209_ (.CLK(clknet_3_5_0_wb_clk_i),
    .D(_0797_),
    .Q(net341));
 sky130_fd_sc_hd__dfxtp_4 _7210_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0798_),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_2 _7211_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0799_),
    .RESET_B(net458),
    .Q(\wbbd_data[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7212_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0800_),
    .RESET_B(net458),
    .Q(\wbbd_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7213_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0801_),
    .RESET_B(net458),
    .Q(\wbbd_data[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7214_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0802_),
    .RESET_B(net458),
    .Q(\wbbd_data[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7215_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0803_),
    .RESET_B(net458),
    .Q(\wbbd_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7216_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0804_),
    .RESET_B(net458),
    .Q(\wbbd_data[5] ));
 sky130_fd_sc_hd__dfrtp_2 _7217_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0805_),
    .RESET_B(net458),
    .Q(\wbbd_data[6] ));
 sky130_fd_sc_hd__dfrtp_2 _7218_ (.CLK(clknet_3_7_0_wb_clk_i),
    .D(_0806_),
    .RESET_B(net458),
    .Q(\wbbd_data[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7219_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0807_),
    .RESET_B(net457),
    .Q(wbbd_sck));
 sky130_fd_sc_hd__dfrtp_4 _7220_ (.CLK(clknet_3_4_0_wb_clk_i),
    .D(_0808_),
    .RESET_B(net457),
    .Q(wbbd_write));
 sky130_fd_sc_hd__dfrtp_2 _7221_ (.CLK(clknet_leaf_73_csclk),
    .D(net1621),
    .RESET_B(net420),
    .Q(\gpio_configure[27][8] ));
 sky130_fd_sc_hd__dfrtp_2 _7222_ (.CLK(clknet_leaf_73_csclk),
    .D(net980),
    .RESET_B(net422),
    .Q(\gpio_configure[27][9] ));
 sky130_fd_sc_hd__dfstp_4 _7223_ (.CLK(clknet_leaf_74_csclk),
    .D(_0811_),
    .SET_B(net422),
    .Q(\gpio_configure[27][10] ));
 sky130_fd_sc_hd__dfrtp_2 _7224_ (.CLK(clknet_leaf_74_csclk),
    .D(net1440),
    .RESET_B(net420),
    .Q(\gpio_configure[27][11] ));
 sky130_fd_sc_hd__dfrtp_2 _7225_ (.CLK(clknet_leaf_74_csclk),
    .D(net1213),
    .RESET_B(net422),
    .Q(\gpio_configure[27][12] ));
 sky130_fd_sc_hd__inv_2 _3240__1 (.A(clknet_2_2_0_mgmt_gpio_in[4]),
    .Y(net461));
 sky130_fd_sc_hd__buf_2 _7227_ (.A(net87),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 _7228_ (.A(net65),
    .X(net315));
 sky130_fd_sc_hd__buf_2 _7229_ (.A(net66),
    .X(net316));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(wb_adr_i[18]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(wb_adr_i[17]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(wb_adr_i[16]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(wb_adr_i[15]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(wb_adr_i[14]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(wb_adr_i[13]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input102 (.A(wb_adr_i[12]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(wb_adr_i[11]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(wb_adr_i[10]),
    .X(net100));
 sky130_fd_sc_hd__buf_8 input99 (.A(wb_adr_i[0]),
    .X(net99));
 sky130_fd_sc_hd__buf_6 input98 (.A(usr2_vdd_pwrgood),
    .X(net98));
 sky130_fd_sc_hd__buf_6 input97 (.A(usr2_vcc_pwrgood),
    .X(net97));
 sky130_fd_sc_hd__buf_6 input96 (.A(usr1_vdd_pwrgood),
    .X(net96));
 sky130_fd_sc_hd__buf_6 input95 (.A(usr1_vcc_pwrgood),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(uart_enabled),
    .X(net94));
 sky130_fd_sc_hd__buf_8 input93 (.A(trap),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(spimemio_flash_io3_oeb),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(spimemio_flash_io3_do),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(spimemio_flash_io2_oeb),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(spimemio_flash_io2_do),
    .X(net89));
 sky130_fd_sc_hd__buf_8 input88 (.A(spimemio_flash_io1_oeb),
    .X(net88));
 sky130_fd_sc_hd__buf_8 input87 (.A(spimemio_flash_io1_do),
    .X(net87));
 sky130_fd_sc_hd__buf_8 input86 (.A(spimemio_flash_io0_oeb),
    .X(net86));
 sky130_fd_sc_hd__buf_6 input85 (.A(spimemio_flash_io0_do),
    .X(net85));
 sky130_fd_sc_hd__buf_6 input84 (.A(spimemio_flash_csb),
    .X(net84));
 sky130_fd_sc_hd__buf_6 input83 (.A(spimemio_flash_clk),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(spi_sdoenb),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(spi_sdo),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input80 (.A(spi_sck),
    .X(net80));
 sky130_fd_sc_hd__buf_6 input79 (.A(spi_enabled),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 input78 (.A(spi_csb),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(ser_tx),
    .X(net77));
 sky130_fd_sc_hd__buf_8 input76 (.A(qspi_enabled),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 input75 (.A(porb),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(pad_flash_io1_di),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(pad_flash_io0_di),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input72 (.A(mgmt_gpio_in[9]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(mgmt_gpio_in[8]),
    .X(net71));
 sky130_fd_sc_hd__buf_8 input70 (.A(mgmt_gpio_in[7]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(mgmt_gpio_in[6]),
    .X(net69));
 sky130_fd_sc_hd__buf_8 input68 (.A(mgmt_gpio_in[5]),
    .X(net68));
 sky130_fd_sc_hd__buf_8 input67 (.A(mgmt_gpio_in[3]),
    .X(net67));
 sky130_fd_sc_hd__buf_8 input66 (.A(mgmt_gpio_in[37]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input65 (.A(mgmt_gpio_in[36]),
    .X(net65));
 sky130_fd_sc_hd__buf_4 input64 (.A(mgmt_gpio_in[35]),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input63 (.A(mgmt_gpio_in[34]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input62 (.A(mgmt_gpio_in[33]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(mgmt_gpio_in[32]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input60 (.A(mgmt_gpio_in[31]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input59 (.A(mgmt_gpio_in[30]),
    .X(net59));
 sky130_fd_sc_hd__buf_8 input58 (.A(mgmt_gpio_in[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(mgmt_gpio_in[29]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input56 (.A(mgmt_gpio_in[28]),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input55 (.A(mgmt_gpio_in[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(mgmt_gpio_in[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(mgmt_gpio_in[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(mgmt_gpio_in[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(mgmt_gpio_in[23]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input50 (.A(mgmt_gpio_in[22]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input49 (.A(mgmt_gpio_in[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(mgmt_gpio_in[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(mgmt_gpio_in[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_6 input46 (.A(mgmt_gpio_in[19]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(mgmt_gpio_in[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(mgmt_gpio_in[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(mgmt_gpio_in[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(mgmt_gpio_in[15]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(mgmt_gpio_in[14]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(mgmt_gpio_in[13]),
    .X(net40));
 sky130_fd_sc_hd__buf_8 input39 (.A(mgmt_gpio_in[12]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input38 (.A(mgmt_gpio_in[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(mgmt_gpio_in[10]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input36 (.A(mgmt_gpio_in[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(mask_rev_in[9]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(mask_rev_in[8]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(mask_rev_in[7]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(mask_rev_in[6]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(mask_rev_in[5]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(mask_rev_in[4]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(mask_rev_in[3]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(mask_rev_in[31]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(mask_rev_in[30]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(mask_rev_in[2]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(mask_rev_in[29]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(mask_rev_in[28]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(mask_rev_in[27]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(mask_rev_in[26]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(mask_rev_in[25]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(mask_rev_in[24]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(mask_rev_in[23]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(mask_rev_in[22]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(mask_rev_in[21]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input16 (.A(mask_rev_in[20]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(mask_rev_in[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(mask_rev_in[19]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(mask_rev_in[18]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(mask_rev_in[17]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(mask_rev_in[16]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(mask_rev_in[15]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(mask_rev_in[14]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(mask_rev_in[13]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(mask_rev_in[12]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(mask_rev_in[11]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(mask_rev_in[10]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(mask_rev_in[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(debug_out),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(debug_oeb),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input1 (.A(debug_mode),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(wb_adr_i[19]),
    .X(net109));
 sky130_fd_sc_hd__buf_8 input110 (.A(wb_adr_i[1]),
    .X(net110));
 sky130_fd_sc_hd__buf_8 input111 (.A(wb_adr_i[20]),
    .X(net111));
 sky130_fd_sc_hd__buf_4 input112 (.A(wb_adr_i[21]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(wb_adr_i[22]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(wb_adr_i[23]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(wb_adr_i[24]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(wb_adr_i[25]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(wb_adr_i[26]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 input118 (.A(wb_adr_i[27]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(wb_adr_i[28]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(wb_adr_i[29]),
    .X(net120));
 sky130_fd_sc_hd__buf_8 input121 (.A(wb_adr_i[2]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(wb_adr_i[30]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(wb_adr_i[31]),
    .X(net123));
 sky130_fd_sc_hd__buf_8 input124 (.A(wb_adr_i[3]),
    .X(net124));
 sky130_fd_sc_hd__buf_8 input125 (.A(wb_adr_i[4]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 input126 (.A(wb_adr_i[5]),
    .X(net126));
 sky130_fd_sc_hd__buf_8 input127 (.A(wb_adr_i[6]),
    .X(net127));
 sky130_fd_sc_hd__buf_8 input128 (.A(wb_adr_i[7]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 input129 (.A(wb_adr_i[8]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 input130 (.A(wb_adr_i[9]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(wb_cyc_i),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 input132 (.A(wb_dat_i[0]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(wb_dat_i[10]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(wb_dat_i[11]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(wb_dat_i[12]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(wb_dat_i[13]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(wb_dat_i[14]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(wb_dat_i[15]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 input139 (.A(wb_dat_i[16]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input140 (.A(wb_dat_i[17]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(wb_dat_i[18]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 input142 (.A(wb_dat_i[19]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 input143 (.A(wb_dat_i[1]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(wb_dat_i[20]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 input145 (.A(wb_dat_i[21]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 input146 (.A(wb_dat_i[22]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(wb_dat_i[23]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(wb_dat_i[24]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 input149 (.A(wb_dat_i[25]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input150 (.A(wb_dat_i[26]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 input151 (.A(wb_dat_i[27]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(wb_dat_i[28]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(wb_dat_i[29]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(wb_dat_i[2]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(wb_dat_i[30]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(wb_dat_i[31]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(wb_dat_i[3]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(wb_dat_i[4]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(wb_dat_i[5]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(wb_dat_i[6]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(wb_dat_i[7]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(wb_dat_i[8]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(wb_dat_i[9]),
    .X(net163));
 sky130_fd_sc_hd__buf_6 input164 (.A(wb_rstn_i),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 input165 (.A(wb_sel_i[0]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 input166 (.A(wb_sel_i[1]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 input167 (.A(wb_sel_i[2]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 input168 (.A(wb_sel_i[3]),
    .X(net168));
 sky130_fd_sc_hd__buf_6 input169 (.A(wb_stb_i),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input170 (.A(wb_we_i),
    .X(net170));
 sky130_fd_sc_hd__buf_8 output171 (.A(net171),
    .X(debug_in));
 sky130_fd_sc_hd__buf_8 output172 (.A(net172),
    .X(irq[0]));
 sky130_fd_sc_hd__buf_8 output173 (.A(net173),
    .X(irq[1]));
 sky130_fd_sc_hd__buf_8 output174 (.A(net174),
    .X(irq[2]));
 sky130_fd_sc_hd__buf_8 output175 (.A(net175),
    .X(mgmt_gpio_oeb[0]));
 sky130_fd_sc_hd__buf_8 output176 (.A(net176),
    .X(mgmt_gpio_oeb[10]));
 sky130_fd_sc_hd__buf_8 output177 (.A(net177),
    .X(mgmt_gpio_oeb[11]));
 sky130_fd_sc_hd__buf_8 output178 (.A(net178),
    .X(mgmt_gpio_oeb[12]));
 sky130_fd_sc_hd__buf_8 output179 (.A(net179),
    .X(mgmt_gpio_oeb[13]));
 sky130_fd_sc_hd__buf_8 output180 (.A(net180),
    .X(mgmt_gpio_oeb[14]));
 sky130_fd_sc_hd__buf_8 output181 (.A(net181),
    .X(mgmt_gpio_oeb[15]));
 sky130_fd_sc_hd__buf_8 output182 (.A(net182),
    .X(mgmt_gpio_oeb[16]));
 sky130_fd_sc_hd__buf_8 output183 (.A(net183),
    .X(mgmt_gpio_oeb[17]));
 sky130_fd_sc_hd__buf_8 output184 (.A(net184),
    .X(mgmt_gpio_oeb[18]));
 sky130_fd_sc_hd__buf_8 output185 (.A(net185),
    .X(mgmt_gpio_oeb[19]));
 sky130_fd_sc_hd__buf_8 output186 (.A(net186),
    .X(mgmt_gpio_oeb[1]));
 sky130_fd_sc_hd__buf_8 output187 (.A(net187),
    .X(mgmt_gpio_oeb[20]));
 sky130_fd_sc_hd__buf_8 output188 (.A(net188),
    .X(mgmt_gpio_oeb[21]));
 sky130_fd_sc_hd__buf_8 output189 (.A(net189),
    .X(mgmt_gpio_oeb[22]));
 sky130_fd_sc_hd__buf_8 output190 (.A(net190),
    .X(mgmt_gpio_oeb[23]));
 sky130_fd_sc_hd__buf_8 output191 (.A(net191),
    .X(mgmt_gpio_oeb[24]));
 sky130_fd_sc_hd__buf_8 output192 (.A(net192),
    .X(mgmt_gpio_oeb[25]));
 sky130_fd_sc_hd__buf_8 output193 (.A(net193),
    .X(mgmt_gpio_oeb[26]));
 sky130_fd_sc_hd__buf_8 output194 (.A(net194),
    .X(mgmt_gpio_oeb[27]));
 sky130_fd_sc_hd__buf_8 output195 (.A(net195),
    .X(mgmt_gpio_oeb[28]));
 sky130_fd_sc_hd__buf_8 output196 (.A(net196),
    .X(mgmt_gpio_oeb[29]));
 sky130_fd_sc_hd__buf_8 output197 (.A(net197),
    .X(mgmt_gpio_oeb[2]));
 sky130_fd_sc_hd__buf_8 output198 (.A(net198),
    .X(mgmt_gpio_oeb[30]));
 sky130_fd_sc_hd__buf_8 output199 (.A(net199),
    .X(mgmt_gpio_oeb[31]));
 sky130_fd_sc_hd__buf_8 output200 (.A(net200),
    .X(mgmt_gpio_oeb[32]));
 sky130_fd_sc_hd__buf_8 output201 (.A(net201),
    .X(mgmt_gpio_oeb[33]));
 sky130_fd_sc_hd__buf_8 output202 (.A(net202),
    .X(mgmt_gpio_oeb[34]));
 sky130_fd_sc_hd__buf_8 output203 (.A(net203),
    .X(mgmt_gpio_oeb[35]));
 sky130_fd_sc_hd__buf_8 output204 (.A(net204),
    .X(mgmt_gpio_oeb[36]));
 sky130_fd_sc_hd__buf_8 output205 (.A(net205),
    .X(mgmt_gpio_oeb[37]));
 sky130_fd_sc_hd__buf_8 output206 (.A(net206),
    .X(mgmt_gpio_oeb[3]));
 sky130_fd_sc_hd__buf_8 output207 (.A(net207),
    .X(mgmt_gpio_oeb[4]));
 sky130_fd_sc_hd__buf_8 output208 (.A(net208),
    .X(mgmt_gpio_oeb[5]));
 sky130_fd_sc_hd__buf_8 output209 (.A(net209),
    .X(mgmt_gpio_oeb[6]));
 sky130_fd_sc_hd__buf_8 output210 (.A(net210),
    .X(mgmt_gpio_oeb[7]));
 sky130_fd_sc_hd__buf_8 output211 (.A(net211),
    .X(mgmt_gpio_oeb[8]));
 sky130_fd_sc_hd__buf_8 output212 (.A(net212),
    .X(mgmt_gpio_oeb[9]));
 sky130_fd_sc_hd__buf_8 output213 (.A(net213),
    .X(mgmt_gpio_out[0]));
 sky130_fd_sc_hd__buf_8 output214 (.A(net214),
    .X(mgmt_gpio_out[10]));
 sky130_fd_sc_hd__buf_8 output215 (.A(net215),
    .X(mgmt_gpio_out[11]));
 sky130_fd_sc_hd__buf_8 output216 (.A(net216),
    .X(mgmt_gpio_out[12]));
 sky130_fd_sc_hd__buf_8 output217 (.A(net217),
    .X(mgmt_gpio_out[13]));
 sky130_fd_sc_hd__clkbuf_4 output218 (.A(net218),
    .X(mgmt_gpio_out[14]));
 sky130_fd_sc_hd__clkbuf_4 output219 (.A(net219),
    .X(mgmt_gpio_out[15]));
 sky130_fd_sc_hd__buf_8 output220 (.A(net220),
    .X(mgmt_gpio_out[16]));
 sky130_fd_sc_hd__buf_8 output221 (.A(net221),
    .X(mgmt_gpio_out[17]));
 sky130_fd_sc_hd__buf_8 output222 (.A(net222),
    .X(mgmt_gpio_out[18]));
 sky130_fd_sc_hd__buf_8 output223 (.A(net223),
    .X(mgmt_gpio_out[19]));
 sky130_fd_sc_hd__buf_8 output224 (.A(net224),
    .X(mgmt_gpio_out[1]));
 sky130_fd_sc_hd__buf_8 output225 (.A(net225),
    .X(mgmt_gpio_out[20]));
 sky130_fd_sc_hd__buf_8 output226 (.A(net226),
    .X(mgmt_gpio_out[21]));
 sky130_fd_sc_hd__buf_8 output227 (.A(net227),
    .X(mgmt_gpio_out[22]));
 sky130_fd_sc_hd__buf_8 output228 (.A(net228),
    .X(mgmt_gpio_out[23]));
 sky130_fd_sc_hd__buf_8 output229 (.A(net229),
    .X(mgmt_gpio_out[24]));
 sky130_fd_sc_hd__buf_8 output230 (.A(net230),
    .X(mgmt_gpio_out[25]));
 sky130_fd_sc_hd__buf_8 output231 (.A(net231),
    .X(mgmt_gpio_out[26]));
 sky130_fd_sc_hd__buf_8 output232 (.A(net232),
    .X(mgmt_gpio_out[27]));
 sky130_fd_sc_hd__buf_8 output233 (.A(net233),
    .X(mgmt_gpio_out[28]));
 sky130_fd_sc_hd__buf_8 output234 (.A(net234),
    .X(mgmt_gpio_out[29]));
 sky130_fd_sc_hd__buf_8 output235 (.A(net235),
    .X(mgmt_gpio_out[2]));
 sky130_fd_sc_hd__buf_8 output236 (.A(net236),
    .X(mgmt_gpio_out[30]));
 sky130_fd_sc_hd__buf_8 output237 (.A(net237),
    .X(mgmt_gpio_out[31]));
 sky130_fd_sc_hd__buf_8 output238 (.A(net238),
    .X(mgmt_gpio_out[32]));
 sky130_fd_sc_hd__buf_8 output239 (.A(net239),
    .X(mgmt_gpio_out[33]));
 sky130_fd_sc_hd__buf_8 output240 (.A(net240),
    .X(mgmt_gpio_out[34]));
 sky130_fd_sc_hd__buf_8 output241 (.A(net241),
    .X(mgmt_gpio_out[35]));
 sky130_fd_sc_hd__buf_8 output242 (.A(net242),
    .X(mgmt_gpio_out[36]));
 sky130_fd_sc_hd__buf_8 output243 (.A(net243),
    .X(mgmt_gpio_out[37]));
 sky130_fd_sc_hd__buf_8 output244 (.A(net244),
    .X(mgmt_gpio_out[3]));
 sky130_fd_sc_hd__buf_8 output245 (.A(net245),
    .X(mgmt_gpio_out[4]));
 sky130_fd_sc_hd__buf_8 output246 (.A(net246),
    .X(mgmt_gpio_out[5]));
 sky130_fd_sc_hd__buf_8 output247 (.A(net247),
    .X(mgmt_gpio_out[6]));
 sky130_fd_sc_hd__buf_8 output248 (.A(net248),
    .X(mgmt_gpio_out[7]));
 sky130_fd_sc_hd__buf_8 output249 (.A(net249),
    .X(mgmt_gpio_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net250),
    .X(mgmt_gpio_out[9]));
 sky130_fd_sc_hd__clkbuf_4 output251 (.A(net251),
    .X(pad_flash_clk));
 sky130_fd_sc_hd__buf_8 output252 (.A(net252),
    .X(pad_flash_clk_oeb));
 sky130_fd_sc_hd__buf_8 output253 (.A(net253),
    .X(pad_flash_csb));
 sky130_fd_sc_hd__buf_8 output254 (.A(net254),
    .X(pad_flash_csb_oeb));
 sky130_fd_sc_hd__buf_8 output255 (.A(net255),
    .X(pad_flash_io0_do));
 sky130_fd_sc_hd__buf_8 output256 (.A(net256),
    .X(pad_flash_io0_ieb));
 sky130_fd_sc_hd__buf_8 output257 (.A(net257),
    .X(pad_flash_io0_oeb));
 sky130_fd_sc_hd__buf_8 output258 (.A(net258),
    .X(pad_flash_io1_do));
 sky130_fd_sc_hd__buf_8 output259 (.A(net259),
    .X(pad_flash_io1_ieb));
 sky130_fd_sc_hd__buf_8 output260 (.A(net260),
    .X(pad_flash_io1_oeb));
 sky130_fd_sc_hd__buf_8 output261 (.A(net261),
    .X(pll90_sel[0]));
 sky130_fd_sc_hd__buf_8 output262 (.A(net262),
    .X(pll90_sel[1]));
 sky130_fd_sc_hd__buf_8 output263 (.A(net263),
    .X(pll90_sel[2]));
 sky130_fd_sc_hd__buf_8 output264 (.A(net264),
    .X(pll_bypass));
 sky130_fd_sc_hd__buf_8 output265 (.A(net265),
    .X(pll_dco_ena));
 sky130_fd_sc_hd__buf_8 output266 (.A(net266),
    .X(pll_div[0]));
 sky130_fd_sc_hd__buf_8 output267 (.A(net267),
    .X(pll_div[1]));
 sky130_fd_sc_hd__buf_8 output268 (.A(net268),
    .X(pll_div[2]));
 sky130_fd_sc_hd__buf_8 output269 (.A(net269),
    .X(pll_div[3]));
 sky130_fd_sc_hd__buf_8 output270 (.A(net270),
    .X(pll_div[4]));
 sky130_fd_sc_hd__buf_8 output271 (.A(net271),
    .X(pll_ena));
 sky130_fd_sc_hd__buf_8 output272 (.A(net272),
    .X(pll_sel[0]));
 sky130_fd_sc_hd__buf_8 output273 (.A(net273),
    .X(pll_sel[1]));
 sky130_fd_sc_hd__buf_8 output274 (.A(net274),
    .X(pll_sel[2]));
 sky130_fd_sc_hd__buf_8 output275 (.A(net275),
    .X(pll_trim[0]));
 sky130_fd_sc_hd__buf_8 output276 (.A(net276),
    .X(pll_trim[10]));
 sky130_fd_sc_hd__buf_8 output277 (.A(net277),
    .X(pll_trim[11]));
 sky130_fd_sc_hd__buf_8 output278 (.A(net278),
    .X(pll_trim[12]));
 sky130_fd_sc_hd__buf_8 output279 (.A(net279),
    .X(pll_trim[13]));
 sky130_fd_sc_hd__buf_8 output280 (.A(net280),
    .X(pll_trim[14]));
 sky130_fd_sc_hd__buf_8 output281 (.A(net281),
    .X(pll_trim[15]));
 sky130_fd_sc_hd__buf_8 output282 (.A(net282),
    .X(pll_trim[16]));
 sky130_fd_sc_hd__buf_8 output283 (.A(net283),
    .X(pll_trim[17]));
 sky130_fd_sc_hd__buf_8 output284 (.A(net284),
    .X(pll_trim[18]));
 sky130_fd_sc_hd__buf_8 output285 (.A(net285),
    .X(pll_trim[19]));
 sky130_fd_sc_hd__buf_8 output286 (.A(net286),
    .X(pll_trim[1]));
 sky130_fd_sc_hd__buf_8 output287 (.A(net287),
    .X(pll_trim[20]));
 sky130_fd_sc_hd__buf_8 output288 (.A(net288),
    .X(pll_trim[21]));
 sky130_fd_sc_hd__buf_8 output289 (.A(net289),
    .X(pll_trim[22]));
 sky130_fd_sc_hd__buf_8 output290 (.A(net290),
    .X(pll_trim[23]));
 sky130_fd_sc_hd__buf_8 output291 (.A(net291),
    .X(pll_trim[24]));
 sky130_fd_sc_hd__buf_8 output292 (.A(net292),
    .X(pll_trim[25]));
 sky130_fd_sc_hd__buf_8 output293 (.A(net293),
    .X(pll_trim[2]));
 sky130_fd_sc_hd__buf_8 output294 (.A(net294),
    .X(pll_trim[3]));
 sky130_fd_sc_hd__buf_8 output295 (.A(net295),
    .X(pll_trim[4]));
 sky130_fd_sc_hd__buf_8 output296 (.A(net296),
    .X(pll_trim[5]));
 sky130_fd_sc_hd__buf_8 output297 (.A(net297),
    .X(pll_trim[6]));
 sky130_fd_sc_hd__buf_8 output298 (.A(net298),
    .X(pll_trim[7]));
 sky130_fd_sc_hd__buf_8 output299 (.A(net299),
    .X(pll_trim[8]));
 sky130_fd_sc_hd__buf_8 output300 (.A(net300),
    .X(pll_trim[9]));
 sky130_fd_sc_hd__buf_8 output301 (.A(net301),
    .X(pwr_ctrl_out[0]));
 sky130_fd_sc_hd__buf_8 output302 (.A(net302),
    .X(pwr_ctrl_out[1]));
 sky130_fd_sc_hd__buf_8 output303 (.A(net303),
    .X(pwr_ctrl_out[2]));
 sky130_fd_sc_hd__buf_8 output304 (.A(net304),
    .X(pwr_ctrl_out[3]));
 sky130_fd_sc_hd__buf_8 output305 (.A(net305),
    .X(reset));
 sky130_fd_sc_hd__buf_8 output306 (.A(net306),
    .X(ser_rx));
 sky130_fd_sc_hd__buf_8 output307 (.A(net307),
    .X(serial_clock));
 sky130_fd_sc_hd__buf_8 output308 (.A(net308),
    .X(serial_data_1));
 sky130_fd_sc_hd__buf_8 output309 (.A(net309),
    .X(serial_data_2));
 sky130_fd_sc_hd__buf_8 output310 (.A(net310),
    .X(serial_load));
 sky130_fd_sc_hd__buf_8 output311 (.A(net311),
    .X(serial_resetn));
 sky130_fd_sc_hd__buf_8 output312 (.A(net312),
    .X(spi_sdi));
 sky130_fd_sc_hd__buf_8 output313 (.A(net313),
    .X(spimemio_flash_io0_di));
 sky130_fd_sc_hd__buf_8 output314 (.A(net314),
    .X(spimemio_flash_io1_di));
 sky130_fd_sc_hd__buf_8 output315 (.A(net315),
    .X(spimemio_flash_io2_di));
 sky130_fd_sc_hd__buf_8 output316 (.A(net316),
    .X(spimemio_flash_io3_di));
 sky130_fd_sc_hd__buf_8 output317 (.A(net317),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_8 output318 (.A(net318),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_8 output319 (.A(net319),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_8 output320 (.A(net320),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_8 output321 (.A(net321),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_8 output322 (.A(net322),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_8 output323 (.A(net323),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_8 output324 (.A(net324),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_8 output325 (.A(net325),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_8 output326 (.A(net326),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_8 output327 (.A(net327),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_8 output328 (.A(net328),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_8 output329 (.A(net329),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_8 output330 (.A(net330),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_8 output331 (.A(net331),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_8 output332 (.A(net332),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_8 output333 (.A(net333),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_8 output334 (.A(net334),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_8 output335 (.A(net335),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_8 output336 (.A(net336),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_8 output337 (.A(net337),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_8 output338 (.A(net338),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_8 output339 (.A(net339),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_8 output340 (.A(net340),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_8 output341 (.A(net341),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_8 output342 (.A(net342),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_8 output343 (.A(net343),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_8 output344 (.A(net344),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_8 output345 (.A(net345),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_8 output346 (.A(net346),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__buf_8 output347 (.A(net347),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_8 output348 (.A(net348),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_8 output349 (.A(net349),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_6 max_cap350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_6 wire351 (.A(_2841_),
    .X(net351));
 sky130_fd_sc_hd__buf_8 fanout352 (.A(_2493_),
    .X(net352));
 sky130_fd_sc_hd__buf_8 fanout353 (.A(_2492_),
    .X(net353));
 sky130_fd_sc_hd__buf_8 load_slew354 (.A(_0893_),
    .X(net354));
 sky130_fd_sc_hd__buf_8 load_slew355 (.A(_0883_),
    .X(net355));
 sky130_fd_sc_hd__buf_8 load_slew356 (.A(_0868_),
    .X(net356));
 sky130_fd_sc_hd__buf_8 load_slew357 (.A(net515),
    .X(net357));
 sky130_fd_sc_hd__buf_8 load_slew358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_8 max_cap359 (.A(net522),
    .X(net359));
 sky130_fd_sc_hd__buf_8 max_cap360 (.A(net609),
    .X(net360));
 sky130_fd_sc_hd__buf_8 fanout361 (.A(_1805_),
    .X(net361));
 sky130_fd_sc_hd__buf_8 fanout362 (.A(net509),
    .X(net362));
 sky130_fd_sc_hd__buf_8 fanout363 (.A(net509),
    .X(net363));
 sky130_fd_sc_hd__buf_8 fanout364 (.A(net562),
    .X(net364));
 sky130_fd_sc_hd__buf_8 fanout365 (.A(net562),
    .X(net365));
 sky130_fd_sc_hd__bufbuf_16 fanout366 (.A(net562),
    .X(net366));
 sky130_fd_sc_hd__buf_8 fanout367 (.A(_1866_),
    .X(net367));
 sky130_fd_sc_hd__buf_8 fanout368 (.A(_1709_),
    .X(net368));
 sky130_fd_sc_hd__buf_8 fanout369 (.A(net465),
    .X(net369));
 sky130_fd_sc_hd__buf_8 fanout370 (.A(net476),
    .X(net370));
 sky130_fd_sc_hd__buf_8 fanout371 (.A(net474),
    .X(net371));
 sky130_fd_sc_hd__buf_8 fanout372 (.A(net592),
    .X(net372));
 sky130_fd_sc_hd__buf_8 fanout373 (.A(net592),
    .X(net373));
 sky130_fd_sc_hd__buf_8 fanout374 (.A(net669),
    .X(net374));
 sky130_fd_sc_hd__buf_8 fanout375 (.A(net469),
    .X(net375));
 sky130_fd_sc_hd__buf_8 fanout376 (.A(net540),
    .X(net376));
 sky130_fd_sc_hd__buf_8 fanout377 (.A(net538),
    .X(net377));
 sky130_fd_sc_hd__buf_8 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_8 fanout379 (.A(net631),
    .X(net379));
 sky130_fd_sc_hd__buf_8 fanout380 (.A(net645),
    .X(net380));
 sky130_fd_sc_hd__buf_8 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_8 fanout382 (.A(net645),
    .X(net382));
 sky130_fd_sc_hd__buf_8 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_8 fanout384 (.A(net598),
    .X(net384));
 sky130_fd_sc_hd__buf_8 fanout385 (.A(net597),
    .X(net385));
 sky130_fd_sc_hd__buf_8 fanout386 (.A(net533),
    .X(net386));
 sky130_fd_sc_hd__buf_8 fanout387 (.A(net597),
    .X(net387));
 sky130_fd_sc_hd__buf_8 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_8 fanout389 (.A(net495),
    .X(net389));
 sky130_fd_sc_hd__buf_8 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_8 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net495),
    .X(net392));
 sky130_fd_sc_hd__buf_8 fanout393 (.A(net503),
    .X(net393));
 sky130_fd_sc_hd__buf_8 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_8 fanout395 (.A(net529),
    .X(net395));
 sky130_fd_sc_hd__buf_8 fanout396 (.A(net529),
    .X(net396));
 sky130_fd_sc_hd__buf_8 fanout397 (.A(net529),
    .X(net397));
 sky130_fd_sc_hd__buf_8 fanout398 (.A(net529),
    .X(net398));
 sky130_fd_sc_hd__buf_8 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_8 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__buf_8 fanout401 (.A(net1347),
    .X(net401));
 sky130_fd_sc_hd__buf_8 fanout402 (.A(net1347),
    .X(net402));
 sky130_fd_sc_hd__buf_8 fanout403 (.A(net1347),
    .X(net403));
 sky130_fd_sc_hd__buf_8 fanout404 (.A(_0830_),
    .X(net404));
 sky130_fd_sc_hd__buf_8 fanout405 (.A(_0819_),
    .X(net405));
 sky130_fd_sc_hd__buf_8 fanout406 (.A(net675),
    .X(net406));
 sky130_fd_sc_hd__buf_8 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_8 fanout408 (.A(\xfer_state[1] ),
    .X(net408));
 sky130_fd_sc_hd__buf_8 fanout409 (.A(\hkspi.state[3] ),
    .X(net409));
 sky130_fd_sc_hd__buf_8 fanout410 (.A(net412),
    .X(net410));
 sky130_fd_sc_hd__buf_8 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_8 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_8 fanout413 (.A(_1426_),
    .X(net413));
 sky130_fd_sc_hd__buf_8 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__buf_8 fanout415 (.A(net423),
    .X(net415));
 sky130_fd_sc_hd__buf_8 fanout416 (.A(net423),
    .X(net416));
 sky130_fd_sc_hd__buf_8 fanout417 (.A(net423),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(net423),
    .X(net418));
 sky130_fd_sc_hd__buf_8 fanout419 (.A(net421),
    .X(net419));
 sky130_fd_sc_hd__buf_8 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_8 fanout421 (.A(net423),
    .X(net421));
 sky130_fd_sc_hd__buf_8 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_8 fanout423 (.A(net456),
    .X(net423));
 sky130_fd_sc_hd__buf_8 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_8 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_8 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_8 fanout427 (.A(net456),
    .X(net427));
 sky130_fd_sc_hd__buf_8 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_8 fanout429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__buf_8 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_8 fanout431 (.A(net456),
    .X(net431));
 sky130_fd_sc_hd__buf_8 fanout432 (.A(net435),
    .X(net432));
 sky130_fd_sc_hd__buf_8 fanout433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_8 fanout435 (.A(net456),
    .X(net435));
 sky130_fd_sc_hd__buf_8 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_8 fanout437 (.A(net456),
    .X(net437));
 sky130_fd_sc_hd__buf_8 fanout438 (.A(net456),
    .X(net438));
 sky130_fd_sc_hd__buf_8 fanout439 (.A(net456),
    .X(net439));
 sky130_fd_sc_hd__buf_8 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__buf_8 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_8 fanout442 (.A(net456),
    .X(net442));
 sky130_fd_sc_hd__buf_8 fanout443 (.A(net455),
    .X(net443));
 sky130_fd_sc_hd__buf_8 fanout444 (.A(net455),
    .X(net444));
 sky130_fd_sc_hd__buf_8 fanout445 (.A(net455),
    .X(net445));
 sky130_fd_sc_hd__buf_8 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__buf_8 fanout447 (.A(net449),
    .X(net447));
 sky130_fd_sc_hd__buf_8 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_8 fanout449 (.A(net455),
    .X(net449));
 sky130_fd_sc_hd__buf_8 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_8 fanout451 (.A(net455),
    .X(net451));
 sky130_fd_sc_hd__buf_8 fanout452 (.A(net454),
    .X(net452));
 sky130_fd_sc_hd__buf_8 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_8 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_8 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_8 fanout456 (.A(net75),
    .X(net456));
 sky130_fd_sc_hd__buf_8 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_8 fanout458 (.A(net164),
    .X(net458));
 sky130_fd_sc_hd__buf_8 fanout459 (.A(net126),
    .X(net459));
 sky130_fd_sc_hd__conb_1 _7172__460 (.HI(net460));
 sky130_fd_sc_hd__inv_2 net399_2 (.A(clknet_2_2_0_mgmt_gpio_in[4]),
    .Y(net462));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_0_mgmt_gpio_in[4]  (.A(mgmt_gpio_in[4]),
    .X(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_0_0_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_1_0_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_1_1_0_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_1_1_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_0_0_mgmt_gpio_in[4]  (.A(clknet_1_0_0_mgmt_gpio_in[4]),
    .X(clknet_2_0_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_1_0_mgmt_gpio_in[4]  (.A(clknet_1_0_0_mgmt_gpio_in[4]),
    .X(clknet_2_1_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_2_0_mgmt_gpio_in[4]  (.A(clknet_1_1_0_mgmt_gpio_in[4]),
    .X(clknet_2_2_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 \clkbuf_2_3_0_mgmt_gpio_in[4]  (.A(clknet_1_1_0_mgmt_gpio_in[4]),
    .X(clknet_2_3_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_2_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_3_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_4_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_5_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_7_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_8_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_10_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_11_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_csclk (.A(clknet_opt_4_0_csclk),
    .X(clknet_leaf_12_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_13_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_14_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_15_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_16_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_17_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_18_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_19_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_20_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_21_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_22_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_23_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_24_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_25_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_26_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_27_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_28_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_29_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_30_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_31_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_32_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_33_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_34_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_35_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_36_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_37_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_38_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_39_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_40_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_42_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_43_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_44_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_45_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_46_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_47_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_48_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_49_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_50_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_51_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_52_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_53_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_54_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_55_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_56_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_57_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_58_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_59_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_60_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_61_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_62_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_63_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_64_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_65_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_67_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_68_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_69_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_70_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_csclk (.A(clknet_opt_1_0_csclk),
    .X(clknet_leaf_71_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_72_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_73_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_74_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_75_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_76_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_csclk (.A(clknet_opt_2_0_csclk),
    .X(clknet_leaf_77_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_78_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_csclk (.A(csclk),
    .X(clknet_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_csclk (.A(clknet_1_0_0_csclk),
    .X(clknet_1_0_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_csclk (.A(clknet_0_csclk),
    .X(clknet_1_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_csclk (.A(clknet_1_1_0_csclk),
    .X(clknet_1_1_1_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_csclk (.A(clknet_1_0_1_csclk),
    .X(clknet_2_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_csclk (.A(clknet_1_1_1_csclk),
    .X(clknet_2_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_csclk (.A(clknet_2_0_0_csclk),
    .X(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_csclk (.A(clknet_2_1_0_csclk),
    .X(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_csclk (.A(clknet_2_2_0_csclk),
    .X(clknet_3_5_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_csclk (.A(clknet_2_3_0_csclk),
    .X(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_opt_1_0_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_opt_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_opt_2_0_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_opt_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_opt_3_0_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_opt_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_opt_4_0_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_opt_4_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0__1132_ (.A(_1132_),
    .X(clknet_0__1132_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f__1132_ (.A(clknet_0__1132_),
    .X(clknet_1_0__leaf__1132_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f__1132_ (.A(clknet_0__1132_),
    .X(clknet_1_1__leaf__1132_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_wbbd_sck (.A(wbbd_sck),
    .X(clknet_0_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_0__leaf_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_1__leaf_wbbd_sck));
 sky130_fd_sc_hd__bufbuf_16 hold1 (.A(net471),
    .X(net463));
 sky130_fd_sc_hd__bufbuf_16 hold2 (.A(net473),
    .X(net464));
 sky130_fd_sc_hd__bufbuf_16 hold3 (.A(net475),
    .X(net465));
 sky130_fd_sc_hd__bufbuf_16 hold4 (.A(_0296_),
    .X(net466));
 sky130_fd_sc_hd__bufbuf_16 hold5 (.A(net535),
    .X(net467));
 sky130_fd_sc_hd__bufbuf_16 hold6 (.A(net537),
    .X(net468));
 sky130_fd_sc_hd__bufbuf_16 hold7 (.A(net539),
    .X(net469));
 sky130_fd_sc_hd__bufbuf_16 hold8 (.A(_0294_),
    .X(net470));
 sky130_fd_sc_hd__bufbuf_16 hold9 (.A(\hkspi.odata[7] ),
    .X(net471));
 sky130_fd_sc_hd__bufbuf_16 hold10 (.A(net463),
    .X(net472));
 sky130_fd_sc_hd__bufbuf_16 hold11 (.A(_1474_),
    .X(net473));
 sky130_fd_sc_hd__bufbuf_16 hold12 (.A(net464),
    .X(net474));
 sky130_fd_sc_hd__bufbuf_16 hold13 (.A(net371),
    .X(net475));
 sky130_fd_sc_hd__bufbuf_16 hold14 (.A(net465),
    .X(net476));
 sky130_fd_sc_hd__bufbuf_16 hold15 (.A(_0705_),
    .X(net477));
 sky130_fd_sc_hd__bufbuf_16 hold16 (.A(\hkspi.addr[1] ),
    .X(net478));
 sky130_fd_sc_hd__bufbuf_16 hold17 (.A(_0857_),
    .X(net479));
 sky130_fd_sc_hd__bufbuf_16 hold18 (.A(net788),
    .X(net480));
 sky130_fd_sc_hd__bufbuf_16 hold19 (.A(_0861_),
    .X(net481));
 sky130_fd_sc_hd__bufbuf_16 hold20 (.A(_0896_),
    .X(net482));
 sky130_fd_sc_hd__bufbuf_16 hold21 (.A(_0944_),
    .X(net483));
 sky130_fd_sc_hd__bufbuf_16 hold22 (.A(_2442_),
    .X(net484));
 sky130_fd_sc_hd__bufbuf_16 hold23 (.A(_0697_),
    .X(net485));
 sky130_fd_sc_hd__bufbuf_16 hold24 (.A(\hkspi.addr[2] ),
    .X(net486));
 sky130_fd_sc_hd__bufbuf_16 hold25 (.A(_0850_),
    .X(net487));
 sky130_fd_sc_hd__bufbuf_16 hold26 (.A(net584),
    .X(net488));
 sky130_fd_sc_hd__bufbuf_16 hold27 (.A(net577),
    .X(net489));
 sky130_fd_sc_hd__bufbuf_16 hold28 (.A(_0884_),
    .X(net490));
 sky130_fd_sc_hd__bufbuf_16 hold29 (.A(_2412_),
    .X(net491));
 sky130_fd_sc_hd__bufbuf_16 hold30 (.A(_0457_),
    .X(net492));
 sky130_fd_sc_hd__bufbuf_16 hold31 (.A(net500),
    .X(net493));
 sky130_fd_sc_hd__bufbuf_16 hold32 (.A(net502),
    .X(net494));
 sky130_fd_sc_hd__bufbuf_16 hold33 (.A(net504),
    .X(net495));
 sky130_fd_sc_hd__bufbuf_16 hold34 (.A(_0612_),
    .X(net496));
 sky130_fd_sc_hd__bufbuf_16 hold35 (.A(net526),
    .X(net497));
 sky130_fd_sc_hd__bufbuf_16 hold36 (.A(net623),
    .X(net498));
 sky130_fd_sc_hd__bufbuf_16 hold37 (.A(_0707_),
    .X(net499));
 sky130_fd_sc_hd__bufbuf_16 hold38 (.A(\hkspi.odata[2] ),
    .X(net500));
 sky130_fd_sc_hd__bufbuf_16 hold39 (.A(net493),
    .X(net501));
 sky130_fd_sc_hd__bufbuf_16 hold40 (.A(_1469_),
    .X(net502));
 sky130_fd_sc_hd__bufbuf_16 hold41 (.A(net494),
    .X(net503));
 sky130_fd_sc_hd__bufbuf_16 hold42 (.A(net393),
    .X(net504));
 sky130_fd_sc_hd__bufbuf_16 hold43 (.A(net495),
    .X(net505));
 sky130_fd_sc_hd__bufbuf_16 hold44 (.A(_0532_),
    .X(net506));
 sky130_fd_sc_hd__bufbuf_16 hold45 (.A(net1273),
    .X(net507));
 sky130_fd_sc_hd__bufbuf_16 hold46 (.A(net561),
    .X(net508));
 sky130_fd_sc_hd__bufbuf_16 hold47 (.A(net364),
    .X(net509));
 sky130_fd_sc_hd__bufbuf_16 hold48 (.A(_2429_),
    .X(net510));
 sky130_fd_sc_hd__bufbuf_16 hold49 (.A(_0588_),
    .X(net511));
 sky130_fd_sc_hd__bufbuf_16 hold50 (.A(\hkspi.addr[6] ),
    .X(net512));
 sky130_fd_sc_hd__bufbuf_16 hold51 (.A(net686),
    .X(net513));
 sky130_fd_sc_hd__bufbuf_16 hold52 (.A(net656),
    .X(net514));
 sky130_fd_sc_hd__bufbuf_16 hold53 (.A(_0864_),
    .X(net515));
 sky130_fd_sc_hd__bufbuf_16 hold54 (.A(_0875_),
    .X(net516));
 sky130_fd_sc_hd__bufbuf_16 hold55 (.A(_2440_),
    .X(net517));
 sky130_fd_sc_hd__bufbuf_16 hold56 (.A(_0676_),
    .X(net518));
 sky130_fd_sc_hd__bufbuf_16 hold57 (.A(net572),
    .X(net519));
 sky130_fd_sc_hd__bufbuf_16 hold58 (.A(_0839_),
    .X(net520));
 sky130_fd_sc_hd__bufbuf_16 hold59 (.A(net636),
    .X(net521));
 sky130_fd_sc_hd__bufbuf_16 hold60 (.A(net638),
    .X(net522));
 sky130_fd_sc_hd__bufbuf_16 hold61 (.A(_0954_),
    .X(net523));
 sky130_fd_sc_hd__bufbuf_16 hold62 (.A(_2446_),
    .X(net524));
 sky130_fd_sc_hd__bufbuf_16 hold63 (.A(_0724_),
    .X(net525));
 sky130_fd_sc_hd__bufbuf_16 hold64 (.A(\hkspi.odata[1] ),
    .X(net526));
 sky130_fd_sc_hd__bufbuf_16 hold65 (.A(net497),
    .X(net527));
 sky130_fd_sc_hd__bufbuf_16 hold66 (.A(net622),
    .X(net528));
 sky130_fd_sc_hd__bufbuf_16 hold67 (.A(net498),
    .X(net529));
 sky130_fd_sc_hd__bufbuf_16 hold68 (.A(_0691_),
    .X(net530));
 sky130_fd_sc_hd__bufbuf_16 hold69 (.A(net594),
    .X(net531));
 sky130_fd_sc_hd__bufbuf_16 hold70 (.A(net596),
    .X(net532));
 sky130_fd_sc_hd__bufbuf_16 hold71 (.A(net387),
    .X(net533));
 sky130_fd_sc_hd__bufbuf_16 hold72 (.A(_0174_),
    .X(net534));
 sky130_fd_sc_hd__bufbuf_16 hold73 (.A(\hkspi.odata[5] ),
    .X(net535));
 sky130_fd_sc_hd__bufbuf_16 hold74 (.A(net467),
    .X(net536));
 sky130_fd_sc_hd__bufbuf_16 hold75 (.A(_1472_),
    .X(net537));
 sky130_fd_sc_hd__bufbuf_16 hold76 (.A(net468),
    .X(net538));
 sky130_fd_sc_hd__bufbuf_16 hold77 (.A(net377),
    .X(net539));
 sky130_fd_sc_hd__bufbuf_16 hold78 (.A(net469),
    .X(net540));
 sky130_fd_sc_hd__bufbuf_16 hold79 (.A(_0455_),
    .X(net541));
 sky130_fd_sc_hd__bufbuf_16 hold80 (.A(\hkspi.addr[0] ),
    .X(net542));
 sky130_fd_sc_hd__bufbuf_16 hold81 (.A(_0859_),
    .X(net543));
 sky130_fd_sc_hd__bufbuf_16 hold82 (.A(net820),
    .X(net544));
 sky130_fd_sc_hd__bufbuf_16 hold83 (.A(_0877_),
    .X(net545));
 sky130_fd_sc_hd__bufbuf_16 hold84 (.A(_0879_),
    .X(net546));
 sky130_fd_sc_hd__bufbuf_16 hold85 (.A(_0900_),
    .X(net547));
 sky130_fd_sc_hd__bufbuf_16 hold86 (.A(_2443_),
    .X(net548));
 sky130_fd_sc_hd__bufbuf_16 hold87 (.A(_0703_),
    .X(net549));
 sky130_fd_sc_hd__bufbuf_16 hold88 (.A(net747),
    .X(net550));
 sky130_fd_sc_hd__bufbuf_16 hold89 (.A(_0855_),
    .X(net551));
 sky130_fd_sc_hd__bufbuf_16 hold90 (.A(_0856_),
    .X(net552));
 sky130_fd_sc_hd__bufbuf_16 hold91 (.A(_0862_),
    .X(net553));
 sky130_fd_sc_hd__bufbuf_16 hold92 (.A(_0865_),
    .X(net554));
 sky130_fd_sc_hd__bufbuf_16 hold93 (.A(_2438_),
    .X(net555));
 sky130_fd_sc_hd__bufbuf_16 hold94 (.A(_0660_),
    .X(net556));
 sky130_fd_sc_hd__bufbuf_16 hold95 (.A(\mgmt_gpio_data[37] ),
    .X(net557));
 sky130_fd_sc_hd__bufbuf_16 hold96 (.A(_0433_),
    .X(net558));
 sky130_fd_sc_hd__bufbuf_16 hold97 (.A(net1272),
    .X(net559));
 sky130_fd_sc_hd__bufbuf_16 hold98 (.A(net507),
    .X(net560));
 sky130_fd_sc_hd__bufbuf_16 hold99 (.A(_1464_),
    .X(net561));
 sky130_fd_sc_hd__bufbuf_16 hold100 (.A(net508),
    .X(net562));
 sky130_fd_sc_hd__bufbuf_16 hold101 (.A(_2424_),
    .X(net563));
 sky130_fd_sc_hd__bufbuf_16 hold102 (.A(_0553_),
    .X(net564));
 sky130_fd_sc_hd__bufbuf_16 hold103 (.A(\hkspi.addr[4] ),
    .X(net565));
 sky130_fd_sc_hd__bufbuf_16 hold104 (.A(_0842_),
    .X(net566));
 sky130_fd_sc_hd__bufbuf_16 hold105 (.A(net607),
    .X(net567));
 sky130_fd_sc_hd__bufbuf_16 hold106 (.A(_0867_),
    .X(net568));
 sky130_fd_sc_hd__bufbuf_16 hold107 (.A(_0903_),
    .X(net569));
 sky130_fd_sc_hd__bufbuf_16 hold108 (.A(_0904_),
    .X(net570));
 sky130_fd_sc_hd__bufbuf_16 hold109 (.A(_0449_),
    .X(net571));
 sky130_fd_sc_hd__bufbuf_16 hold110 (.A(\hkspi.addr[3] ),
    .X(net572));
 sky130_fd_sc_hd__bufbuf_16 hold111 (.A(net519),
    .X(net573));
 sky130_fd_sc_hd__bufbuf_16 hold112 (.A(_0852_),
    .X(net574));
 sky130_fd_sc_hd__bufbuf_16 hold113 (.A(_0853_),
    .X(net575));
 sky130_fd_sc_hd__bufbuf_16 hold114 (.A(_0854_),
    .X(net576));
 sky130_fd_sc_hd__bufbuf_16 hold115 (.A(_0881_),
    .X(net577));
 sky130_fd_sc_hd__bufbuf_16 hold116 (.A(net489),
    .X(net578));
 sky130_fd_sc_hd__bufbuf_16 hold117 (.A(_0888_),
    .X(net579));
 sky130_fd_sc_hd__bufbuf_16 hold118 (.A(_0583_),
    .X(net580));
 sky130_fd_sc_hd__bufbuf_16 hold119 (.A(\gpio_configure[31][5] ),
    .X(net581));
 sky130_fd_sc_hd__bufbuf_16 hold120 (.A(_0695_),
    .X(net582));
 sky130_fd_sc_hd__bufbuf_16 hold121 (.A(\wbbd_addr[2] ),
    .X(net583));
 sky130_fd_sc_hd__bufbuf_16 hold122 (.A(_0851_),
    .X(net584));
 sky130_fd_sc_hd__bufbuf_16 hold123 (.A(net488),
    .X(net585));
 sky130_fd_sc_hd__bufbuf_16 hold124 (.A(_0873_),
    .X(net586));
 sky130_fd_sc_hd__bufbuf_16 hold125 (.A(_0910_),
    .X(net587));
 sky130_fd_sc_hd__bufbuf_16 hold126 (.A(_0930_),
    .X(net588));
 sky130_fd_sc_hd__bufbuf_16 hold127 (.A(_0684_),
    .X(net589));
 sky130_fd_sc_hd__bufbuf_16 hold128 (.A(net666),
    .X(net590));
 sky130_fd_sc_hd__bufbuf_16 hold129 (.A(net668),
    .X(net591));
 sky130_fd_sc_hd__bufbuf_16 hold130 (.A(net670),
    .X(net592));
 sky130_fd_sc_hd__bufbuf_16 hold131 (.A(net1697),
    .X(net593));
 sky130_fd_sc_hd__bufbuf_16 hold132 (.A(\hkspi.odata[3] ),
    .X(net594));
 sky130_fd_sc_hd__bufbuf_16 hold133 (.A(net531),
    .X(net595));
 sky130_fd_sc_hd__bufbuf_16 hold134 (.A(net614),
    .X(net596));
 sky130_fd_sc_hd__bufbuf_16 hold135 (.A(net532),
    .X(net597));
 sky130_fd_sc_hd__bufbuf_16 hold136 (.A(net385),
    .X(net598));
 sky130_fd_sc_hd__bufbuf_16 hold137 (.A(_0416_),
    .X(net599));
 sky130_fd_sc_hd__bufbuf_16 hold138 (.A(\gpio_configure[19][5] ),
    .X(net600));
 sky130_fd_sc_hd__bufbuf_16 hold139 (.A(_0599_),
    .X(net601));
 sky130_fd_sc_hd__bufbuf_16 hold140 (.A(\gpio_configure[37][3] ),
    .X(net602));
 sky130_fd_sc_hd__bufbuf_16 hold141 (.A(_0741_),
    .X(net603));
 sky130_fd_sc_hd__bufbuf_16 hold142 (.A(\gpio_configure[33][5] ),
    .X(net604));
 sky130_fd_sc_hd__bufbuf_16 hold143 (.A(_0711_),
    .X(net605));
 sky130_fd_sc_hd__bufbuf_16 hold144 (.A(\wbbd_addr[5] ),
    .X(net606));
 sky130_fd_sc_hd__bufbuf_16 hold145 (.A(_0843_),
    .X(net607));
 sky130_fd_sc_hd__bufbuf_16 hold146 (.A(net567),
    .X(net608));
 sky130_fd_sc_hd__bufbuf_16 hold147 (.A(_0849_),
    .X(net609));
 sky130_fd_sc_hd__bufbuf_16 hold148 (.A(_0948_),
    .X(net610));
 sky130_fd_sc_hd__bufbuf_16 hold149 (.A(_2431_),
    .X(net611));
 sky130_fd_sc_hd__bufbuf_16 hold150 (.A(_0605_),
    .X(net612));
 sky130_fd_sc_hd__bufbuf_16 hold151 (.A(\wbbd_data[3] ),
    .X(net613));
 sky130_fd_sc_hd__bufbuf_16 hold152 (.A(_1470_),
    .X(net614));
 sky130_fd_sc_hd__bufbuf_16 hold153 (.A(_0733_),
    .X(net615));
 sky130_fd_sc_hd__bufbuf_16 hold154 (.A(wbbd_write),
    .X(net616));
 sky130_fd_sc_hd__bufbuf_16 hold155 (.A(_1463_),
    .X(net617));
 sky130_fd_sc_hd__bufbuf_16 hold156 (.A(_0645_),
    .X(net618));
 sky130_fd_sc_hd__bufbuf_16 hold157 (.A(\gpio_configure[28][2] ),
    .X(net619));
 sky130_fd_sc_hd__bufbuf_16 hold158 (.A(_0668_),
    .X(net620));
 sky130_fd_sc_hd__bufbuf_16 hold159 (.A(\wbbd_data[1] ),
    .X(net621));
 sky130_fd_sc_hd__bufbuf_16 hold160 (.A(_1468_),
    .X(net622));
 sky130_fd_sc_hd__bufbuf_16 hold161 (.A(net528),
    .X(net623));
 sky130_fd_sc_hd__bufbuf_16 hold162 (.A(_0113_),
    .X(net624));
 sky130_fd_sc_hd__bufbuf_16 hold163 (.A(\gpio_configure[26][3] ),
    .X(net625));
 sky130_fd_sc_hd__bufbuf_16 hold164 (.A(_0653_),
    .X(net626));
 sky130_fd_sc_hd__bufbuf_16 hold165 (.A(net232),
    .X(net627));
 sky130_fd_sc_hd__bufbuf_16 hold166 (.A(_0125_),
    .X(net628));
 sky130_fd_sc_hd__bufbuf_16 hold167 (.A(net642),
    .X(net629));
 sky130_fd_sc_hd__bufbuf_16 hold168 (.A(net664),
    .X(net630));
 sky130_fd_sc_hd__bufbuf_16 hold169 (.A(net646),
    .X(net631));
 sky130_fd_sc_hd__bufbuf_16 hold170 (.A(_0415_),
    .X(net632));
 sky130_fd_sc_hd__bufbuf_16 hold171 (.A(\gpio_configure[1][3] ),
    .X(net633));
 sky130_fd_sc_hd__bufbuf_16 hold172 (.A(_0453_),
    .X(net634));
 sky130_fd_sc_hd__bufbuf_16 hold173 (.A(\wbbd_addr[4] ),
    .X(net635));
 sky130_fd_sc_hd__bufbuf_16 hold174 (.A(_0840_),
    .X(net636));
 sky130_fd_sc_hd__bufbuf_16 hold175 (.A(net521),
    .X(net637));
 sky130_fd_sc_hd__bufbuf_16 hold176 (.A(_0898_),
    .X(net638));
 sky130_fd_sc_hd__bufbuf_16 hold177 (.A(net522),
    .X(net639));
 sky130_fd_sc_hd__bufbuf_16 hold178 (.A(_1135_),
    .X(net640));
 sky130_fd_sc_hd__bufbuf_16 hold179 (.A(_0412_),
    .X(net641));
 sky130_fd_sc_hd__bufbuf_16 hold180 (.A(\hkspi.odata[4] ),
    .X(net642));
 sky130_fd_sc_hd__bufbuf_16 hold181 (.A(net629),
    .X(net643));
 sky130_fd_sc_hd__bufbuf_16 hold182 (.A(net663),
    .X(net644));
 sky130_fd_sc_hd__bufbuf_16 hold183 (.A(net630),
    .X(net645));
 sky130_fd_sc_hd__bufbuf_16 hold184 (.A(net380),
    .X(net646));
 sky130_fd_sc_hd__bufbuf_16 hold185 (.A(net631),
    .X(net647));
 sky130_fd_sc_hd__bufbuf_16 hold186 (.A(_0630_),
    .X(net648));
 sky130_fd_sc_hd__bufbuf_16 hold187 (.A(\gpio_configure[15][5] ),
    .X(net649));
 sky130_fd_sc_hd__bufbuf_16 hold188 (.A(_0567_),
    .X(net650));
 sky130_fd_sc_hd__bufbuf_16 hold189 (.A(\gpio_configure[20][4] ),
    .X(net651));
 sky130_fd_sc_hd__bufbuf_16 hold190 (.A(_0606_),
    .X(net652));
 sky130_fd_sc_hd__bufbuf_16 hold191 (.A(\hkspi.addr[5] ),
    .X(net653));
 sky130_fd_sc_hd__bufbuf_16 hold192 (.A(_0846_),
    .X(net654));
 sky130_fd_sc_hd__bufbuf_16 hold193 (.A(_0847_),
    .X(net655));
 sky130_fd_sc_hd__bufbuf_16 hold194 (.A(_0848_),
    .X(net656));
 sky130_fd_sc_hd__bufbuf_16 hold195 (.A(net514),
    .X(net657));
 sky130_fd_sc_hd__bufbuf_16 hold196 (.A(_0923_),
    .X(net658));
 sky130_fd_sc_hd__bufbuf_16 hold197 (.A(_0629_),
    .X(net659));
 sky130_fd_sc_hd__bufbuf_16 hold198 (.A(\gpio_configure[0][3] ),
    .X(net660));
 sky130_fd_sc_hd__bufbuf_16 hold199 (.A(_0445_),
    .X(net661));
 sky130_fd_sc_hd__bufbuf_16 hold200 (.A(\wbbd_data[4] ),
    .X(net662));
 sky130_fd_sc_hd__bufbuf_16 hold201 (.A(_1471_),
    .X(net663));
 sky130_fd_sc_hd__bufbuf_16 hold202 (.A(net644),
    .X(net664));
 sky130_fd_sc_hd__bufbuf_16 hold203 (.A(_0231_),
    .X(net665));
 sky130_fd_sc_hd__bufbuf_16 hold204 (.A(\hkspi.odata[6] ),
    .X(net666));
 sky130_fd_sc_hd__bufbuf_16 hold205 (.A(net590),
    .X(net667));
 sky130_fd_sc_hd__bufbuf_16 hold206 (.A(_1473_),
    .X(net668));
 sky130_fd_sc_hd__bufbuf_16 hold207 (.A(net591),
    .X(net669));
 sky130_fd_sc_hd__bufbuf_16 hold208 (.A(net374),
    .X(net670));
 sky130_fd_sc_hd__bufbuf_16 hold209 (.A(net592),
    .X(net671));
 sky130_fd_sc_hd__bufbuf_16 hold210 (.A(_0736_),
    .X(net672));
 sky130_fd_sc_hd__bufbuf_16 hold211 (.A(\gpio_configure[5][12] ),
    .X(net673));
 sky130_fd_sc_hd__bufbuf_16 hold212 (.A(_0175_),
    .X(net674));
 sky130_fd_sc_hd__bufbuf_16 hold213 (.A(wbbd_busy),
    .X(net675));
 sky130_fd_sc_hd__bufbuf_16 hold214 (.A(net406),
    .X(net676));
 sky130_fd_sc_hd__bufbuf_16 hold215 (.A(net1274),
    .X(net677));
 sky130_fd_sc_hd__bufbuf_16 hold216 (.A(_2410_),
    .X(net678));
 sky130_fd_sc_hd__bufbuf_16 hold217 (.A(_0437_),
    .X(net679));
 sky130_fd_sc_hd__bufbuf_16 hold218 (.A(\gpio_configure[34][4] ),
    .X(net680));
 sky130_fd_sc_hd__bufbuf_16 hold219 (.A(_0718_),
    .X(net681));
 sky130_fd_sc_hd__bufbuf_16 hold220 (.A(\gpio_configure[17][3] ),
    .X(net682));
 sky130_fd_sc_hd__bufbuf_16 hold221 (.A(\gpio_configure[30][3] ),
    .X(net683));
 sky130_fd_sc_hd__bufbuf_16 hold222 (.A(\hkspi.addr[7] ),
    .X(net684));
 sky130_fd_sc_hd__bufbuf_16 hold223 (.A(_0844_),
    .X(net685));
 sky130_fd_sc_hd__bufbuf_16 hold224 (.A(_0845_),
    .X(net686));
 sky130_fd_sc_hd__bufbuf_16 hold225 (.A(_0866_),
    .X(net687));
 sky130_fd_sc_hd__bufbuf_16 hold226 (.A(_0933_),
    .X(net688));
 sky130_fd_sc_hd__bufbuf_16 hold227 (.A(_0110_),
    .X(net689));
 sky130_fd_sc_hd__bufbuf_16 hold228 (.A(\gpio_configure[21][3] ),
    .X(net690));
 sky130_fd_sc_hd__bufbuf_16 hold229 (.A(_0613_),
    .X(net691));
 sky130_fd_sc_hd__bufbuf_16 hold230 (.A(\gpio_configure[17][4] ),
    .X(net692));
 sky130_fd_sc_hd__bufbuf_16 hold231 (.A(_0582_),
    .X(net693));
 sky130_fd_sc_hd__bufbuf_16 hold232 (.A(\gpio_configure[9][11] ),
    .X(net694));
 sky130_fd_sc_hd__bufbuf_16 hold233 (.A(_0210_),
    .X(net695));
 sky130_fd_sc_hd__bufbuf_16 hold234 (.A(\gpio_configure[31][3] ),
    .X(net696));
 sky130_fd_sc_hd__bufbuf_16 hold235 (.A(\gpio_configure[28][3] ),
    .X(net697));
 sky130_fd_sc_hd__bufbuf_16 hold236 (.A(_0669_),
    .X(net698));
 sky130_fd_sc_hd__bufbuf_16 hold237 (.A(\gpio_configure[11][4] ),
    .X(net699));
 sky130_fd_sc_hd__bufbuf_16 hold238 (.A(_0534_),
    .X(net700));
 sky130_fd_sc_hd__bufbuf_16 hold239 (.A(\gpio_configure[27][3] ),
    .X(net701));
 sky130_fd_sc_hd__bufbuf_16 hold240 (.A(\gpio_configure[22][3] ),
    .X(net702));
 sky130_fd_sc_hd__bufbuf_16 hold241 (.A(_0621_),
    .X(net703));
 sky130_fd_sc_hd__bufbuf_16 hold242 (.A(\gpio_configure[11][11] ),
    .X(net704));
 sky130_fd_sc_hd__bufbuf_16 hold243 (.A(_0220_),
    .X(net705));
 sky130_fd_sc_hd__bufbuf_16 hold244 (.A(\gpio_configure[35][3] ),
    .X(net706));
 sky130_fd_sc_hd__bufbuf_16 hold245 (.A(_0725_),
    .X(net707));
 sky130_fd_sc_hd__bufbuf_16 hold246 (.A(\mgmt_gpio_data_buf[6] ),
    .X(net708));
 sky130_fd_sc_hd__bufbuf_16 hold247 (.A(_0440_),
    .X(net709));
 sky130_fd_sc_hd__bufbuf_16 hold248 (.A(\gpio_configure[27][4] ),
    .X(net710));
 sky130_fd_sc_hd__bufbuf_16 hold249 (.A(_0662_),
    .X(net711));
 sky130_fd_sc_hd__bufbuf_16 hold250 (.A(\gpio_configure[29][4] ),
    .X(net712));
 sky130_fd_sc_hd__bufbuf_16 hold251 (.A(_0678_),
    .X(net713));
 sky130_fd_sc_hd__bufbuf_16 hold252 (.A(net233),
    .X(net714));
 sky130_fd_sc_hd__bufbuf_16 hold253 (.A(_0126_),
    .X(net715));
 sky130_fd_sc_hd__bufbuf_16 hold254 (.A(net228),
    .X(net716));
 sky130_fd_sc_hd__bufbuf_16 hold255 (.A(_0279_),
    .X(net717));
 sky130_fd_sc_hd__bufbuf_16 hold256 (.A(\gpio_configure[1][6] ),
    .X(net718));
 sky130_fd_sc_hd__bufbuf_16 hold257 (.A(_0456_),
    .X(net719));
 sky130_fd_sc_hd__bufbuf_16 hold258 (.A(\gpio_configure[19][3] ),
    .X(net720));
 sky130_fd_sc_hd__bufbuf_16 hold259 (.A(_0597_),
    .X(net721));
 sky130_fd_sc_hd__bufbuf_16 hold260 (.A(\gpio_configure[15][6] ),
    .X(net722));
 sky130_fd_sc_hd__bufbuf_16 hold261 (.A(_0568_),
    .X(net723));
 sky130_fd_sc_hd__bufbuf_16 hold262 (.A(\gpio_configure[11][3] ),
    .X(net724));
 sky130_fd_sc_hd__bufbuf_16 hold263 (.A(_0533_),
    .X(net725));
 sky130_fd_sc_hd__bufbuf_16 hold264 (.A(\gpio_configure[2][5] ),
    .X(net726));
 sky130_fd_sc_hd__bufbuf_16 hold265 (.A(_0463_),
    .X(net727));
 sky130_fd_sc_hd__bufbuf_16 hold266 (.A(\gpio_configure[24][3] ),
    .X(net728));
 sky130_fd_sc_hd__bufbuf_16 hold267 (.A(\mgmt_gpio_data_buf[12] ),
    .X(net729));
 sky130_fd_sc_hd__bufbuf_16 hold268 (.A(_0134_),
    .X(net730));
 sky130_fd_sc_hd__bufbuf_16 hold269 (.A(\gpio_configure[30][4] ),
    .X(net731));
 sky130_fd_sc_hd__bufbuf_16 hold270 (.A(_0686_),
    .X(net732));
 sky130_fd_sc_hd__bufbuf_16 hold271 (.A(\gpio_configure[24][4] ),
    .X(net733));
 sky130_fd_sc_hd__bufbuf_16 hold272 (.A(_0638_),
    .X(net734));
 sky130_fd_sc_hd__bufbuf_16 hold273 (.A(net226),
    .X(net735));
 sky130_fd_sc_hd__bufbuf_16 hold274 (.A(_0277_),
    .X(net736));
 sky130_fd_sc_hd__bufbuf_16 hold275 (.A(\gpio_configure[19][4] ),
    .X(net737));
 sky130_fd_sc_hd__bufbuf_16 hold276 (.A(_0598_),
    .X(net738));
 sky130_fd_sc_hd__bufbuf_16 hold277 (.A(\gpio_configure[0][4] ),
    .X(net739));
 sky130_fd_sc_hd__bufbuf_16 hold278 (.A(_0446_),
    .X(net740));
 sky130_fd_sc_hd__bufbuf_16 hold279 (.A(\gpio_configure[16][4] ),
    .X(net741));
 sky130_fd_sc_hd__bufbuf_16 hold280 (.A(_0574_),
    .X(net742));
 sky130_fd_sc_hd__bufbuf_16 hold281 (.A(\mgmt_gpio_data[15] ),
    .X(net743));
 sky130_fd_sc_hd__bufbuf_16 hold282 (.A(_0121_),
    .X(net744));
 sky130_fd_sc_hd__bufbuf_16 hold283 (.A(\gpio_configure[14][4] ),
    .X(net745));
 sky130_fd_sc_hd__bufbuf_16 hold284 (.A(_0558_),
    .X(net746));
 sky130_fd_sc_hd__bufbuf_16 hold285 (.A(\wbbd_addr[3] ),
    .X(net747));
 sky130_fd_sc_hd__bufbuf_16 hold286 (.A(net550),
    .X(net748));
 sky130_fd_sc_hd__bufbuf_16 hold287 (.A(_0905_),
    .X(net749));
 sky130_fd_sc_hd__bufbuf_16 hold288 (.A(_0906_),
    .X(net750));
 sky130_fd_sc_hd__bufbuf_16 hold289 (.A(_0651_),
    .X(net751));
 sky130_fd_sc_hd__bufbuf_16 hold290 (.A(\gpio_configure[29][3] ),
    .X(net752));
 sky130_fd_sc_hd__bufbuf_16 hold291 (.A(\gpio_configure[13][6] ),
    .X(net753));
 sky130_fd_sc_hd__bufbuf_16 hold292 (.A(_0552_),
    .X(net754));
 sky130_fd_sc_hd__bufbuf_16 hold293 (.A(\mgmt_gpio_data_buf[4] ),
    .X(net755));
 sky130_fd_sc_hd__bufbuf_16 hold294 (.A(_0438_),
    .X(net756));
 sky130_fd_sc_hd__bufbuf_16 hold295 (.A(\gpio_configure[13][3] ),
    .X(net757));
 sky130_fd_sc_hd__bufbuf_16 hold296 (.A(_0549_),
    .X(net758));
 sky130_fd_sc_hd__bufbuf_16 hold297 (.A(\gpio_configure[21][4] ),
    .X(net759));
 sky130_fd_sc_hd__bufbuf_16 hold298 (.A(_0614_),
    .X(net760));
 sky130_fd_sc_hd__bufbuf_16 hold299 (.A(\gpio_configure[28][4] ),
    .X(net761));
 sky130_fd_sc_hd__bufbuf_16 hold300 (.A(_0670_),
    .X(net762));
 sky130_fd_sc_hd__bufbuf_16 hold301 (.A(\gpio_configure[9][4] ),
    .X(net763));
 sky130_fd_sc_hd__bufbuf_16 hold302 (.A(_0518_),
    .X(net764));
 sky130_fd_sc_hd__bufbuf_16 hold303 (.A(\gpio_configure[18][4] ),
    .X(net765));
 sky130_fd_sc_hd__bufbuf_16 hold304 (.A(_0590_),
    .X(net766));
 sky130_fd_sc_hd__bufbuf_16 hold305 (.A(\gpio_configure[4][11] ),
    .X(net767));
 sky130_fd_sc_hd__bufbuf_16 hold306 (.A(_0161_),
    .X(net768));
 sky130_fd_sc_hd__bufbuf_16 hold307 (.A(\gpio_configure[27][6] ),
    .X(net769));
 sky130_fd_sc_hd__bufbuf_16 hold308 (.A(_0664_),
    .X(net770));
 sky130_fd_sc_hd__bufbuf_16 hold309 (.A(net230),
    .X(net771));
 sky130_fd_sc_hd__bufbuf_16 hold310 (.A(_0123_),
    .X(net772));
 sky130_fd_sc_hd__bufbuf_16 hold311 (.A(\gpio_configure[9][1] ),
    .X(net773));
 sky130_fd_sc_hd__bufbuf_16 hold312 (.A(\gpio_configure[16][11] ),
    .X(net774));
 sky130_fd_sc_hd__bufbuf_16 hold313 (.A(_0235_),
    .X(net775));
 sky130_fd_sc_hd__bufbuf_16 hold314 (.A(\gpio_configure[16][1] ),
    .X(net776));
 sky130_fd_sc_hd__bufbuf_16 hold315 (.A(\gpio_configure[7][1] ),
    .X(net777));
 sky130_fd_sc_hd__bufbuf_16 hold316 (.A(_0499_),
    .X(net778));
 sky130_fd_sc_hd__bufbuf_16 hold317 (.A(net1728),
    .X(net779));
 sky130_fd_sc_hd__bufbuf_16 hold318 (.A(_0290_),
    .X(net780));
 sky130_fd_sc_hd__bufbuf_16 hold319 (.A(net237),
    .X(net781));
 sky130_fd_sc_hd__bufbuf_16 hold320 (.A(_0129_),
    .X(net782));
 sky130_fd_sc_hd__bufbuf_16 hold321 (.A(\mgmt_gpio_data_buf[9] ),
    .X(net783));
 sky130_fd_sc_hd__bufbuf_16 hold322 (.A(_0131_),
    .X(net784));
 sky130_fd_sc_hd__bufbuf_16 hold323 (.A(\gpio_configure[3][9] ),
    .X(net785));
 sky130_fd_sc_hd__bufbuf_16 hold324 (.A(_0154_),
    .X(net786));
 sky130_fd_sc_hd__bufbuf_16 hold325 (.A(\wbbd_addr[1] ),
    .X(net787));
 sky130_fd_sc_hd__bufbuf_16 hold326 (.A(_0858_),
    .X(net788));
 sky130_fd_sc_hd__bufbuf_16 hold327 (.A(net480),
    .X(net789));
 sky130_fd_sc_hd__bufbuf_16 hold328 (.A(_0931_),
    .X(net790));
 sky130_fd_sc_hd__bufbuf_16 hold329 (.A(_0956_),
    .X(net791));
 sky130_fd_sc_hd__bufbuf_16 hold330 (.A(_1095_),
    .X(net792));
 sky130_fd_sc_hd__bufbuf_16 hold331 (.A(_0223_),
    .X(net793));
 sky130_fd_sc_hd__bufbuf_16 hold332 (.A(\gpio_configure[10][1] ),
    .X(net794));
 sky130_fd_sc_hd__bufbuf_16 hold333 (.A(\gpio_configure[14][1] ),
    .X(net795));
 sky130_fd_sc_hd__bufbuf_16 hold334 (.A(_0555_),
    .X(net796));
 sky130_fd_sc_hd__bufbuf_16 hold335 (.A(\gpio_configure[9][7] ),
    .X(net797));
 sky130_fd_sc_hd__bufbuf_16 hold336 (.A(_0521_),
    .X(net798));
 sky130_fd_sc_hd__bufbuf_16 hold337 (.A(\gpio_configure[8][7] ),
    .X(net799));
 sky130_fd_sc_hd__bufbuf_16 hold338 (.A(_0513_),
    .X(net800));
 sky130_fd_sc_hd__bufbuf_16 hold339 (.A(\gpio_configure[29][1] ),
    .X(net801));
 sky130_fd_sc_hd__bufbuf_16 hold340 (.A(\gpio_configure[2][3] ),
    .X(net802));
 sky130_fd_sc_hd__bufbuf_16 hold341 (.A(\gpio_configure[34][1] ),
    .X(net803));
 sky130_fd_sc_hd__bufbuf_16 hold342 (.A(\gpio_configure[25][9] ),
    .X(net804));
 sky130_fd_sc_hd__bufbuf_16 hold343 (.A(_0258_),
    .X(net805));
 sky130_fd_sc_hd__bufbuf_16 hold344 (.A(\gpio_configure[5][9] ),
    .X(net806));
 sky130_fd_sc_hd__bufbuf_16 hold345 (.A(_0172_),
    .X(net807));
 sky130_fd_sc_hd__bufbuf_16 hold346 (.A(\gpio_configure[23][1] ),
    .X(net808));
 sky130_fd_sc_hd__bufbuf_16 hold347 (.A(\gpio_configure[7][7] ),
    .X(net809));
 sky130_fd_sc_hd__bufbuf_16 hold348 (.A(_0505_),
    .X(net810));
 sky130_fd_sc_hd__bufbuf_16 hold349 (.A(\gpio_configure[36][7] ),
    .X(net811));
 sky130_fd_sc_hd__bufbuf_16 hold350 (.A(_0737_),
    .X(net812));
 sky130_fd_sc_hd__bufbuf_16 hold351 (.A(\gpio_configure[18][1] ),
    .X(net813));
 sky130_fd_sc_hd__bufbuf_16 hold352 (.A(_0587_),
    .X(net814));
 sky130_fd_sc_hd__bufbuf_16 hold353 (.A(net302),
    .X(net815));
 sky130_fd_sc_hd__bufbuf_16 hold354 (.A(_0410_),
    .X(net816));
 sky130_fd_sc_hd__bufbuf_16 hold355 (.A(\mgmt_gpio_data_buf[15] ),
    .X(net817));
 sky130_fd_sc_hd__bufbuf_16 hold356 (.A(_0137_),
    .X(net818));
 sky130_fd_sc_hd__bufbuf_16 hold357 (.A(\wbbd_addr[0] ),
    .X(net819));
 sky130_fd_sc_hd__bufbuf_16 hold358 (.A(_0860_),
    .X(net820));
 sky130_fd_sc_hd__bufbuf_16 hold359 (.A(_0420_),
    .X(net821));
 sky130_fd_sc_hd__bufbuf_16 hold360 (.A(\gpio_configure[30][1] ),
    .X(net822));
 sky130_fd_sc_hd__bufbuf_16 hold361 (.A(\gpio_configure[20][1] ),
    .X(net823));
 sky130_fd_sc_hd__bufbuf_16 hold362 (.A(\gpio_configure[35][1] ),
    .X(net824));
 sky130_fd_sc_hd__bufbuf_16 hold363 (.A(\gpio_configure[25][7] ),
    .X(net825));
 sky130_fd_sc_hd__bufbuf_16 hold364 (.A(_0649_),
    .X(net826));
 sky130_fd_sc_hd__bufbuf_16 hold365 (.A(\gpio_configure[25][1] ),
    .X(net827));
 sky130_fd_sc_hd__bufbuf_16 hold366 (.A(\gpio_configure[4][7] ),
    .X(net828));
 sky130_fd_sc_hd__bufbuf_16 hold367 (.A(_0481_),
    .X(net829));
 sky130_fd_sc_hd__bufbuf_16 hold368 (.A(\gpio_configure[14][7] ),
    .X(net830));
 sky130_fd_sc_hd__bufbuf_16 hold369 (.A(_0561_),
    .X(net831));
 sky130_fd_sc_hd__bufbuf_16 hold370 (.A(\gpio_configure[16][7] ),
    .X(net832));
 sky130_fd_sc_hd__bufbuf_16 hold371 (.A(_0577_),
    .X(net833));
 sky130_fd_sc_hd__bufbuf_16 hold372 (.A(net283),
    .X(net834));
 sky130_fd_sc_hd__bufbuf_16 hold373 (.A(\gpio_configure[22][1] ),
    .X(net835));
 sky130_fd_sc_hd__bufbuf_16 hold374 (.A(\gpio_configure[9][5] ),
    .X(net836));
 sky130_fd_sc_hd__bufbuf_16 hold375 (.A(_0519_),
    .X(net837));
 sky130_fd_sc_hd__bufbuf_16 hold376 (.A(\gpio_configure[36][11] ),
    .X(net838));
 sky130_fd_sc_hd__bufbuf_16 hold377 (.A(\gpio_configure[3][7] ),
    .X(net839));
 sky130_fd_sc_hd__bufbuf_16 hold378 (.A(_0473_),
    .X(net840));
 sky130_fd_sc_hd__bufbuf_16 hold379 (.A(\gpio_configure[11][1] ),
    .X(net841));
 sky130_fd_sc_hd__bufbuf_16 hold380 (.A(\gpio_configure[18][7] ),
    .X(net842));
 sky130_fd_sc_hd__bufbuf_16 hold381 (.A(_0593_),
    .X(net843));
 sky130_fd_sc_hd__bufbuf_16 hold382 (.A(\gpio_configure[13][1] ),
    .X(net844));
 sky130_fd_sc_hd__bufbuf_16 hold383 (.A(\gpio_configure[37][1] ),
    .X(net845));
 sky130_fd_sc_hd__bufbuf_16 hold384 (.A(net234),
    .X(net846));
 sky130_fd_sc_hd__bufbuf_16 hold385 (.A(_0127_),
    .X(net847));
 sky130_fd_sc_hd__bufbuf_16 hold386 (.A(\gpio_configure[5][7] ),
    .X(net848));
 sky130_fd_sc_hd__bufbuf_16 hold387 (.A(_0489_),
    .X(net849));
 sky130_fd_sc_hd__bufbuf_16 hold388 (.A(\gpio_configure[34][5] ),
    .X(net850));
 sky130_fd_sc_hd__bufbuf_16 hold389 (.A(_0719_),
    .X(net851));
 sky130_fd_sc_hd__bufbuf_16 hold390 (.A(\gpio_configure[37][7] ),
    .X(net852));
 sky130_fd_sc_hd__bufbuf_16 hold391 (.A(_0745_),
    .X(net853));
 sky130_fd_sc_hd__bufbuf_16 hold392 (.A(\gpio_configure[1][1] ),
    .X(net854));
 sky130_fd_sc_hd__bufbuf_16 hold393 (.A(\gpio_configure[3][5] ),
    .X(net855));
 sky130_fd_sc_hd__bufbuf_16 hold394 (.A(_0471_),
    .X(net856));
 sky130_fd_sc_hd__bufbuf_16 hold395 (.A(\gpio_configure[0][1] ),
    .X(net857));
 sky130_fd_sc_hd__bufbuf_16 hold396 (.A(_0443_),
    .X(net858));
 sky130_fd_sc_hd__bufbuf_16 hold397 (.A(\gpio_configure[17][1] ),
    .X(net859));
 sky130_fd_sc_hd__bufbuf_16 hold398 (.A(\gpio_configure[11][7] ),
    .X(net860));
 sky130_fd_sc_hd__bufbuf_16 hold399 (.A(_0537_),
    .X(net861));
 sky130_fd_sc_hd__bufbuf_16 hold400 (.A(\gpio_configure[28][7] ),
    .X(net862));
 sky130_fd_sc_hd__bufbuf_16 hold401 (.A(_0673_),
    .X(net863));
 sky130_fd_sc_hd__bufbuf_16 hold402 (.A(\gpio_configure[26][5] ),
    .X(net864));
 sky130_fd_sc_hd__bufbuf_16 hold403 (.A(_0655_),
    .X(net865));
 sky130_fd_sc_hd__bufbuf_16 hold404 (.A(\gpio_configure[8][5] ),
    .X(net866));
 sky130_fd_sc_hd__bufbuf_16 hold405 (.A(_0511_),
    .X(net867));
 sky130_fd_sc_hd__bufbuf_16 hold406 (.A(\gpio_configure[22][7] ),
    .X(net868));
 sky130_fd_sc_hd__bufbuf_16 hold407 (.A(_0625_),
    .X(net869));
 sky130_fd_sc_hd__bufbuf_16 hold408 (.A(net281),
    .X(net870));
 sky130_fd_sc_hd__bufbuf_16 hold409 (.A(\gpio_configure[16][5] ),
    .X(net871));
 sky130_fd_sc_hd__bufbuf_16 hold410 (.A(_0575_),
    .X(net872));
 sky130_fd_sc_hd__bufbuf_16 hold411 (.A(\mgmt_gpio_data_buf[13] ),
    .X(net873));
 sky130_fd_sc_hd__bufbuf_16 hold412 (.A(_0135_),
    .X(net874));
 sky130_fd_sc_hd__bufbuf_16 hold413 (.A(\gpio_configure[19][9] ),
    .X(net875));
 sky130_fd_sc_hd__bufbuf_16 hold414 (.A(_0328_),
    .X(net876));
 sky130_fd_sc_hd__bufbuf_16 hold415 (.A(\gpio_configure[28][1] ),
    .X(net877));
 sky130_fd_sc_hd__bufbuf_16 hold416 (.A(_0667_),
    .X(net878));
 sky130_fd_sc_hd__bufbuf_16 hold417 (.A(net290),
    .X(net879));
 sky130_fd_sc_hd__bufbuf_16 hold418 (.A(\gpio_configure[30][7] ),
    .X(net880));
 sky130_fd_sc_hd__bufbuf_16 hold419 (.A(_0689_),
    .X(net881));
 sky130_fd_sc_hd__bufbuf_16 hold420 (.A(\gpio_configure[27][1] ),
    .X(net882));
 sky130_fd_sc_hd__bufbuf_16 hold421 (.A(\gpio_configure[20][7] ),
    .X(net883));
 sky130_fd_sc_hd__bufbuf_16 hold422 (.A(_0609_),
    .X(net884));
 sky130_fd_sc_hd__bufbuf_16 hold423 (.A(\gpio_configure[23][7] ),
    .X(net885));
 sky130_fd_sc_hd__bufbuf_16 hold424 (.A(_0633_),
    .X(net886));
 sky130_fd_sc_hd__bufbuf_16 hold425 (.A(clk2_output_dest),
    .X(net887));
 sky130_fd_sc_hd__bufbuf_16 hold426 (.A(_0424_),
    .X(net888));
 sky130_fd_sc_hd__bufbuf_16 hold427 (.A(\gpio_configure[35][7] ),
    .X(net889));
 sky130_fd_sc_hd__bufbuf_16 hold428 (.A(_0729_),
    .X(net890));
 sky130_fd_sc_hd__bufbuf_16 hold429 (.A(\mgmt_gpio_data_buf[7] ),
    .X(net891));
 sky130_fd_sc_hd__bufbuf_16 hold430 (.A(_0441_),
    .X(net892));
 sky130_fd_sc_hd__bufbuf_16 hold431 (.A(\gpio_configure[26][2] ),
    .X(net893));
 sky130_fd_sc_hd__bufbuf_16 hold432 (.A(_0652_),
    .X(net894));
 sky130_fd_sc_hd__bufbuf_16 hold433 (.A(\gpio_configure[13][4] ),
    .X(net895));
 sky130_fd_sc_hd__bufbuf_16 hold434 (.A(_0550_),
    .X(net896));
 sky130_fd_sc_hd__bufbuf_16 hold435 (.A(\gpio_configure[29][7] ),
    .X(net897));
 sky130_fd_sc_hd__bufbuf_16 hold436 (.A(_0681_),
    .X(net898));
 sky130_fd_sc_hd__bufbuf_16 hold437 (.A(\gpio_configure[34][2] ),
    .X(net899));
 sky130_fd_sc_hd__bufbuf_16 hold438 (.A(_0716_),
    .X(net900));
 sky130_fd_sc_hd__bufbuf_16 hold439 (.A(\gpio_configure[34][7] ),
    .X(net901));
 sky130_fd_sc_hd__bufbuf_16 hold440 (.A(_0721_),
    .X(net902));
 sky130_fd_sc_hd__bufbuf_16 hold441 (.A(\gpio_configure[21][1] ),
    .X(net903));
 sky130_fd_sc_hd__bufbuf_16 hold442 (.A(\gpio_configure[10][5] ),
    .X(net904));
 sky130_fd_sc_hd__bufbuf_16 hold443 (.A(_0527_),
    .X(net905));
 sky130_fd_sc_hd__bufbuf_16 hold444 (.A(\gpio_configure[6][4] ),
    .X(net906));
 sky130_fd_sc_hd__bufbuf_16 hold445 (.A(_0494_),
    .X(net907));
 sky130_fd_sc_hd__bufbuf_16 hold446 (.A(net244),
    .X(net908));
 sky130_fd_sc_hd__bufbuf_16 hold447 (.A(_0283_),
    .X(net909));
 sky130_fd_sc_hd__bufbuf_16 hold448 (.A(\gpio_configure[19][1] ),
    .X(net910));
 sky130_fd_sc_hd__bufbuf_16 hold449 (.A(\gpio_configure[7][5] ),
    .X(net911));
 sky130_fd_sc_hd__bufbuf_16 hold450 (.A(_0503_),
    .X(net912));
 sky130_fd_sc_hd__bufbuf_16 hold451 (.A(\gpio_configure[36][5] ),
    .X(net913));
 sky130_fd_sc_hd__bufbuf_16 hold452 (.A(_0735_),
    .X(net914));
 sky130_fd_sc_hd__bufbuf_16 hold453 (.A(\gpio_configure[21][9] ),
    .X(net915));
 sky130_fd_sc_hd__bufbuf_16 hold454 (.A(_0348_),
    .X(net916));
 sky130_fd_sc_hd__bufbuf_16 hold455 (.A(\gpio_configure[24][1] ),
    .X(net917));
 sky130_fd_sc_hd__bufbuf_16 hold456 (.A(\gpio_configure[25][5] ),
    .X(net918));
 sky130_fd_sc_hd__bufbuf_16 hold457 (.A(_0647_),
    .X(net919));
 sky130_fd_sc_hd__bufbuf_16 hold458 (.A(\mgmt_gpio_data_buf[20] ),
    .X(net920));
 sky130_fd_sc_hd__bufbuf_16 hold459 (.A(_1519_),
    .X(net921));
 sky130_fd_sc_hd__bufbuf_16 hold460 (.A(_0276_),
    .X(net922));
 sky130_fd_sc_hd__bufbuf_16 hold461 (.A(\gpio_configure[36][1] ),
    .X(net923));
 sky130_fd_sc_hd__bufbuf_16 hold462 (.A(\gpio_configure[26][4] ),
    .X(net924));
 sky130_fd_sc_hd__bufbuf_16 hold463 (.A(_0654_),
    .X(net925));
 sky130_fd_sc_hd__bufbuf_16 hold464 (.A(\gpio_configure[37][5] ),
    .X(net926));
 sky130_fd_sc_hd__bufbuf_16 hold465 (.A(_0743_),
    .X(net927));
 sky130_fd_sc_hd__bufbuf_16 hold466 (.A(net287),
    .X(net928));
 sky130_fd_sc_hd__bufbuf_16 hold467 (.A(_0404_),
    .X(net929));
 sky130_fd_sc_hd__bufbuf_16 hold468 (.A(\gpio_configure[4][5] ),
    .X(net930));
 sky130_fd_sc_hd__bufbuf_16 hold469 (.A(_0479_),
    .X(net931));
 sky130_fd_sc_hd__bufbuf_16 hold470 (.A(net278),
    .X(net932));
 sky130_fd_sc_hd__bufbuf_16 hold471 (.A(_0100_),
    .X(net933));
 sky130_fd_sc_hd__bufbuf_16 hold472 (.A(\gpio_configure[21][7] ),
    .X(net934));
 sky130_fd_sc_hd__bufbuf_16 hold473 (.A(_0617_),
    .X(net935));
 sky130_fd_sc_hd__bufbuf_16 hold474 (.A(\gpio_configure[19][7] ),
    .X(net936));
 sky130_fd_sc_hd__bufbuf_16 hold475 (.A(_0601_),
    .X(net937));
 sky130_fd_sc_hd__bufbuf_16 hold476 (.A(\gpio_configure[14][5] ),
    .X(net938));
 sky130_fd_sc_hd__bufbuf_16 hold477 (.A(_0559_),
    .X(net939));
 sky130_fd_sc_hd__bufbuf_16 hold478 (.A(\gpio_configure[15][4] ),
    .X(net940));
 sky130_fd_sc_hd__bufbuf_16 hold479 (.A(_0566_),
    .X(net941));
 sky130_fd_sc_hd__bufbuf_16 hold480 (.A(\gpio_configure[33][7] ),
    .X(net942));
 sky130_fd_sc_hd__bufbuf_16 hold481 (.A(_0713_),
    .X(net943));
 sky130_fd_sc_hd__bufbuf_16 hold482 (.A(\gpio_configure[17][7] ),
    .X(net944));
 sky130_fd_sc_hd__bufbuf_16 hold483 (.A(_0585_),
    .X(net945));
 sky130_fd_sc_hd__bufbuf_16 hold484 (.A(\gpio_configure[26][7] ),
    .X(net946));
 sky130_fd_sc_hd__bufbuf_16 hold485 (.A(_0657_),
    .X(net947));
 sky130_fd_sc_hd__bufbuf_16 hold486 (.A(\gpio_configure[27][7] ),
    .X(net948));
 sky130_fd_sc_hd__bufbuf_16 hold487 (.A(_0665_),
    .X(net949));
 sky130_fd_sc_hd__bufbuf_16 hold488 (.A(net298),
    .X(net950));
 sky130_fd_sc_hd__bufbuf_16 hold489 (.A(\gpio_configure[14][9] ),
    .X(net951));
 sky130_fd_sc_hd__bufbuf_16 hold490 (.A(_0298_),
    .X(net952));
 sky130_fd_sc_hd__bufbuf_16 hold491 (.A(\mgmt_gpio_data[33] ),
    .X(net953));
 sky130_fd_sc_hd__bufbuf_16 hold492 (.A(_0429_),
    .X(net954));
 sky130_fd_sc_hd__bufbuf_16 hold493 (.A(\gpio_configure[15][7] ),
    .X(net955));
 sky130_fd_sc_hd__bufbuf_16 hold494 (.A(_0569_),
    .X(net956));
 sky130_fd_sc_hd__bufbuf_16 hold495 (.A(\gpio_configure[6][9] ),
    .X(net957));
 sky130_fd_sc_hd__bufbuf_16 hold496 (.A(_0185_),
    .X(net958));
 sky130_fd_sc_hd__bufbuf_16 hold497 (.A(\gpio_configure[33][9] ),
    .X(net959));
 sky130_fd_sc_hd__bufbuf_16 hold498 (.A(_0343_),
    .X(net960));
 sky130_fd_sc_hd__bufbuf_16 hold499 (.A(\gpio_configure[12][7] ),
    .X(net961));
 sky130_fd_sc_hd__bufbuf_16 hold500 (.A(_0545_),
    .X(net962));
 sky130_fd_sc_hd__bufbuf_16 hold501 (.A(\gpio_configure[22][9] ),
    .X(net963));
 sky130_fd_sc_hd__bufbuf_16 hold502 (.A(_0358_),
    .X(net964));
 sky130_fd_sc_hd__bufbuf_16 hold503 (.A(\gpio_configure[10][9] ),
    .X(net965));
 sky130_fd_sc_hd__bufbuf_16 hold504 (.A(_0213_),
    .X(net966));
 sky130_fd_sc_hd__bufbuf_16 hold505 (.A(\gpio_configure[24][7] ),
    .X(net967));
 sky130_fd_sc_hd__bufbuf_16 hold506 (.A(_0641_),
    .X(net968));
 sky130_fd_sc_hd__bufbuf_16 hold507 (.A(\gpio_configure[4][1] ),
    .X(net969));
 sky130_fd_sc_hd__bufbuf_16 hold508 (.A(\gpio_configure[15][1] ),
    .X(net970));
 sky130_fd_sc_hd__bufbuf_16 hold509 (.A(net231),
    .X(net971));
 sky130_fd_sc_hd__bufbuf_16 hold510 (.A(_0124_),
    .X(net972));
 sky130_fd_sc_hd__bufbuf_16 hold511 (.A(\gpio_configure[7][2] ),
    .X(net973));
 sky130_fd_sc_hd__bufbuf_16 hold512 (.A(_0500_),
    .X(net974));
 sky130_fd_sc_hd__bufbuf_16 hold513 (.A(\gpio_configure[8][9] ),
    .X(net975));
 sky130_fd_sc_hd__bufbuf_16 hold514 (.A(_0203_),
    .X(net976));
 sky130_fd_sc_hd__bufbuf_16 hold515 (.A(\gpio_configure[16][2] ),
    .X(net977));
 sky130_fd_sc_hd__bufbuf_16 hold516 (.A(_0572_),
    .X(net978));
 sky130_fd_sc_hd__bufbuf_16 hold517 (.A(\gpio_configure[27][9] ),
    .X(net979));
 sky130_fd_sc_hd__bufbuf_16 hold518 (.A(_0810_),
    .X(net980));
 sky130_fd_sc_hd__bufbuf_16 hold519 (.A(\gpio_configure[2][7] ),
    .X(net981));
 sky130_fd_sc_hd__bufbuf_16 hold520 (.A(_0465_),
    .X(net982));
 sky130_fd_sc_hd__bufbuf_16 hold521 (.A(\mgmt_gpio_data_buf[22] ),
    .X(net983));
 sky130_fd_sc_hd__bufbuf_16 hold522 (.A(_0295_),
    .X(net984));
 sky130_fd_sc_hd__bufbuf_16 hold523 (.A(\mgmt_gpio_data[6] ),
    .X(net985));
 sky130_fd_sc_hd__bufbuf_16 hold524 (.A(_0286_),
    .X(net986));
 sky130_fd_sc_hd__bufbuf_16 hold525 (.A(\mgmt_gpio_data_buf[10] ),
    .X(net987));
 sky130_fd_sc_hd__bufbuf_16 hold526 (.A(_0132_),
    .X(net988));
 sky130_fd_sc_hd__bufbuf_16 hold527 (.A(\gpio_configure[15][9] ),
    .X(net989));
 sky130_fd_sc_hd__bufbuf_16 hold528 (.A(_0303_),
    .X(net990));
 sky130_fd_sc_hd__bufbuf_16 hold529 (.A(\gpio_configure[6][7] ),
    .X(net991));
 sky130_fd_sc_hd__bufbuf_16 hold530 (.A(_0497_),
    .X(net992));
 sky130_fd_sc_hd__bufbuf_16 hold531 (.A(\gpio_configure[9][9] ),
    .X(net993));
 sky130_fd_sc_hd__bufbuf_16 hold532 (.A(_0208_),
    .X(net994));
 sky130_fd_sc_hd__bufbuf_16 hold533 (.A(\gpio_configure[37][2] ),
    .X(net995));
 sky130_fd_sc_hd__bufbuf_16 hold534 (.A(_0740_),
    .X(net996));
 sky130_fd_sc_hd__bufbuf_16 hold535 (.A(\gpio_configure[16][9] ),
    .X(net997));
 sky130_fd_sc_hd__bufbuf_16 hold536 (.A(_0233_),
    .X(net998));
 sky130_fd_sc_hd__bufbuf_16 hold537 (.A(net236),
    .X(net999));
 sky130_fd_sc_hd__bufbuf_16 hold538 (.A(_0128_),
    .X(net1000));
 sky130_fd_sc_hd__bufbuf_16 hold539 (.A(\gpio_configure[4][6] ),
    .X(net1001));
 sky130_fd_sc_hd__bufbuf_16 hold540 (.A(_0480_),
    .X(net1002));
 sky130_fd_sc_hd__bufbuf_16 hold541 (.A(net240),
    .X(net1003));
 sky130_fd_sc_hd__bufbuf_16 hold542 (.A(_0430_),
    .X(net1004));
 sky130_fd_sc_hd__bufbuf_16 hold543 (.A(\gpio_configure[32][2] ),
    .X(net1005));
 sky130_fd_sc_hd__bufbuf_16 hold544 (.A(_0700_),
    .X(net1006));
 sky130_fd_sc_hd__bufbuf_16 hold545 (.A(\gpio_configure[9][6] ),
    .X(net1007));
 sky130_fd_sc_hd__bufbuf_16 hold546 (.A(_0520_),
    .X(net1008));
 sky130_fd_sc_hd__bufbuf_16 hold547 (.A(\gpio_configure[32][1] ),
    .X(net1009));
 sky130_fd_sc_hd__bufbuf_16 hold548 (.A(net245),
    .X(net1010));
 sky130_fd_sc_hd__bufbuf_16 hold549 (.A(_0284_),
    .X(net1011));
 sky130_fd_sc_hd__bufbuf_16 hold550 (.A(\gpio_configure[14][2] ),
    .X(net1012));
 sky130_fd_sc_hd__bufbuf_16 hold551 (.A(_0556_),
    .X(net1013));
 sky130_fd_sc_hd__bufbuf_16 hold552 (.A(\gpio_configure[5][5] ),
    .X(net1014));
 sky130_fd_sc_hd__bufbuf_16 hold553 (.A(_0487_),
    .X(net1015));
 sky130_fd_sc_hd__bufbuf_16 hold554 (.A(\mgmt_gpio_data_buf[18] ),
    .X(net1016));
 sky130_fd_sc_hd__bufbuf_16 hold555 (.A(_0291_),
    .X(net1017));
 sky130_fd_sc_hd__bufbuf_16 hold556 (.A(\gpio_configure[2][1] ),
    .X(net1018));
 sky130_fd_sc_hd__bufbuf_16 hold557 (.A(\gpio_configure[7][9] ),
    .X(net1019));
 sky130_fd_sc_hd__bufbuf_16 hold558 (.A(_0198_),
    .X(net1020));
 sky130_fd_sc_hd__bufbuf_16 hold559 (.A(\gpio_configure[8][1] ),
    .X(net1021));
 sky130_fd_sc_hd__bufbuf_16 hold560 (.A(\gpio_configure[16][6] ),
    .X(net1022));
 sky130_fd_sc_hd__bufbuf_16 hold561 (.A(_0576_),
    .X(net1023));
 sky130_fd_sc_hd__bufbuf_16 hold562 (.A(\gpio_configure[12][5] ),
    .X(net1024));
 sky130_fd_sc_hd__bufbuf_16 hold563 (.A(_0543_),
    .X(net1025));
 sky130_fd_sc_hd__bufbuf_16 hold564 (.A(\gpio_configure[33][3] ),
    .X(net1026));
 sky130_fd_sc_hd__bufbuf_16 hold565 (.A(_0709_),
    .X(net1027));
 sky130_fd_sc_hd__bufbuf_16 hold566 (.A(\gpio_configure[35][9] ),
    .X(net1028));
 sky130_fd_sc_hd__bufbuf_16 hold567 (.A(_0323_),
    .X(net1029));
 sky130_fd_sc_hd__bufbuf_16 hold568 (.A(\gpio_configure[34][9] ),
    .X(net1030));
 sky130_fd_sc_hd__bufbuf_16 hold569 (.A(_0333_),
    .X(net1031));
 sky130_fd_sc_hd__bufbuf_16 hold570 (.A(\gpio_configure[18][5] ),
    .X(net1032));
 sky130_fd_sc_hd__bufbuf_16 hold571 (.A(_0591_),
    .X(net1033));
 sky130_fd_sc_hd__bufbuf_16 hold572 (.A(\gpio_configure[4][3] ),
    .X(net1034));
 sky130_fd_sc_hd__bufbuf_16 hold573 (.A(\gpio_configure[7][3] ),
    .X(net1035));
 sky130_fd_sc_hd__bufbuf_16 hold574 (.A(_0501_),
    .X(net1036));
 sky130_fd_sc_hd__bufbuf_16 hold575 (.A(serial_bb_data_1),
    .X(net1037));
 sky130_fd_sc_hd__bufbuf_16 hold576 (.A(_0418_),
    .X(net1038));
 sky130_fd_sc_hd__bufbuf_16 hold577 (.A(\gpio_configure[23][5] ),
    .X(net1039));
 sky130_fd_sc_hd__bufbuf_16 hold578 (.A(_0631_),
    .X(net1040));
 sky130_fd_sc_hd__bufbuf_16 hold579 (.A(\gpio_configure[13][5] ),
    .X(net1041));
 sky130_fd_sc_hd__bufbuf_16 hold580 (.A(_0551_),
    .X(net1042));
 sky130_fd_sc_hd__bufbuf_16 hold581 (.A(\gpio_configure[6][5] ),
    .X(net1043));
 sky130_fd_sc_hd__bufbuf_16 hold582 (.A(_0495_),
    .X(net1044));
 sky130_fd_sc_hd__bufbuf_16 hold583 (.A(\gpio_configure[5][3] ),
    .X(net1045));
 sky130_fd_sc_hd__bufbuf_16 hold584 (.A(\gpio_configure[32][3] ),
    .X(net1046));
 sky130_fd_sc_hd__bufbuf_16 hold585 (.A(\gpio_configure[7][6] ),
    .X(net1047));
 sky130_fd_sc_hd__bufbuf_16 hold586 (.A(_0504_),
    .X(net1048));
 sky130_fd_sc_hd__bufbuf_16 hold587 (.A(\gpio_configure[3][1] ),
    .X(net1049));
 sky130_fd_sc_hd__bufbuf_16 hold588 (.A(_0467_),
    .X(net1050));
 sky130_fd_sc_hd__bufbuf_16 hold589 (.A(\gpio_configure[8][6] ),
    .X(net1051));
 sky130_fd_sc_hd__bufbuf_16 hold590 (.A(_0512_),
    .X(net1052));
 sky130_fd_sc_hd__bufbuf_16 hold591 (.A(\gpio_configure[9][3] ),
    .X(net1053));
 sky130_fd_sc_hd__bufbuf_16 hold592 (.A(_0517_),
    .X(net1054));
 sky130_fd_sc_hd__bufbuf_16 hold593 (.A(\gpio_configure[10][7] ),
    .X(net1055));
 sky130_fd_sc_hd__bufbuf_16 hold594 (.A(_0529_),
    .X(net1056));
 sky130_fd_sc_hd__bufbuf_16 hold595 (.A(\gpio_configure[36][9] ),
    .X(net1057));
 sky130_fd_sc_hd__bufbuf_16 hold596 (.A(_0238_),
    .X(net1058));
 sky130_fd_sc_hd__bufbuf_16 hold597 (.A(\gpio_configure[25][6] ),
    .X(net1059));
 sky130_fd_sc_hd__bufbuf_16 hold598 (.A(_0648_),
    .X(net1060));
 sky130_fd_sc_hd__bufbuf_16 hold599 (.A(\gpio_configure[3][6] ),
    .X(net1061));
 sky130_fd_sc_hd__bufbuf_16 hold600 (.A(_0472_),
    .X(net1062));
 sky130_fd_sc_hd__bufbuf_16 hold601 (.A(\gpio_configure[34][3] ),
    .X(net1063));
 sky130_fd_sc_hd__bufbuf_16 hold602 (.A(_0717_),
    .X(net1064));
 sky130_fd_sc_hd__bufbuf_16 hold603 (.A(\gpio_configure[37][6] ),
    .X(net1065));
 sky130_fd_sc_hd__bufbuf_16 hold604 (.A(_0744_),
    .X(net1066));
 sky130_fd_sc_hd__bufbuf_16 hold605 (.A(net263),
    .X(net1067));
 sky130_fd_sc_hd__bufbuf_16 hold606 (.A(_0399_),
    .X(net1068));
 sky130_fd_sc_hd__bufbuf_16 hold607 (.A(\gpio_configure[29][9] ),
    .X(net1069));
 sky130_fd_sc_hd__bufbuf_16 hold608 (.A(_0253_),
    .X(net1070));
 sky130_fd_sc_hd__bufbuf_16 hold609 (.A(\gpio_configure[17][9] ),
    .X(net1071));
 sky130_fd_sc_hd__bufbuf_16 hold610 (.A(_0313_),
    .X(net1072));
 sky130_fd_sc_hd__bufbuf_16 hold611 (.A(\gpio_configure[37][9] ),
    .X(net1073));
 sky130_fd_sc_hd__bufbuf_16 hold612 (.A(_0308_),
    .X(net1074));
 sky130_fd_sc_hd__bufbuf_16 hold613 (.A(net279),
    .X(net1075));
 sky130_fd_sc_hd__bufbuf_16 hold614 (.A(net288),
    .X(net1076));
 sky130_fd_sc_hd__bufbuf_16 hold615 (.A(\gpio_configure[22][5] ),
    .X(net1077));
 sky130_fd_sc_hd__bufbuf_16 hold616 (.A(_0623_),
    .X(net1078));
 sky130_fd_sc_hd__bufbuf_16 hold617 (.A(\gpio_configure[16][3] ),
    .X(net1079));
 sky130_fd_sc_hd__bufbuf_16 hold618 (.A(_0573_),
    .X(net1080));
 sky130_fd_sc_hd__bufbuf_16 hold619 (.A(net296),
    .X(net1081));
 sky130_fd_sc_hd__bufbuf_16 hold620 (.A(\gpio_configure[1][4] ),
    .X(net1082));
 sky130_fd_sc_hd__bufbuf_16 hold621 (.A(_0454_),
    .X(net1083));
 sky130_fd_sc_hd__bufbuf_16 hold622 (.A(\gpio_configure[11][6] ),
    .X(net1084));
 sky130_fd_sc_hd__bufbuf_16 hold623 (.A(_0536_),
    .X(net1085));
 sky130_fd_sc_hd__bufbuf_16 hold624 (.A(\gpio_configure[10][6] ),
    .X(net1086));
 sky130_fd_sc_hd__bufbuf_16 hold625 (.A(_0528_),
    .X(net1087));
 sky130_fd_sc_hd__bufbuf_16 hold626 (.A(net280),
    .X(net1088));
 sky130_fd_sc_hd__bufbuf_16 hold627 (.A(\gpio_configure[5][1] ),
    .X(net1089));
 sky130_fd_sc_hd__bufbuf_16 hold628 (.A(\gpio_configure[18][6] ),
    .X(net1090));
 sky130_fd_sc_hd__bufbuf_16 hold629 (.A(\gpio_configure[18][3] ),
    .X(net1091));
 sky130_fd_sc_hd__bufbuf_16 hold630 (.A(\gpio_configure[14][3] ),
    .X(net1092));
 sky130_fd_sc_hd__bufbuf_16 hold631 (.A(_0557_),
    .X(net1093));
 sky130_fd_sc_hd__bufbuf_16 hold632 (.A(\gpio_configure[20][5] ),
    .X(net1094));
 sky130_fd_sc_hd__bufbuf_16 hold633 (.A(_0607_),
    .X(net1095));
 sky130_fd_sc_hd__bufbuf_16 hold634 (.A(\gpio_configure[30][5] ),
    .X(net1096));
 sky130_fd_sc_hd__bufbuf_16 hold635 (.A(_0687_),
    .X(net1097));
 sky130_fd_sc_hd__bufbuf_16 hold636 (.A(\gpio_configure[3][3] ),
    .X(net1098));
 sky130_fd_sc_hd__bufbuf_16 hold637 (.A(\gpio_configure[13][9] ),
    .X(net1099));
 sky130_fd_sc_hd__bufbuf_16 hold638 (.A(_0228_),
    .X(net1100));
 sky130_fd_sc_hd__bufbuf_16 hold639 (.A(\gpio_configure[31][6] ),
    .X(net1101));
 sky130_fd_sc_hd__bufbuf_16 hold640 (.A(_0696_),
    .X(net1102));
 sky130_fd_sc_hd__bufbuf_16 hold641 (.A(net1727),
    .X(net1103));
 sky130_fd_sc_hd__bufbuf_16 hold642 (.A(_0292_),
    .X(net1104));
 sky130_fd_sc_hd__bufbuf_16 hold643 (.A(\gpio_configure[23][6] ),
    .X(net1105));
 sky130_fd_sc_hd__bufbuf_16 hold644 (.A(_0632_),
    .X(net1106));
 sky130_fd_sc_hd__bufbuf_16 hold645 (.A(\gpio_configure[32][6] ),
    .X(net1107));
 sky130_fd_sc_hd__bufbuf_16 hold646 (.A(_0704_),
    .X(net1108));
 sky130_fd_sc_hd__bufbuf_16 hold647 (.A(\gpio_configure[29][6] ),
    .X(net1109));
 sky130_fd_sc_hd__bufbuf_16 hold648 (.A(_0680_),
    .X(net1110));
 sky130_fd_sc_hd__bufbuf_16 hold649 (.A(\gpio_configure[0][5] ),
    .X(net1111));
 sky130_fd_sc_hd__bufbuf_16 hold650 (.A(_0447_),
    .X(net1112));
 sky130_fd_sc_hd__bufbuf_16 hold651 (.A(\gpio_configure[34][6] ),
    .X(net1113));
 sky130_fd_sc_hd__bufbuf_16 hold652 (.A(_0720_),
    .X(net1114));
 sky130_fd_sc_hd__bufbuf_16 hold653 (.A(\gpio_configure[22][6] ),
    .X(net1115));
 sky130_fd_sc_hd__bufbuf_16 hold654 (.A(_0624_),
    .X(net1116));
 sky130_fd_sc_hd__bufbuf_16 hold655 (.A(\gpio_configure[24][5] ),
    .X(net1117));
 sky130_fd_sc_hd__bufbuf_16 hold656 (.A(_0639_),
    .X(net1118));
 sky130_fd_sc_hd__bufbuf_16 hold657 (.A(\gpio_configure[4][9] ),
    .X(net1119));
 sky130_fd_sc_hd__bufbuf_16 hold658 (.A(_0159_),
    .X(net1120));
 sky130_fd_sc_hd__bufbuf_16 hold659 (.A(\gpio_configure[5][6] ),
    .X(net1121));
 sky130_fd_sc_hd__bufbuf_16 hold660 (.A(_0488_),
    .X(net1122));
 sky130_fd_sc_hd__bufbuf_16 hold661 (.A(\gpio_configure[35][5] ),
    .X(net1123));
 sky130_fd_sc_hd__bufbuf_16 hold662 (.A(_0727_),
    .X(net1124));
 sky130_fd_sc_hd__bufbuf_16 hold663 (.A(\gpio_configure[8][3] ),
    .X(net1125));
 sky130_fd_sc_hd__bufbuf_16 hold664 (.A(_0509_),
    .X(net1126));
 sky130_fd_sc_hd__bufbuf_16 hold665 (.A(\gpio_configure[20][2] ),
    .X(net1127));
 sky130_fd_sc_hd__bufbuf_16 hold666 (.A(_0604_),
    .X(net1128));
 sky130_fd_sc_hd__bufbuf_16 hold667 (.A(\gpio_configure[29][5] ),
    .X(net1129));
 sky130_fd_sc_hd__bufbuf_16 hold668 (.A(_0679_),
    .X(net1130));
 sky130_fd_sc_hd__bufbuf_16 hold669 (.A(\gpio_configure[23][10] ),
    .X(net1131));
 sky130_fd_sc_hd__bufbuf_16 hold670 (.A(\gpio_configure[28][5] ),
    .X(net1132));
 sky130_fd_sc_hd__bufbuf_16 hold671 (.A(_0671_),
    .X(net1133));
 sky130_fd_sc_hd__bufbuf_16 hold672 (.A(serial_bb_data_2),
    .X(net1134));
 sky130_fd_sc_hd__bufbuf_16 hold673 (.A(_0419_),
    .X(net1135));
 sky130_fd_sc_hd__bufbuf_16 hold674 (.A(\gpio_configure[1][10] ),
    .X(net1136));
 sky130_fd_sc_hd__bufbuf_16 hold675 (.A(_0145_),
    .X(net1137));
 sky130_fd_sc_hd__bufbuf_16 hold676 (.A(\gpio_configure[17][2] ),
    .X(net1138));
 sky130_fd_sc_hd__bufbuf_16 hold677 (.A(_0580_),
    .X(net1139));
 sky130_fd_sc_hd__bufbuf_16 hold678 (.A(\gpio_configure[6][10] ),
    .X(net1140));
 sky130_fd_sc_hd__bufbuf_16 hold679 (.A(net289),
    .X(net1141));
 sky130_fd_sc_hd__bufbuf_16 hold680 (.A(net303),
    .X(net1142));
 sky130_fd_sc_hd__bufbuf_16 hold681 (.A(\gpio_configure[11][9] ),
    .X(net1143));
 sky130_fd_sc_hd__bufbuf_16 hold682 (.A(_0218_),
    .X(net1144));
 sky130_fd_sc_hd__bufbuf_16 hold683 (.A(\gpio_configure[23][2] ),
    .X(net1145));
 sky130_fd_sc_hd__bufbuf_16 hold684 (.A(_0628_),
    .X(net1146));
 sky130_fd_sc_hd__bufbuf_16 hold685 (.A(\gpio_configure[20][6] ),
    .X(net1147));
 sky130_fd_sc_hd__bufbuf_16 hold686 (.A(_0608_),
    .X(net1148));
 sky130_fd_sc_hd__bufbuf_16 hold687 (.A(\mgmt_gpio_data_buf[2] ),
    .X(net1149));
 sky130_fd_sc_hd__bufbuf_16 hold688 (.A(_0436_),
    .X(net1150));
 sky130_fd_sc_hd__bufbuf_16 hold689 (.A(\gpio_configure[25][10] ),
    .X(net1151));
 sky130_fd_sc_hd__bufbuf_16 hold690 (.A(\gpio_configure[14][10] ),
    .X(net1152));
 sky130_fd_sc_hd__bufbuf_16 hold691 (.A(\gpio_configure[21][5] ),
    .X(net1153));
 sky130_fd_sc_hd__bufbuf_16 hold692 (.A(_0615_),
    .X(net1154));
 sky130_fd_sc_hd__bufbuf_16 hold693 (.A(\gpio_configure[26][6] ),
    .X(net1155));
 sky130_fd_sc_hd__bufbuf_16 hold694 (.A(_0656_),
    .X(net1156));
 sky130_fd_sc_hd__bufbuf_16 hold695 (.A(\gpio_configure[12][1] ),
    .X(net1157));
 sky130_fd_sc_hd__bufbuf_16 hold696 (.A(\gpio_configure[19][6] ),
    .X(net1158));
 sky130_fd_sc_hd__bufbuf_16 hold697 (.A(_0600_),
    .X(net1159));
 sky130_fd_sc_hd__bufbuf_16 hold698 (.A(\gpio_configure[33][6] ),
    .X(net1160));
 sky130_fd_sc_hd__bufbuf_16 hold699 (.A(_0712_),
    .X(net1161));
 sky130_fd_sc_hd__bufbuf_16 hold700 (.A(\mgmt_gpio_data_buf[5] ),
    .X(net1162));
 sky130_fd_sc_hd__bufbuf_16 hold701 (.A(_0439_),
    .X(net1163));
 sky130_fd_sc_hd__bufbuf_16 hold702 (.A(\gpio_configure[24][2] ),
    .X(net1164));
 sky130_fd_sc_hd__bufbuf_16 hold703 (.A(_0636_),
    .X(net1165));
 sky130_fd_sc_hd__bufbuf_16 hold704 (.A(serial_bb_resetn),
    .X(net1166));
 sky130_fd_sc_hd__bufbuf_16 hold705 (.A(_0417_),
    .X(net1167));
 sky130_fd_sc_hd__bufbuf_16 hold706 (.A(\gpio_configure[0][6] ),
    .X(net1168));
 sky130_fd_sc_hd__bufbuf_16 hold707 (.A(_0448_),
    .X(net1169));
 sky130_fd_sc_hd__bufbuf_16 hold708 (.A(\gpio_configure[30][6] ),
    .X(net1170));
 sky130_fd_sc_hd__bufbuf_16 hold709 (.A(_0688_),
    .X(net1171));
 sky130_fd_sc_hd__bufbuf_16 hold710 (.A(\gpio_configure[11][5] ),
    .X(net1172));
 sky130_fd_sc_hd__bufbuf_16 hold711 (.A(_0535_),
    .X(net1173));
 sky130_fd_sc_hd__bufbuf_16 hold712 (.A(\gpio_configure[8][10] ),
    .X(net1174));
 sky130_fd_sc_hd__bufbuf_16 hold713 (.A(\gpio_configure[28][6] ),
    .X(net1175));
 sky130_fd_sc_hd__bufbuf_16 hold714 (.A(_0672_),
    .X(net1176));
 sky130_fd_sc_hd__bufbuf_16 hold715 (.A(\mgmt_gpio_data_buf[11] ),
    .X(net1177));
 sky130_fd_sc_hd__bufbuf_16 hold716 (.A(_0133_),
    .X(net1178));
 sky130_fd_sc_hd__bufbuf_16 hold717 (.A(\gpio_configure[19][2] ),
    .X(net1179));
 sky130_fd_sc_hd__bufbuf_16 hold718 (.A(_0596_),
    .X(net1180));
 sky130_fd_sc_hd__bufbuf_16 hold719 (.A(\mgmt_gpio_data[9] ),
    .X(net1181));
 sky130_fd_sc_hd__bufbuf_16 hold720 (.A(_0115_),
    .X(net1182));
 sky130_fd_sc_hd__bufbuf_16 hold721 (.A(\gpio_configure[24][6] ),
    .X(net1183));
 sky130_fd_sc_hd__bufbuf_16 hold722 (.A(_0640_),
    .X(net1184));
 sky130_fd_sc_hd__bufbuf_16 hold723 (.A(\gpio_configure[35][6] ),
    .X(net1185));
 sky130_fd_sc_hd__bufbuf_16 hold724 (.A(_0728_),
    .X(net1186));
 sky130_fd_sc_hd__bufbuf_16 hold725 (.A(clk1_output_dest),
    .X(net1187));
 sky130_fd_sc_hd__bufbuf_16 hold726 (.A(_0423_),
    .X(net1188));
 sky130_fd_sc_hd__bufbuf_16 hold727 (.A(net221),
    .X(net1189));
 sky130_fd_sc_hd__bufbuf_16 hold728 (.A(_0273_),
    .X(net1190));
 sky130_fd_sc_hd__bufbuf_16 hold729 (.A(\gpio_configure[21][6] ),
    .X(net1191));
 sky130_fd_sc_hd__bufbuf_16 hold730 (.A(_0616_),
    .X(net1192));
 sky130_fd_sc_hd__bufbuf_16 hold731 (.A(\gpio_configure[28][12] ),
    .X(net1193));
 sky130_fd_sc_hd__bufbuf_16 hold732 (.A(_0266_),
    .X(net1194));
 sky130_fd_sc_hd__bufbuf_16 hold733 (.A(\gpio_configure[30][12] ),
    .X(net1195));
 sky130_fd_sc_hd__bufbuf_16 hold734 (.A(_0378_),
    .X(net1196));
 sky130_fd_sc_hd__bufbuf_16 hold735 (.A(\gpio_configure[7][4] ),
    .X(net1197));
 sky130_fd_sc_hd__bufbuf_16 hold736 (.A(_0502_),
    .X(net1198));
 sky130_fd_sc_hd__bufbuf_16 hold737 (.A(\gpio_configure[6][6] ),
    .X(net1199));
 sky130_fd_sc_hd__bufbuf_16 hold738 (.A(_0496_),
    .X(net1200));
 sky130_fd_sc_hd__bufbuf_16 hold739 (.A(\gpio_configure[19][12] ),
    .X(net1201));
 sky130_fd_sc_hd__bufbuf_16 hold740 (.A(_0331_),
    .X(net1202));
 sky130_fd_sc_hd__bufbuf_16 hold741 (.A(\gpio_configure[6][1] ),
    .X(net1203));
 sky130_fd_sc_hd__bufbuf_16 hold742 (.A(\gpio_configure[15][11] ),
    .X(net1204));
 sky130_fd_sc_hd__bufbuf_16 hold743 (.A(_0305_),
    .X(net1205));
 sky130_fd_sc_hd__bufbuf_16 hold744 (.A(\gpio_configure[24][12] ),
    .X(net1206));
 sky130_fd_sc_hd__bufbuf_16 hold745 (.A(_0251_),
    .X(net1207));
 sky130_fd_sc_hd__bufbuf_16 hold746 (.A(\gpio_configure[14][6] ),
    .X(net1208));
 sky130_fd_sc_hd__bufbuf_16 hold747 (.A(_0560_),
    .X(net1209));
 sky130_fd_sc_hd__bufbuf_16 hold748 (.A(\gpio_configure[20][12] ),
    .X(net1210));
 sky130_fd_sc_hd__bufbuf_16 hold749 (.A(_0341_),
    .X(net1211));
 sky130_fd_sc_hd__bufbuf_16 hold750 (.A(\gpio_configure[27][12] ),
    .X(net1212));
 sky130_fd_sc_hd__bufbuf_16 hold751 (.A(_0813_),
    .X(net1213));
 sky130_fd_sc_hd__bufbuf_16 hold752 (.A(\gpio_configure[12][6] ),
    .X(net1214));
 sky130_fd_sc_hd__bufbuf_16 hold753 (.A(_0544_),
    .X(net1215));
 sky130_fd_sc_hd__bufbuf_16 hold754 (.A(\gpio_configure[31][12] ),
    .X(net1216));
 sky130_fd_sc_hd__bufbuf_16 hold755 (.A(_0246_),
    .X(net1217));
 sky130_fd_sc_hd__bufbuf_16 hold756 (.A(\gpio_configure[0][2] ),
    .X(net1218));
 sky130_fd_sc_hd__bufbuf_16 hold757 (.A(_0444_),
    .X(net1219));
 sky130_fd_sc_hd__bufbuf_16 hold758 (.A(net1344),
    .X(net1220));
 sky130_fd_sc_hd__bufbuf_16 hold759 (.A(net1346),
    .X(net1221));
 sky130_fd_sc_hd__bufbuf_16 hold760 (.A(_0130_),
    .X(net1222));
 sky130_fd_sc_hd__bufbuf_16 hold761 (.A(\gpio_configure[8][11] ),
    .X(net1223));
 sky130_fd_sc_hd__bufbuf_16 hold762 (.A(_0205_),
    .X(net1224));
 sky130_fd_sc_hd__bufbuf_16 hold763 (.A(\gpio_configure[21][12] ),
    .X(net1225));
 sky130_fd_sc_hd__bufbuf_16 hold764 (.A(_0351_),
    .X(net1226));
 sky130_fd_sc_hd__bufbuf_16 hold765 (.A(\gpio_configure[27][5] ),
    .X(net1227));
 sky130_fd_sc_hd__bufbuf_16 hold766 (.A(_0663_),
    .X(net1228));
 sky130_fd_sc_hd__bufbuf_16 hold767 (.A(\gpio_configure[2][6] ),
    .X(net1229));
 sky130_fd_sc_hd__bufbuf_16 hold768 (.A(_0464_),
    .X(net1230));
 sky130_fd_sc_hd__bufbuf_16 hold769 (.A(net295),
    .X(net1231));
 sky130_fd_sc_hd__bufbuf_16 hold770 (.A(net216),
    .X(net1232));
 sky130_fd_sc_hd__bufbuf_16 hold771 (.A(_0118_),
    .X(net1233));
 sky130_fd_sc_hd__bufbuf_16 hold772 (.A(\gpio_configure[14][11] ),
    .X(net1234));
 sky130_fd_sc_hd__bufbuf_16 hold773 (.A(_0300_),
    .X(net1235));
 sky130_fd_sc_hd__bufbuf_16 hold774 (.A(\gpio_configure[17][6] ),
    .X(net1236));
 sky130_fd_sc_hd__bufbuf_16 hold775 (.A(_0584_),
    .X(net1237));
 sky130_fd_sc_hd__bufbuf_16 hold776 (.A(\gpio_configure[22][2] ),
    .X(net1238));
 sky130_fd_sc_hd__bufbuf_16 hold777 (.A(_0620_),
    .X(net1239));
 sky130_fd_sc_hd__bufbuf_16 hold778 (.A(\gpio_configure[6][3] ),
    .X(net1240));
 sky130_fd_sc_hd__bufbuf_16 hold779 (.A(_0493_),
    .X(net1241));
 sky130_fd_sc_hd__bufbuf_16 hold780 (.A(\gpio_configure[6][11] ),
    .X(net1242));
 sky130_fd_sc_hd__bufbuf_16 hold781 (.A(_0187_),
    .X(net1243));
 sky130_fd_sc_hd__bufbuf_16 hold782 (.A(\gpio_configure[15][3] ),
    .X(net1244));
 sky130_fd_sc_hd__bufbuf_16 hold783 (.A(_0565_),
    .X(net1245));
 sky130_fd_sc_hd__bufbuf_16 hold784 (.A(\gpio_configure[15][2] ),
    .X(net1246));
 sky130_fd_sc_hd__bufbuf_16 hold785 (.A(_0564_),
    .X(net1247));
 sky130_fd_sc_hd__bufbuf_16 hold786 (.A(\gpio_configure[3][11] ),
    .X(net1248));
 sky130_fd_sc_hd__bufbuf_16 hold787 (.A(net262),
    .X(net1249));
 sky130_fd_sc_hd__bufbuf_16 hold788 (.A(\gpio_configure[18][12] ),
    .X(net1250));
 sky130_fd_sc_hd__bufbuf_16 hold789 (.A(_0321_),
    .X(net1251));
 sky130_fd_sc_hd__bufbuf_16 hold790 (.A(\gpio_configure[22][12] ),
    .X(net1252));
 sky130_fd_sc_hd__bufbuf_16 hold791 (.A(_0361_),
    .X(net1253));
 sky130_fd_sc_hd__bufbuf_16 hold792 (.A(\gpio_configure[0][11] ),
    .X(net1254));
 sky130_fd_sc_hd__bufbuf_16 hold793 (.A(\gpio_configure[10][3] ),
    .X(net1255));
 sky130_fd_sc_hd__bufbuf_16 hold794 (.A(\gpio_configure[11][12] ),
    .X(net1256));
 sky130_fd_sc_hd__bufbuf_16 hold795 (.A(_0221_),
    .X(net1257));
 sky130_fd_sc_hd__bufbuf_16 hold796 (.A(\gpio_configure[12][3] ),
    .X(net1258));
 sky130_fd_sc_hd__bufbuf_16 hold797 (.A(_0541_),
    .X(net1259));
 sky130_fd_sc_hd__bufbuf_16 hold798 (.A(\gpio_configure[21][11] ),
    .X(net1260));
 sky130_fd_sc_hd__bufbuf_16 hold799 (.A(_0350_),
    .X(net1261));
 sky130_fd_sc_hd__bufbuf_16 hold800 (.A(\gpio_configure[22][11] ),
    .X(net1262));
 sky130_fd_sc_hd__bufbuf_16 hold801 (.A(_0360_),
    .X(net1263));
 sky130_fd_sc_hd__bufbuf_16 hold802 (.A(\mgmt_gpio_data[13] ),
    .X(net1264));
 sky130_fd_sc_hd__bufbuf_16 hold803 (.A(_0119_),
    .X(net1265));
 sky130_fd_sc_hd__bufbuf_16 hold804 (.A(\gpio_configure[25][11] ),
    .X(net1266));
 sky130_fd_sc_hd__bufbuf_16 hold805 (.A(_0260_),
    .X(net1267));
 sky130_fd_sc_hd__bufbuf_16 hold806 (.A(\gpio_configure[9][12] ),
    .X(net1268));
 sky130_fd_sc_hd__bufbuf_16 hold807 (.A(_0211_),
    .X(net1269));
 sky130_fd_sc_hd__bufbuf_16 hold808 (.A(\gpio_configure[12][11] ),
    .X(net1270));
 sky130_fd_sc_hd__bufbuf_16 hold809 (.A(_0225_),
    .X(net1271));
 sky130_fd_sc_hd__bufbuf_16 hold810 (.A(\hkspi.wrstb ),
    .X(net1272));
 sky130_fd_sc_hd__bufbuf_16 hold811 (.A(net559),
    .X(net1273));
 sky130_fd_sc_hd__bufbuf_16 hold812 (.A(_1465_),
    .X(net1274));
 sky130_fd_sc_hd__bufbuf_16 hold813 (.A(net677),
    .X(net1275));
 sky130_fd_sc_hd__bufbuf_16 hold814 (.A(_0293_),
    .X(net1276));
 sky130_fd_sc_hd__bufbuf_16 hold815 (.A(\gpio_configure[16][12] ),
    .X(net1277));
 sky130_fd_sc_hd__bufbuf_16 hold816 (.A(_0236_),
    .X(net1278));
 sky130_fd_sc_hd__bufbuf_16 hold817 (.A(\gpio_configure[13][11] ),
    .X(net1279));
 sky130_fd_sc_hd__bufbuf_16 hold818 (.A(_0230_),
    .X(net1280));
 sky130_fd_sc_hd__bufbuf_16 hold819 (.A(\gpio_configure[32][4] ),
    .X(net1281));
 sky130_fd_sc_hd__bufbuf_16 hold820 (.A(_0702_),
    .X(net1282));
 sky130_fd_sc_hd__bufbuf_16 hold821 (.A(\gpio_configure[26][12] ),
    .X(net1283));
 sky130_fd_sc_hd__bufbuf_16 hold822 (.A(_0271_),
    .X(net1284));
 sky130_fd_sc_hd__bufbuf_16 hold823 (.A(net270),
    .X(net1285));
 sky130_fd_sc_hd__bufbuf_16 hold824 (.A(_0393_),
    .X(net1286));
 sky130_fd_sc_hd__bufbuf_16 hold825 (.A(\gpio_configure[33][2] ),
    .X(net1287));
 sky130_fd_sc_hd__bufbuf_16 hold826 (.A(_0708_),
    .X(net1288));
 sky130_fd_sc_hd__bufbuf_16 hold827 (.A(\gpio_configure[5][4] ),
    .X(net1289));
 sky130_fd_sc_hd__bufbuf_16 hold828 (.A(_0486_),
    .X(net1290));
 sky130_fd_sc_hd__bufbuf_16 hold829 (.A(\gpio_configure[7][11] ),
    .X(net1291));
 sky130_fd_sc_hd__bufbuf_16 hold830 (.A(_0200_),
    .X(net1292));
 sky130_fd_sc_hd__bufbuf_16 hold831 (.A(\gpio_configure[33][12] ),
    .X(net1293));
 sky130_fd_sc_hd__bufbuf_16 hold832 (.A(_0346_),
    .X(net1294));
 sky130_fd_sc_hd__bufbuf_16 hold833 (.A(\gpio_configure[33][4] ),
    .X(net1295));
 sky130_fd_sc_hd__bufbuf_16 hold834 (.A(_0710_),
    .X(net1296));
 sky130_fd_sc_hd__bufbuf_16 hold835 (.A(\gpio_configure[34][11] ),
    .X(net1297));
 sky130_fd_sc_hd__bufbuf_16 hold836 (.A(_0335_),
    .X(net1298));
 sky130_fd_sc_hd__bufbuf_16 hold837 (.A(\gpio_configure[8][4] ),
    .X(net1299));
 sky130_fd_sc_hd__bufbuf_16 hold838 (.A(_0510_),
    .X(net1300));
 sky130_fd_sc_hd__bufbuf_16 hold839 (.A(\gpio_configure[36][4] ),
    .X(net1301));
 sky130_fd_sc_hd__bufbuf_16 hold840 (.A(_0734_),
    .X(net1302));
 sky130_fd_sc_hd__bufbuf_16 hold841 (.A(\gpio_configure[37][11] ),
    .X(net1303));
 sky130_fd_sc_hd__bufbuf_16 hold842 (.A(_0310_),
    .X(net1304));
 sky130_fd_sc_hd__bufbuf_16 hold843 (.A(\gpio_configure[3][4] ),
    .X(net1305));
 sky130_fd_sc_hd__bufbuf_16 hold844 (.A(_0470_),
    .X(net1306));
 sky130_fd_sc_hd__bufbuf_16 hold845 (.A(\gpio_configure[10][4] ),
    .X(net1307));
 sky130_fd_sc_hd__bufbuf_16 hold846 (.A(_0526_),
    .X(net1308));
 sky130_fd_sc_hd__bufbuf_16 hold847 (.A(net248),
    .X(net1309));
 sky130_fd_sc_hd__bufbuf_16 hold848 (.A(_0287_),
    .X(net1310));
 sky130_fd_sc_hd__bufbuf_16 hold849 (.A(\gpio_configure[12][4] ),
    .X(net1311));
 sky130_fd_sc_hd__bufbuf_16 hold850 (.A(_0542_),
    .X(net1312));
 sky130_fd_sc_hd__bufbuf_16 hold851 (.A(\gpio_configure[4][4] ),
    .X(net1313));
 sky130_fd_sc_hd__bufbuf_16 hold852 (.A(_0478_),
    .X(net1314));
 sky130_fd_sc_hd__bufbuf_16 hold853 (.A(\gpio_configure[25][4] ),
    .X(net1315));
 sky130_fd_sc_hd__bufbuf_16 hold854 (.A(_0646_),
    .X(net1316));
 sky130_fd_sc_hd__bufbuf_16 hold855 (.A(\gpio_configure[2][4] ),
    .X(net1317));
 sky130_fd_sc_hd__bufbuf_16 hold856 (.A(_0462_),
    .X(net1318));
 sky130_fd_sc_hd__bufbuf_16 hold857 (.A(\gpio_configure[22][4] ),
    .X(net1319));
 sky130_fd_sc_hd__bufbuf_16 hold858 (.A(_0622_),
    .X(net1320));
 sky130_fd_sc_hd__bufbuf_16 hold859 (.A(\gpio_configure[31][2] ),
    .X(net1321));
 sky130_fd_sc_hd__bufbuf_16 hold860 (.A(_0692_),
    .X(net1322));
 sky130_fd_sc_hd__bufbuf_16 hold861 (.A(\gpio_configure[29][11] ),
    .X(net1323));
 sky130_fd_sc_hd__bufbuf_16 hold862 (.A(_0255_),
    .X(net1324));
 sky130_fd_sc_hd__bufbuf_16 hold863 (.A(\gpio_configure[37][4] ),
    .X(net1325));
 sky130_fd_sc_hd__bufbuf_16 hold864 (.A(_0742_),
    .X(net1326));
 sky130_fd_sc_hd__bufbuf_16 hold865 (.A(\gpio_configure[35][11] ),
    .X(net1327));
 sky130_fd_sc_hd__bufbuf_16 hold866 (.A(_0325_),
    .X(net1328));
 sky130_fd_sc_hd__bufbuf_16 hold867 (.A(\gpio_configure[15][10] ),
    .X(net1329));
 sky130_fd_sc_hd__bufbuf_16 hold868 (.A(\gpio_configure[35][4] ),
    .X(net1330));
 sky130_fd_sc_hd__bufbuf_16 hold869 (.A(_0726_),
    .X(net1331));
 sky130_fd_sc_hd__bufbuf_16 hold870 (.A(\gpio_configure[17][11] ),
    .X(net1332));
 sky130_fd_sc_hd__bufbuf_16 hold871 (.A(_0315_),
    .X(net1333));
 sky130_fd_sc_hd__bufbuf_16 hold872 (.A(\gpio_configure[17][12] ),
    .X(net1334));
 sky130_fd_sc_hd__bufbuf_16 hold873 (.A(_0316_),
    .X(net1335));
 sky130_fd_sc_hd__bufbuf_16 hold874 (.A(net227),
    .X(net1336));
 sky130_fd_sc_hd__bufbuf_16 hold875 (.A(_0278_),
    .X(net1337));
 sky130_fd_sc_hd__bufbuf_16 hold876 (.A(\mgmt_gpio_data[10] ),
    .X(net1338));
 sky130_fd_sc_hd__bufbuf_16 hold877 (.A(_0116_),
    .X(net1339));
 sky130_fd_sc_hd__bufbuf_16 hold878 (.A(\gpio_configure[4][12] ),
    .X(net1340));
 sky130_fd_sc_hd__bufbuf_16 hold879 (.A(_0162_),
    .X(net1341));
 sky130_fd_sc_hd__bufbuf_16 hold880 (.A(\mgmt_gpio_data[36] ),
    .X(net1342));
 sky130_fd_sc_hd__bufbuf_16 hold881 (.A(_0432_),
    .X(net1343));
 sky130_fd_sc_hd__bufbuf_16 hold882 (.A(\wbbd_data[0] ),
    .X(net1344));
 sky130_fd_sc_hd__bufbuf_16 hold883 (.A(net1220),
    .X(net1345));
 sky130_fd_sc_hd__bufbuf_16 hold884 (.A(_1467_),
    .X(net1346));
 sky130_fd_sc_hd__bufbuf_16 hold885 (.A(net1221),
    .X(net1347));
 sky130_fd_sc_hd__bufbuf_16 hold886 (.A(_0546_),
    .X(net1348));
 sky130_fd_sc_hd__bufbuf_16 hold887 (.A(net222),
    .X(net1349));
 sky130_fd_sc_hd__bufbuf_16 hold888 (.A(_0274_),
    .X(net1350));
 sky130_fd_sc_hd__bufbuf_16 hold889 (.A(\mgmt_gpio_data[14] ),
    .X(net1351));
 sky130_fd_sc_hd__bufbuf_16 hold890 (.A(_0120_),
    .X(net1352));
 sky130_fd_sc_hd__bufbuf_16 hold891 (.A(\gpio_configure[1][9] ),
    .X(net1353));
 sky130_fd_sc_hd__bufbuf_16 hold892 (.A(_0144_),
    .X(net1354));
 sky130_fd_sc_hd__bufbuf_16 hold893 (.A(\gpio_configure[2][9] ),
    .X(net1355));
 sky130_fd_sc_hd__bufbuf_16 hold894 (.A(_0149_),
    .X(net1356));
 sky130_fd_sc_hd__bufbuf_16 hold895 (.A(\gpio_configure[31][9] ),
    .X(net1357));
 sky130_fd_sc_hd__bufbuf_16 hold896 (.A(_0243_),
    .X(net1358));
 sky130_fd_sc_hd__bufbuf_16 hold897 (.A(\gpio_configure[28][9] ),
    .X(net1359));
 sky130_fd_sc_hd__bufbuf_16 hold898 (.A(_0263_),
    .X(net1360));
 sky130_fd_sc_hd__bufbuf_16 hold899 (.A(\gpio_configure[0][9] ),
    .X(net1361));
 sky130_fd_sc_hd__bufbuf_16 hold900 (.A(_0139_),
    .X(net1362));
 sky130_fd_sc_hd__bufbuf_16 hold901 (.A(\gpio_configure[30][9] ),
    .X(net1363));
 sky130_fd_sc_hd__bufbuf_16 hold902 (.A(_0375_),
    .X(net1364));
 sky130_fd_sc_hd__bufbuf_16 hold903 (.A(net285),
    .X(net1365));
 sky130_fd_sc_hd__bufbuf_16 hold904 (.A(_0403_),
    .X(net1366));
 sky130_fd_sc_hd__bufbuf_16 hold905 (.A(\gpio_configure[35][8] ),
    .X(net1367));
 sky130_fd_sc_hd__bufbuf_16 hold906 (.A(_0322_),
    .X(net1368));
 sky130_fd_sc_hd__bufbuf_16 hold907 (.A(\gpio_configure[20][9] ),
    .X(net1369));
 sky130_fd_sc_hd__bufbuf_16 hold908 (.A(_0338_),
    .X(net1370));
 sky130_fd_sc_hd__bufbuf_16 hold909 (.A(net286),
    .X(net1371));
 sky130_fd_sc_hd__bufbuf_16 hold910 (.A(\gpio_configure[24][9] ),
    .X(net1372));
 sky130_fd_sc_hd__bufbuf_16 hold911 (.A(_0248_),
    .X(net1373));
 sky130_fd_sc_hd__bufbuf_16 hold912 (.A(\mgmt_gpio_data_buf[1] ),
    .X(net1374));
 sky130_fd_sc_hd__bufbuf_16 hold913 (.A(_0435_),
    .X(net1375));
 sky130_fd_sc_hd__bufbuf_16 hold914 (.A(\gpio_configure[32][9] ),
    .X(net1376));
 sky130_fd_sc_hd__bufbuf_16 hold915 (.A(_0353_),
    .X(net1377));
 sky130_fd_sc_hd__bufbuf_16 hold916 (.A(net223),
    .X(net1378));
 sky130_fd_sc_hd__bufbuf_16 hold917 (.A(_0275_),
    .X(net1379));
 sky130_fd_sc_hd__bufbuf_16 hold918 (.A(\gpio_configure[15][0] ),
    .X(net1380));
 sky130_fd_sc_hd__bufbuf_16 hold919 (.A(net273),
    .X(net1381));
 sky130_fd_sc_hd__bufbuf_16 hold920 (.A(net300),
    .X(net1382));
 sky130_fd_sc_hd__bufbuf_16 hold921 (.A(net235),
    .X(net1383));
 sky130_fd_sc_hd__bufbuf_16 hold922 (.A(_0282_),
    .X(net1384));
 sky130_fd_sc_hd__bufbuf_16 hold923 (.A(\gpio_configure[35][0] ),
    .X(net1385));
 sky130_fd_sc_hd__bufbuf_16 hold924 (.A(\gpio_configure[25][0] ),
    .X(net1386));
 sky130_fd_sc_hd__bufbuf_16 hold925 (.A(\gpio_configure[35][12] ),
    .X(net1387));
 sky130_fd_sc_hd__bufbuf_16 hold926 (.A(_0326_),
    .X(net1388));
 sky130_fd_sc_hd__bufbuf_16 hold927 (.A(net265),
    .X(net1389));
 sky130_fd_sc_hd__bufbuf_16 hold928 (.A(\gpio_configure[23][9] ),
    .X(net1390));
 sky130_fd_sc_hd__bufbuf_16 hold929 (.A(_0363_),
    .X(net1391));
 sky130_fd_sc_hd__bufbuf_16 hold930 (.A(net246),
    .X(net1392));
 sky130_fd_sc_hd__bufbuf_16 hold931 (.A(_0285_),
    .X(net1393));
 sky130_fd_sc_hd__bufbuf_16 hold932 (.A(net267),
    .X(net1394));
 sky130_fd_sc_hd__bufbuf_16 hold933 (.A(_0390_),
    .X(net1395));
 sky130_fd_sc_hd__bufbuf_16 hold934 (.A(\gpio_configure[18][9] ),
    .X(net1396));
 sky130_fd_sc_hd__bufbuf_16 hold935 (.A(_0318_),
    .X(net1397));
 sky130_fd_sc_hd__bufbuf_16 hold936 (.A(irq_2_inputsrc),
    .X(net1398));
 sky130_fd_sc_hd__bufbuf_16 hold937 (.A(_0427_),
    .X(net1399));
 sky130_fd_sc_hd__bufbuf_16 hold938 (.A(\gpio_configure[25][2] ),
    .X(net1400));
 sky130_fd_sc_hd__bufbuf_16 hold939 (.A(_0644_),
    .X(net1401));
 sky130_fd_sc_hd__bufbuf_16 hold940 (.A(\gpio_configure[26][9] ),
    .X(net1402));
 sky130_fd_sc_hd__bufbuf_16 hold941 (.A(_0268_),
    .X(net1403));
 sky130_fd_sc_hd__bufbuf_16 hold942 (.A(\gpio_configure[17][10] ),
    .X(net1404));
 sky130_fd_sc_hd__bufbuf_16 hold943 (.A(net215),
    .X(net1405));
 sky130_fd_sc_hd__bufbuf_16 hold944 (.A(_0117_),
    .X(net1406));
 sky130_fd_sc_hd__bufbuf_16 hold945 (.A(\gpio_configure[4][2] ),
    .X(net1407));
 sky130_fd_sc_hd__bufbuf_16 hold946 (.A(_0476_),
    .X(net1408));
 sky130_fd_sc_hd__bufbuf_16 hold947 (.A(\gpio_configure[35][10] ),
    .X(net1409));
 sky130_fd_sc_hd__bufbuf_16 hold948 (.A(\mgmt_gpio_data[8] ),
    .X(net1410));
 sky130_fd_sc_hd__bufbuf_16 hold949 (.A(_0114_),
    .X(net1411));
 sky130_fd_sc_hd__bufbuf_16 hold950 (.A(\gpio_configure[13][10] ),
    .X(net1412));
 sky130_fd_sc_hd__bufbuf_16 hold951 (.A(_0229_),
    .X(net1413));
 sky130_fd_sc_hd__bufbuf_16 hold952 (.A(\gpio_configure[7][10] ),
    .X(net1414));
 sky130_fd_sc_hd__bufbuf_16 hold953 (.A(net220),
    .X(net1415));
 sky130_fd_sc_hd__bufbuf_16 hold954 (.A(_0272_),
    .X(net1416));
 sky130_fd_sc_hd__bufbuf_16 hold955 (.A(\gpio_configure[10][10] ),
    .X(net1417));
 sky130_fd_sc_hd__bufbuf_16 hold956 (.A(\mgmt_gpio_data_buf[16] ),
    .X(net1418));
 sky130_fd_sc_hd__bufbuf_16 hold957 (.A(_0289_),
    .X(net1419));
 sky130_fd_sc_hd__bufbuf_16 hold958 (.A(\gpio_configure[3][10] ),
    .X(net1420));
 sky130_fd_sc_hd__bufbuf_16 hold959 (.A(_0155_),
    .X(net1421));
 sky130_fd_sc_hd__bufbuf_16 hold960 (.A(\gpio_configure[8][0] ),
    .X(net1422));
 sky130_fd_sc_hd__bufbuf_16 hold961 (.A(\gpio_configure[34][0] ),
    .X(net1423));
 sky130_fd_sc_hd__bufbuf_16 hold962 (.A(\gpio_configure[9][0] ),
    .X(net1424));
 sky130_fd_sc_hd__bufbuf_16 hold963 (.A(\mgmt_gpio_data_buf[0] ),
    .X(net1425));
 sky130_fd_sc_hd__bufbuf_16 hold964 (.A(_0434_),
    .X(net1426));
 sky130_fd_sc_hd__bufbuf_16 hold965 (.A(\gpio_configure[5][0] ),
    .X(net1427));
 sky130_fd_sc_hd__bufbuf_16 hold966 (.A(\gpio_configure[31][11] ),
    .X(net1428));
 sky130_fd_sc_hd__bufbuf_16 hold967 (.A(_0245_),
    .X(net1429));
 sky130_fd_sc_hd__bufbuf_16 hold968 (.A(\gpio_configure[36][10] ),
    .X(net1430));
 sky130_fd_sc_hd__bufbuf_16 hold969 (.A(_0239_),
    .X(net1431));
 sky130_fd_sc_hd__bufbuf_16 hold970 (.A(\gpio_configure[30][11] ),
    .X(net1432));
 sky130_fd_sc_hd__bufbuf_16 hold971 (.A(_0377_),
    .X(net1433));
 sky130_fd_sc_hd__bufbuf_16 hold972 (.A(\gpio_configure[28][11] ),
    .X(net1434));
 sky130_fd_sc_hd__bufbuf_16 hold973 (.A(_0265_),
    .X(net1435));
 sky130_fd_sc_hd__bufbuf_16 hold974 (.A(\gpio_configure[2][0] ),
    .X(net1436));
 sky130_fd_sc_hd__bufbuf_16 hold975 (.A(\gpio_configure[16][0] ),
    .X(net1437));
 sky130_fd_sc_hd__bufbuf_16 hold976 (.A(\gpio_configure[32][0] ),
    .X(net1438));
 sky130_fd_sc_hd__bufbuf_16 hold977 (.A(\gpio_configure[27][11] ),
    .X(net1439));
 sky130_fd_sc_hd__bufbuf_16 hold978 (.A(_0812_),
    .X(net1440));
 sky130_fd_sc_hd__bufbuf_16 hold979 (.A(\gpio_configure[12][10] ),
    .X(net1441));
 sky130_fd_sc_hd__bufbuf_16 hold980 (.A(net261),
    .X(net1442));
 sky130_fd_sc_hd__bufbuf_16 hold981 (.A(_0397_),
    .X(net1443));
 sky130_fd_sc_hd__bufbuf_16 hold982 (.A(net229),
    .X(net1444));
 sky130_fd_sc_hd__bufbuf_16 hold983 (.A(_0122_),
    .X(net1445));
 sky130_fd_sc_hd__bufbuf_16 hold984 (.A(\gpio_configure[33][0] ),
    .X(net1446));
 sky130_fd_sc_hd__bufbuf_16 hold985 (.A(\gpio_configure[1][0] ),
    .X(net1447));
 sky130_fd_sc_hd__bufbuf_16 hold986 (.A(\gpio_configure[5][10] ),
    .X(net1448));
 sky130_fd_sc_hd__bufbuf_16 hold987 (.A(_0173_),
    .X(net1449));
 sky130_fd_sc_hd__bufbuf_16 hold988 (.A(\gpio_configure[36][0] ),
    .X(net1450));
 sky130_fd_sc_hd__bufbuf_16 hold989 (.A(\gpio_configure[1][11] ),
    .X(net1451));
 sky130_fd_sc_hd__bufbuf_16 hold990 (.A(\gpio_configure[19][11] ),
    .X(net1452));
 sky130_fd_sc_hd__bufbuf_16 hold991 (.A(_0330_),
    .X(net1453));
 sky130_fd_sc_hd__bufbuf_16 hold992 (.A(\gpio_configure[24][10] ),
    .X(net1454));
 sky130_fd_sc_hd__bufbuf_16 hold993 (.A(\gpio_configure[20][11] ),
    .X(net1455));
 sky130_fd_sc_hd__bufbuf_16 hold994 (.A(_0340_),
    .X(net1456));
 sky130_fd_sc_hd__bufbuf_16 hold995 (.A(\gpio_configure[27][10] ),
    .X(net1457));
 sky130_fd_sc_hd__bufbuf_16 hold996 (.A(\gpio_configure[30][10] ),
    .X(net1458));
 sky130_fd_sc_hd__bufbuf_16 hold997 (.A(net276),
    .X(net1459));
 sky130_fd_sc_hd__bufbuf_16 hold998 (.A(\gpio_configure[0][10] ),
    .X(net1460));
 sky130_fd_sc_hd__bufbuf_16 hold999 (.A(_0140_),
    .X(net1461));
 sky130_fd_sc_hd__bufbuf_16 hold1000 (.A(\gpio_configure[23][11] ),
    .X(net1462));
 sky130_fd_sc_hd__bufbuf_16 hold1001 (.A(_0365_),
    .X(net1463));
 sky130_fd_sc_hd__bufbuf_16 hold1002 (.A(\gpio_configure[28][10] ),
    .X(net1464));
 sky130_fd_sc_hd__bufbuf_16 hold1003 (.A(\gpio_configure[37][0] ),
    .X(net1465));
 sky130_fd_sc_hd__bufbuf_16 hold1004 (.A(\gpio_configure[19][10] ),
    .X(net1466));
 sky130_fd_sc_hd__bufbuf_16 hold1005 (.A(net277),
    .X(net1467));
 sky130_fd_sc_hd__bufbuf_16 hold1006 (.A(\gpio_configure[2][11] ),
    .X(net1468));
 sky130_fd_sc_hd__bufbuf_16 hold1007 (.A(_0151_),
    .X(net1469));
 sky130_fd_sc_hd__bufbuf_16 hold1008 (.A(\gpio_configure[20][10] ),
    .X(net1470));
 sky130_fd_sc_hd__bufbuf_16 hold1009 (.A(\gpio_configure[31][10] ),
    .X(net1471));
 sky130_fd_sc_hd__bufbuf_16 hold1010 (.A(\mgmt_gpio_data[35] ),
    .X(net1472));
 sky130_fd_sc_hd__bufbuf_16 hold1011 (.A(_0431_),
    .X(net1473));
 sky130_fd_sc_hd__bufbuf_16 hold1012 (.A(\gpio_configure[32][11] ),
    .X(net1474));
 sky130_fd_sc_hd__bufbuf_16 hold1013 (.A(_0355_),
    .X(net1475));
 sky130_fd_sc_hd__bufbuf_16 hold1014 (.A(net269),
    .X(net1476));
 sky130_fd_sc_hd__bufbuf_16 hold1015 (.A(_0392_),
    .X(net1477));
 sky130_fd_sc_hd__bufbuf_16 hold1016 (.A(net294),
    .X(net1478));
 sky130_fd_sc_hd__bufbuf_16 hold1017 (.A(\gpio_configure[18][11] ),
    .X(net1479));
 sky130_fd_sc_hd__bufbuf_16 hold1018 (.A(_0320_),
    .X(net1480));
 sky130_fd_sc_hd__bufbuf_16 hold1019 (.A(\gpio_configure[24][11] ),
    .X(net1481));
 sky130_fd_sc_hd__bufbuf_16 hold1020 (.A(_0250_),
    .X(net1482));
 sky130_fd_sc_hd__bufbuf_16 hold1021 (.A(\gpio_configure[14][0] ),
    .X(net1483));
 sky130_fd_sc_hd__bufbuf_16 hold1022 (.A(\gpio_configure[32][12] ),
    .X(net1484));
 sky130_fd_sc_hd__bufbuf_16 hold1023 (.A(_0356_),
    .X(net1485));
 sky130_fd_sc_hd__bufbuf_16 hold1024 (.A(\gpio_configure[12][0] ),
    .X(net1486));
 sky130_fd_sc_hd__bufbuf_16 hold1025 (.A(\gpio_configure[7][0] ),
    .X(net1487));
 sky130_fd_sc_hd__bufbuf_16 hold1026 (.A(net274),
    .X(net1488));
 sky130_fd_sc_hd__bufbuf_16 hold1027 (.A(_0396_),
    .X(net1489));
 sky130_fd_sc_hd__bufbuf_16 hold1028 (.A(\gpio_configure[32][10] ),
    .X(net1490));
 sky130_fd_sc_hd__bufbuf_16 hold1029 (.A(\gpio_configure[4][0] ),
    .X(net1491));
 sky130_fd_sc_hd__bufbuf_16 hold1030 (.A(\gpio_configure[8][12] ),
    .X(net1492));
 sky130_fd_sc_hd__bufbuf_16 hold1031 (.A(_0206_),
    .X(net1493));
 sky130_fd_sc_hd__bufbuf_16 hold1032 (.A(\gpio_configure[26][10] ),
    .X(net1494));
 sky130_fd_sc_hd__bufbuf_16 hold1033 (.A(\gpio_configure[26][11] ),
    .X(net1495));
 sky130_fd_sc_hd__bufbuf_16 hold1034 (.A(_0270_),
    .X(net1496));
 sky130_fd_sc_hd__bufbuf_16 hold1035 (.A(\gpio_configure[18][10] ),
    .X(net1497));
 sky130_fd_sc_hd__bufbuf_16 hold1036 (.A(\gpio_configure[15][12] ),
    .X(net1498));
 sky130_fd_sc_hd__bufbuf_16 hold1037 (.A(_0306_),
    .X(net1499));
 sky130_fd_sc_hd__bufbuf_16 hold1038 (.A(net293),
    .X(net1500));
 sky130_fd_sc_hd__bufbuf_16 hold1039 (.A(\gpio_configure[6][12] ),
    .X(net1501));
 sky130_fd_sc_hd__bufbuf_16 hold1040 (.A(_0188_),
    .X(net1502));
 sky130_fd_sc_hd__bufbuf_16 hold1041 (.A(net284),
    .X(net1503));
 sky130_fd_sc_hd__bufbuf_16 hold1042 (.A(\gpio_configure[10][0] ),
    .X(net1504));
 sky130_fd_sc_hd__bufbuf_16 hold1043 (.A(\gpio_configure[3][12] ),
    .X(net1505));
 sky130_fd_sc_hd__bufbuf_16 hold1044 (.A(_0157_),
    .X(net1506));
 sky130_fd_sc_hd__bufbuf_16 hold1045 (.A(\gpio_configure[21][10] ),
    .X(net1507));
 sky130_fd_sc_hd__bufbuf_16 hold1046 (.A(\gpio_configure[14][12] ),
    .X(net1508));
 sky130_fd_sc_hd__bufbuf_16 hold1047 (.A(_0301_),
    .X(net1509));
 sky130_fd_sc_hd__bufbuf_16 hold1048 (.A(\gpio_configure[2][12] ),
    .X(net1510));
 sky130_fd_sc_hd__bufbuf_16 hold1049 (.A(_0152_),
    .X(net1511));
 sky130_fd_sc_hd__bufbuf_16 hold1050 (.A(\gpio_configure[10][11] ),
    .X(net1512));
 sky130_fd_sc_hd__bufbuf_16 hold1051 (.A(_0215_),
    .X(net1513));
 sky130_fd_sc_hd__bufbuf_16 hold1052 (.A(\gpio_configure[10][12] ),
    .X(net1514));
 sky130_fd_sc_hd__bufbuf_16 hold1053 (.A(_0216_),
    .X(net1515));
 sky130_fd_sc_hd__bufbuf_16 hold1054 (.A(\gpio_configure[23][12] ),
    .X(net1516));
 sky130_fd_sc_hd__bufbuf_16 hold1055 (.A(_0366_),
    .X(net1517));
 sky130_fd_sc_hd__bufbuf_16 hold1056 (.A(\gpio_configure[1][12] ),
    .X(net1518));
 sky130_fd_sc_hd__bufbuf_16 hold1057 (.A(\gpio_configure[0][12] ),
    .X(net1519));
 sky130_fd_sc_hd__bufbuf_16 hold1058 (.A(\gpio_configure[25][12] ),
    .X(net1520));
 sky130_fd_sc_hd__bufbuf_16 hold1059 (.A(_0261_),
    .X(net1521));
 sky130_fd_sc_hd__bufbuf_16 hold1060 (.A(net268),
    .X(net1522));
 sky130_fd_sc_hd__bufbuf_16 hold1061 (.A(net291),
    .X(net1523));
 sky130_fd_sc_hd__bufbuf_16 hold1062 (.A(\gpio_configure[21][0] ),
    .X(net1524));
 sky130_fd_sc_hd__bufbuf_16 hold1063 (.A(\gpio_configure[12][12] ),
    .X(net1525));
 sky130_fd_sc_hd__bufbuf_16 hold1064 (.A(_0226_),
    .X(net1526));
 sky130_fd_sc_hd__bufbuf_16 hold1065 (.A(\gpio_configure[7][12] ),
    .X(net1527));
 sky130_fd_sc_hd__bufbuf_16 hold1066 (.A(_0201_),
    .X(net1528));
 sky130_fd_sc_hd__bufbuf_16 hold1067 (.A(trap_output_dest),
    .X(net1529));
 sky130_fd_sc_hd__bufbuf_16 hold1068 (.A(_0425_),
    .X(net1530));
 sky130_fd_sc_hd__bufbuf_16 hold1069 (.A(\gpio_configure[17][8] ),
    .X(net1531));
 sky130_fd_sc_hd__bufbuf_16 hold1070 (.A(_0312_),
    .X(net1532));
 sky130_fd_sc_hd__bufbuf_16 hold1071 (.A(\gpio_configure[18][0] ),
    .X(net1533));
 sky130_fd_sc_hd__bufbuf_16 hold1072 (.A(\gpio_configure[11][0] ),
    .X(net1534));
 sky130_fd_sc_hd__bufbuf_16 hold1073 (.A(net301),
    .X(net1535));
 sky130_fd_sc_hd__bufbuf_16 hold1074 (.A(_0409_),
    .X(net1536));
 sky130_fd_sc_hd__bufbuf_16 hold1075 (.A(\gpio_configure[6][0] ),
    .X(net1537));
 sky130_fd_sc_hd__bufbuf_16 hold1076 (.A(\gpio_configure[0][0] ),
    .X(net1538));
 sky130_fd_sc_hd__bufbuf_16 hold1077 (.A(\gpio_configure[26][0] ),
    .X(net1539));
 sky130_fd_sc_hd__bufbuf_16 hold1078 (.A(\gpio_configure[23][0] ),
    .X(net1540));
 sky130_fd_sc_hd__bufbuf_16 hold1079 (.A(\gpio_configure[29][0] ),
    .X(net1541));
 sky130_fd_sc_hd__bufbuf_16 hold1080 (.A(\gpio_configure[20][0] ),
    .X(net1542));
 sky130_fd_sc_hd__bufbuf_16 hold1081 (.A(\mgmt_gpio_data[1] ),
    .X(net1543));
 sky130_fd_sc_hd__bufbuf_16 hold1082 (.A(_0281_),
    .X(net1544));
 sky130_fd_sc_hd__bufbuf_16 hold1083 (.A(\gpio_configure[19][0] ),
    .X(net1545));
 sky130_fd_sc_hd__bufbuf_16 hold1084 (.A(net264),
    .X(net1546));
 sky130_fd_sc_hd__bufbuf_16 hold1085 (.A(\gpio_configure[1][2] ),
    .X(net1547));
 sky130_fd_sc_hd__bufbuf_16 hold1086 (.A(_0452_),
    .X(net1548));
 sky130_fd_sc_hd__bufbuf_16 hold1087 (.A(\gpio_configure[30][0] ),
    .X(net1549));
 sky130_fd_sc_hd__bufbuf_16 hold1088 (.A(\gpio_configure[33][11] ),
    .X(net1550));
 sky130_fd_sc_hd__bufbuf_16 hold1089 (.A(_0345_),
    .X(net1551));
 sky130_fd_sc_hd__bufbuf_16 hold1090 (.A(\gpio_configure[33][10] ),
    .X(net1552));
 sky130_fd_sc_hd__bufbuf_16 hold1091 (.A(_0344_),
    .X(net1553));
 sky130_fd_sc_hd__bufbuf_16 hold1092 (.A(\gpio_configure[31][0] ),
    .X(net1554));
 sky130_fd_sc_hd__bufbuf_16 hold1093 (.A(\gpio_configure[16][8] ),
    .X(net1555));
 sky130_fd_sc_hd__bufbuf_16 hold1094 (.A(_0232_),
    .X(net1556));
 sky130_fd_sc_hd__bufbuf_16 hold1095 (.A(\gpio_configure[17][0] ),
    .X(net1557));
 sky130_fd_sc_hd__bufbuf_16 hold1096 (.A(\gpio_configure[22][10] ),
    .X(net1558));
 sky130_fd_sc_hd__bufbuf_16 hold1097 (.A(\gpio_configure[36][12] ),
    .X(net1559));
 sky130_fd_sc_hd__bufbuf_16 hold1098 (.A(\gpio_configure[24][0] ),
    .X(net1560));
 sky130_fd_sc_hd__bufbuf_16 hold1099 (.A(\gpio_configure[2][8] ),
    .X(net1561));
 sky130_fd_sc_hd__bufbuf_16 hold1100 (.A(_0148_),
    .X(net1562));
 sky130_fd_sc_hd__bufbuf_16 hold1101 (.A(\gpio_configure[29][12] ),
    .X(net1563));
 sky130_fd_sc_hd__bufbuf_16 hold1102 (.A(_0256_),
    .X(net1564));
 sky130_fd_sc_hd__bufbuf_16 hold1103 (.A(\gpio_configure[29][10] ),
    .X(net1565));
 sky130_fd_sc_hd__bufbuf_16 hold1104 (.A(\gpio_configure[34][12] ),
    .X(net1566));
 sky130_fd_sc_hd__bufbuf_16 hold1105 (.A(_0336_),
    .X(net1567));
 sky130_fd_sc_hd__bufbuf_16 hold1106 (.A(\gpio_configure[27][0] ),
    .X(net1568));
 sky130_fd_sc_hd__bufbuf_16 hold1107 (.A(\gpio_configure[31][4] ),
    .X(net1569));
 sky130_fd_sc_hd__bufbuf_16 hold1108 (.A(_0694_),
    .X(net1570));
 sky130_fd_sc_hd__bufbuf_16 hold1109 (.A(\gpio_configure[11][8] ),
    .X(net1571));
 sky130_fd_sc_hd__bufbuf_16 hold1110 (.A(_0217_),
    .X(net1572));
 sky130_fd_sc_hd__bufbuf_16 hold1111 (.A(\gpio_configure[28][0] ),
    .X(net1573));
 sky130_fd_sc_hd__bufbuf_16 hold1112 (.A(\gpio_configure[22][0] ),
    .X(net1574));
 sky130_fd_sc_hd__bufbuf_16 hold1113 (.A(\gpio_configure[3][0] ),
    .X(net1575));
 sky130_fd_sc_hd__bufbuf_16 hold1114 (.A(\gpio_configure[23][8] ),
    .X(net1576));
 sky130_fd_sc_hd__bufbuf_16 hold1115 (.A(_0362_),
    .X(net1577));
 sky130_fd_sc_hd__bufbuf_16 hold1116 (.A(\gpio_configure[11][10] ),
    .X(net1578));
 sky130_fd_sc_hd__bufbuf_16 hold1117 (.A(\gpio_configure[16][10] ),
    .X(net1579));
 sky130_fd_sc_hd__bufbuf_16 hold1118 (.A(\gpio_configure[4][10] ),
    .X(net1580));
 sky130_fd_sc_hd__bufbuf_16 hold1119 (.A(\gpio_configure[34][8] ),
    .X(net1581));
 sky130_fd_sc_hd__bufbuf_16 hold1120 (.A(_0332_),
    .X(net1582));
 sky130_fd_sc_hd__bufbuf_16 hold1121 (.A(\gpio_configure[4][8] ),
    .X(net1583));
 sky130_fd_sc_hd__bufbuf_16 hold1122 (.A(_0158_),
    .X(net1584));
 sky130_fd_sc_hd__bufbuf_16 hold1123 (.A(\gpio_configure[9][2] ),
    .X(net1585));
 sky130_fd_sc_hd__bufbuf_16 hold1124 (.A(_0516_),
    .X(net1586));
 sky130_fd_sc_hd__bufbuf_16 hold1125 (.A(\gpio_configure[6][8] ),
    .X(net1587));
 sky130_fd_sc_hd__bufbuf_16 hold1126 (.A(_0184_),
    .X(net1588));
 sky130_fd_sc_hd__bufbuf_16 hold1127 (.A(\gpio_configure[3][8] ),
    .X(net1589));
 sky130_fd_sc_hd__bufbuf_16 hold1128 (.A(_0153_),
    .X(net1590));
 sky130_fd_sc_hd__bufbuf_16 hold1129 (.A(\gpio_configure[9][8] ),
    .X(net1591));
 sky130_fd_sc_hd__bufbuf_16 hold1130 (.A(_0207_),
    .X(net1592));
 sky130_fd_sc_hd__bufbuf_16 hold1131 (.A(\gpio_configure[36][2] ),
    .X(net1593));
 sky130_fd_sc_hd__bufbuf_16 hold1132 (.A(_0732_),
    .X(net1594));
 sky130_fd_sc_hd__bufbuf_16 hold1133 (.A(net172),
    .X(net1595));
 sky130_fd_sc_hd__bufbuf_16 hold1134 (.A(_0414_),
    .X(net1596));
 sky130_fd_sc_hd__bufbuf_16 hold1135 (.A(\gpio_configure[9][10] ),
    .X(net1597));
 sky130_fd_sc_hd__bufbuf_16 hold1136 (.A(\gpio_configure[5][2] ),
    .X(net1598));
 sky130_fd_sc_hd__bufbuf_16 hold1137 (.A(_0484_),
    .X(net1599));
 sky130_fd_sc_hd__bufbuf_16 hold1138 (.A(\gpio_configure[7][8] ),
    .X(net1600));
 sky130_fd_sc_hd__bufbuf_16 hold1139 (.A(_0197_),
    .X(net1601));
 sky130_fd_sc_hd__bufbuf_16 hold1140 (.A(\gpio_configure[10][8] ),
    .X(net1602));
 sky130_fd_sc_hd__bufbuf_16 hold1141 (.A(_0212_),
    .X(net1603));
 sky130_fd_sc_hd__bufbuf_16 hold1142 (.A(\gpio_configure[25][8] ),
    .X(net1604));
 sky130_fd_sc_hd__bufbuf_16 hold1143 (.A(_0257_),
    .X(net1605));
 sky130_fd_sc_hd__bufbuf_16 hold1144 (.A(\gpio_configure[13][8] ),
    .X(net1606));
 sky130_fd_sc_hd__bufbuf_16 hold1145 (.A(_0227_),
    .X(net1607));
 sky130_fd_sc_hd__bufbuf_16 hold1146 (.A(\gpio_configure[10][2] ),
    .X(net1608));
 sky130_fd_sc_hd__bufbuf_16 hold1147 (.A(_0524_),
    .X(net1609));
 sky130_fd_sc_hd__bufbuf_16 hold1148 (.A(\gpio_configure[3][2] ),
    .X(net1610));
 sky130_fd_sc_hd__bufbuf_16 hold1149 (.A(_0468_),
    .X(net1611));
 sky130_fd_sc_hd__bufbuf_16 hold1150 (.A(\gpio_configure[37][8] ),
    .X(net1612));
 sky130_fd_sc_hd__bufbuf_16 hold1151 (.A(_0307_),
    .X(net1613));
 sky130_fd_sc_hd__bufbuf_16 hold1152 (.A(\gpio_configure[8][2] ),
    .X(net1614));
 sky130_fd_sc_hd__bufbuf_16 hold1153 (.A(_0508_),
    .X(net1615));
 sky130_fd_sc_hd__bufbuf_16 hold1154 (.A(\gpio_configure[31][8] ),
    .X(net1616));
 sky130_fd_sc_hd__bufbuf_16 hold1155 (.A(_0242_),
    .X(net1617));
 sky130_fd_sc_hd__bufbuf_16 hold1156 (.A(\gpio_configure[6][2] ),
    .X(net1618));
 sky130_fd_sc_hd__bufbuf_16 hold1157 (.A(_0492_),
    .X(net1619));
 sky130_fd_sc_hd__bufbuf_16 hold1158 (.A(\gpio_configure[27][8] ),
    .X(net1620));
 sky130_fd_sc_hd__bufbuf_16 hold1159 (.A(_0809_),
    .X(net1621));
 sky130_fd_sc_hd__bufbuf_16 hold1160 (.A(\gpio_configure[2][2] ),
    .X(net1622));
 sky130_fd_sc_hd__bufbuf_16 hold1161 (.A(_0460_),
    .X(net1623));
 sky130_fd_sc_hd__bufbuf_16 hold1162 (.A(\gpio_configure[34][10] ),
    .X(net1624));
 sky130_fd_sc_hd__bufbuf_16 hold1163 (.A(\gpio_configure[14][8] ),
    .X(net1625));
 sky130_fd_sc_hd__bufbuf_16 hold1164 (.A(_0297_),
    .X(net1626));
 sky130_fd_sc_hd__bufbuf_16 hold1165 (.A(\gpio_configure[28][8] ),
    .X(net1627));
 sky130_fd_sc_hd__bufbuf_16 hold1166 (.A(_0262_),
    .X(net1628));
 sky130_fd_sc_hd__bufbuf_16 hold1167 (.A(\gpio_configure[12][8] ),
    .X(net1629));
 sky130_fd_sc_hd__bufbuf_16 hold1168 (.A(_0222_),
    .X(net1630));
 sky130_fd_sc_hd__bufbuf_16 hold1169 (.A(\gpio_configure[37][10] ),
    .X(net1631));
 sky130_fd_sc_hd__bufbuf_16 hold1170 (.A(_0309_),
    .X(net1632));
 sky130_fd_sc_hd__bufbuf_16 hold1171 (.A(net282),
    .X(net1633));
 sky130_fd_sc_hd__bufbuf_16 hold1172 (.A(_0400_),
    .X(net1634));
 sky130_fd_sc_hd__bufbuf_16 hold1173 (.A(\gpio_configure[36][8] ),
    .X(net1635));
 sky130_fd_sc_hd__bufbuf_16 hold1174 (.A(_0237_),
    .X(net1636));
 sky130_fd_sc_hd__bufbuf_16 hold1175 (.A(\gpio_configure[18][8] ),
    .X(net1637));
 sky130_fd_sc_hd__bufbuf_16 hold1176 (.A(_0317_),
    .X(net1638));
 sky130_fd_sc_hd__bufbuf_16 hold1177 (.A(\gpio_configure[26][8] ),
    .X(net1639));
 sky130_fd_sc_hd__bufbuf_16 hold1178 (.A(_0267_),
    .X(net1640));
 sky130_fd_sc_hd__bufbuf_16 hold1179 (.A(\gpio_configure[5][8] ),
    .X(net1641));
 sky130_fd_sc_hd__bufbuf_16 hold1180 (.A(_0171_),
    .X(net1642));
 sky130_fd_sc_hd__bufbuf_16 hold1181 (.A(\gpio_configure[12][2] ),
    .X(net1643));
 sky130_fd_sc_hd__bufbuf_16 hold1182 (.A(_0540_),
    .X(net1644));
 sky130_fd_sc_hd__bufbuf_16 hold1183 (.A(hkspi_disable),
    .X(net1645));
 sky130_fd_sc_hd__bufbuf_16 hold1184 (.A(_0422_),
    .X(net1646));
 sky130_fd_sc_hd__bufbuf_16 hold1185 (.A(\gpio_configure[30][8] ),
    .X(net1647));
 sky130_fd_sc_hd__bufbuf_16 hold1186 (.A(_0374_),
    .X(net1648));
 sky130_fd_sc_hd__bufbuf_16 hold1187 (.A(\gpio_configure[13][2] ),
    .X(net1649));
 sky130_fd_sc_hd__bufbuf_16 hold1188 (.A(_0548_),
    .X(net1650));
 sky130_fd_sc_hd__bufbuf_16 hold1189 (.A(net272),
    .X(net1651));
 sky130_fd_sc_hd__bufbuf_16 hold1190 (.A(_0394_),
    .X(net1652));
 sky130_fd_sc_hd__bufbuf_16 hold1191 (.A(\gpio_configure[2][10] ),
    .X(net1653));
 sky130_fd_sc_hd__bufbuf_16 hold1192 (.A(\gpio_configure[20][8] ),
    .X(net1654));
 sky130_fd_sc_hd__bufbuf_16 hold1193 (.A(_0337_),
    .X(net1655));
 sky130_fd_sc_hd__bufbuf_16 hold1194 (.A(\gpio_configure[19][8] ),
    .X(net1656));
 sky130_fd_sc_hd__bufbuf_16 hold1195 (.A(_0327_),
    .X(net1657));
 sky130_fd_sc_hd__bufbuf_16 hold1196 (.A(net266),
    .X(net1658));
 sky130_fd_sc_hd__bufbuf_16 hold1197 (.A(_0389_),
    .X(net1659));
 sky130_fd_sc_hd__bufbuf_16 hold1198 (.A(serial_xfer),
    .X(net1660));
 sky130_fd_sc_hd__bufbuf_16 hold1199 (.A(_0421_),
    .X(net1661));
 sky130_fd_sc_hd__bufbuf_16 hold1200 (.A(reset_reg),
    .X(net1662));
 sky130_fd_sc_hd__bufbuf_16 hold1201 (.A(_0413_),
    .X(net1663));
 sky130_fd_sc_hd__bufbuf_16 hold1202 (.A(\gpio_configure[37][12] ),
    .X(net1664));
 sky130_fd_sc_hd__bufbuf_16 hold1203 (.A(net299),
    .X(net1665));
 sky130_fd_sc_hd__bufbuf_16 hold1204 (.A(_0096_),
    .X(net1666));
 sky130_fd_sc_hd__bufbuf_16 hold1205 (.A(\gpio_configure[8][8] ),
    .X(net1667));
 sky130_fd_sc_hd__bufbuf_16 hold1206 (.A(_0202_),
    .X(net1668));
 sky130_fd_sc_hd__bufbuf_16 hold1207 (.A(net271),
    .X(net1669));
 sky130_fd_sc_hd__bufbuf_16 hold1208 (.A(_0387_),
    .X(net1670));
 sky130_fd_sc_hd__bufbuf_16 hold1209 (.A(\mgmt_gpio_data[32] ),
    .X(net1671));
 sky130_fd_sc_hd__bufbuf_16 hold1210 (.A(_0428_),
    .X(net1672));
 sky130_fd_sc_hd__bufbuf_16 hold1211 (.A(\gpio_configure[21][8] ),
    .X(net1673));
 sky130_fd_sc_hd__bufbuf_16 hold1212 (.A(_0347_),
    .X(net1674));
 sky130_fd_sc_hd__bufbuf_16 hold1213 (.A(\gpio_configure[1][8] ),
    .X(net1675));
 sky130_fd_sc_hd__bufbuf_16 hold1214 (.A(_0143_),
    .X(net1676));
 sky130_fd_sc_hd__bufbuf_16 hold1215 (.A(\gpio_configure[22][8] ),
    .X(net1677));
 sky130_fd_sc_hd__bufbuf_16 hold1216 (.A(_0357_),
    .X(net1678));
 sky130_fd_sc_hd__bufbuf_16 hold1217 (.A(\gpio_configure[15][8] ),
    .X(net1679));
 sky130_fd_sc_hd__bufbuf_16 hold1218 (.A(_0302_),
    .X(net1680));
 sky130_fd_sc_hd__bufbuf_16 hold1219 (.A(net275),
    .X(net1681));
 sky130_fd_sc_hd__bufbuf_16 hold1220 (.A(\gpio_configure[33][8] ),
    .X(net1682));
 sky130_fd_sc_hd__bufbuf_16 hold1221 (.A(_0342_),
    .X(net1683));
 sky130_fd_sc_hd__bufbuf_16 hold1222 (.A(\gpio_configure[29][8] ),
    .X(net1684));
 sky130_fd_sc_hd__bufbuf_16 hold1223 (.A(_0252_),
    .X(net1685));
 sky130_fd_sc_hd__bufbuf_16 hold1224 (.A(irq_1_inputsrc),
    .X(net1686));
 sky130_fd_sc_hd__bufbuf_16 hold1225 (.A(_0426_),
    .X(net1687));
 sky130_fd_sc_hd__bufbuf_16 hold1226 (.A(\mgmt_gpio_data[0] ),
    .X(net1688));
 sky130_fd_sc_hd__bufbuf_16 hold1227 (.A(_0280_),
    .X(net1689));
 sky130_fd_sc_hd__bufbuf_16 hold1228 (.A(\gpio_configure[24][8] ),
    .X(net1690));
 sky130_fd_sc_hd__bufbuf_16 hold1229 (.A(_0247_),
    .X(net1691));
 sky130_fd_sc_hd__bufbuf_16 hold1230 (.A(\gpio_configure[0][8] ),
    .X(net1692));
 sky130_fd_sc_hd__bufbuf_16 hold1231 (.A(_0138_),
    .X(net1693));
 sky130_fd_sc_hd__bufbuf_16 hold1232 (.A(\gpio_configure[32][8] ),
    .X(net1694));
 sky130_fd_sc_hd__bufbuf_16 hold1233 (.A(_0352_),
    .X(net1695));
 sky130_fd_sc_hd__bufbuf_16 hold1234 (.A(\mgmt_gpio_data_buf[14] ),
    .X(net1696));
 sky130_fd_sc_hd__bufbuf_16 hold1235 (.A(_0136_),
    .X(net1697));
 sky130_fd_sc_hd__bufbuf_16 hold1236 (.A(\mgmt_gpio_data_buf[21] ),
    .X(net1698));
 sky130_fd_sc_hd__bufbuf_16 hold1237 (.A(\mgmt_gpio_data_buf[8] ),
    .X(net1699));
 sky130_fd_sc_hd__bufbuf_16 hold1238 (.A(\mgmt_gpio_data_buf[3] ),
    .X(net1700));
 sky130_fd_sc_hd__bufbuf_16 hold1239 (.A(\mgmt_gpio_data_buf[23] ),
    .X(net1701));
 sky130_fd_sc_hd__bufbuf_16 hold1240 (.A(net225),
    .X(net1702));
 sky130_fd_sc_hd__bufbuf_16 hold1241 (.A(\gpio_configure[31][7] ),
    .X(net1703));
 sky130_fd_sc_hd__bufbuf_16 hold1242 (.A(\gpio_configure[1][7] ),
    .X(net1704));
 sky130_fd_sc_hd__bufbuf_16 hold1243 (.A(\gpio_configure[32][7] ),
    .X(net1705));
 sky130_fd_sc_hd__bufbuf_16 hold1244 (.A(\gpio_configure[12][9] ),
    .X(net1706));
 sky130_fd_sc_hd__bufbuf_16 hold1245 (.A(serial_bb_load),
    .X(net1707));
 sky130_fd_sc_hd__bufbuf_16 hold1246 (.A(\gpio_configure[32][5] ),
    .X(net1708));
 sky130_fd_sc_hd__bufbuf_16 hold1247 (.A(\gpio_configure[0][7] ),
    .X(net1709));
 sky130_fd_sc_hd__bufbuf_16 hold1248 (.A(\gpio_configure[5][11] ),
    .X(net1710));
 sky130_fd_sc_hd__bufbuf_16 hold1249 (.A(\gpio_configure[13][12] ),
    .X(net1711));
 sky130_fd_sc_hd__bufbuf_16 hold1250 (.A(\gpio_configure[27][2] ),
    .X(net1712));
 sky130_fd_sc_hd__bufbuf_16 hold1251 (.A(\gpio_configure[30][2] ),
    .X(net1713));
 sky130_fd_sc_hd__bufbuf_16 hold1252 (.A(\gpio_configure[13][7] ),
    .X(net1714));
 sky130_fd_sc_hd__bufbuf_16 hold1253 (.A(\gpio_configure[17][5] ),
    .X(net1715));
 sky130_fd_sc_hd__bufbuf_16 hold1254 (.A(\gpio_configure[35][2] ),
    .X(net1716));
 sky130_fd_sc_hd__bufbuf_16 hold1255 (.A(\gpio_configure[1][5] ),
    .X(net1717));
 sky130_fd_sc_hd__bufbuf_16 hold1256 (.A(serial_bb_clock),
    .X(net1718));
 sky130_fd_sc_hd__bufbuf_16 hold1257 (.A(\gpio_configure[29][2] ),
    .X(net1719));
 sky130_fd_sc_hd__bufbuf_16 hold1258 (.A(\gpio_configure[23][4] ),
    .X(net1720));
 sky130_fd_sc_hd__bufbuf_16 hold1259 (.A(\gpio_configure[36][6] ),
    .X(net1721));
 sky130_fd_sc_hd__bufbuf_16 hold1260 (.A(\gpio_configure[18][2] ),
    .X(net1722));
 sky130_fd_sc_hd__bufbuf_16 hold1261 (.A(net304),
    .X(net1723));
 sky130_fd_sc_hd__bufbuf_16 hold1262 (.A(\gpio_configure[11][2] ),
    .X(net1724));
 sky130_fd_sc_hd__bufbuf_16 hold1263 (.A(\gpio_configure[21][2] ),
    .X(net1725));
 sky130_fd_sc_hd__bufbuf_16 hold1264 (.A(\gpio_configure[25][3] ),
    .X(net1726));
 sky130_fd_sc_hd__bufbuf_16 hold1265 (.A(\mgmt_gpio_data_buf[19] ),
    .X(net1727));
 sky130_fd_sc_hd__bufbuf_16 hold1266 (.A(\mgmt_gpio_data_buf[17] ),
    .X(net1728));
 sky130_fd_sc_hd__bufbuf_16 hold1267 (.A(\gpio_configure[33][1] ),
    .X(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0106_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0371_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_1189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_1271_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_1534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_2426_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_2509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_2519_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_2530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_2532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_2532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_2533_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_2560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_2563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_2802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_2817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_2817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_3188_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(debug_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(debug_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(debug_out));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(\gpio_configure[14][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(\gpio_configure[17][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(\gpio_configure[18][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\gpio_configure[18][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\gpio_configure[18][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\gpio_configure[25][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\gpio_configure[28][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\gpio_configure[30][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\gpio_configure[36][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\hkspi.addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\hkspi.addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\hkspi.addr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\hkspi.count[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\hkspi.pre_pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(mask_rev_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(mask_rev_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(mask_rev_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(mask_rev_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(mask_rev_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(mask_rev_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(mask_rev_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(mask_rev_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(mask_rev_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(mask_rev_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(mask_rev_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(mask_rev_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(mask_rev_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(mask_rev_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(mask_rev_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(mask_rev_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(mask_rev_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(mask_rev_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\mgmt_gpio_data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(\pad_count_1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(pad_flash_io0_di));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(pad_flash_io1_di));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(ser_tx));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(serial_load_pre));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(spi_csb));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(spi_sck));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(spi_sdoenb));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(spimemio_flash_io3_do));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(spimemio_flash_io3_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(wb_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(wb_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(wb_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(wb_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(wb_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(wb_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(wb_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(wb_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(wb_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(wb_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(wb_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(wb_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(wb_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(wb_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(wb_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(wb_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(wb_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(wb_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(wb_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(wb_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(wb_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(wb_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(wb_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(wb_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(wb_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net1665));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net1669));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net1681));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net1717));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(_1046_));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(_1094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(_2513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(_2752_));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(\hkspi.addr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(\hkspi.count[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(mask_rev_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(\xfer_count[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(net1656));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(_0109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(_2522_));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(_2826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(\gpio_configure[32][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(\hkspi.count[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(\hkspi.count[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(net1104));
 sky130_fd_sc_hd__fill_1 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_771 ();
endmodule
