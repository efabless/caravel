magic
tech sky130A
magscale 1 2
timestamp 1637517609
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< error_s >>
rect 673388 990096 673420 992100
rect 673708 989776 673740 991780
rect 14347 602956 14630 602979
rect 14347 602256 14630 602280
rect 24204 600834 24270 600837
rect 21493 600820 24270 600834
rect 8262 599198 8551 599222
rect 17475 598150 17744 598174
rect 17424 597830 17795 597852
rect 8262 597508 8551 597532
rect 17104 597510 17475 597532
rect 17475 596460 17744 596484
rect 17424 596140 17795 596162
rect 8262 595818 8551 595841
rect 17104 595820 17475 595842
rect 17475 594770 17744 594794
rect 17424 594450 17795 594472
rect 8262 594128 8551 594152
rect 17104 594130 17475 594152
rect 17475 593080 17744 593104
rect 17424 592760 17795 592782
rect 8294 592438 8551 592462
rect 17104 592440 17475 592462
rect 17475 591390 17744 591414
rect 17424 591070 17795 591092
rect 8294 590748 8551 590770
rect 17104 590750 17475 590772
rect 17475 589700 17744 589724
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 953022 710788 965190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use open_source  open_source_0 hexdigits
timestamp 1635801696
transform 1 0 205230 0 1 2174
box 752 5164 29030 16242
use copyright_block_a  copyright_block_a_0
timestamp 1636248774
transform 1 0 149582 0 1 16298
box -262 -9464 35048 2764
use caravan_logo  caravan_logo_0
timestamp 1636751500
transform 1 0 255642 0 1 5786
box 2240 2560 37000 11520
use housekeeping  housekeeping_0
timestamp 1637412603
transform 1 0 602468 0 1 95484
box 0 0 60046 110190
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1636217749
transform -1 0 709467 0 1 131400
box -38 0 6018 2224
use caravel_clocking  caravel_clocking_0
timestamp 1637348273
transform 1 0 649886 0 1 70896
box -38 -48 20000 12000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1637411465
transform -1 0 710203 0 1 118400
box 882 167 34000 13000
use simple_por  simple_por_0
timestamp 1606688983
transform 1 0 624040 0 1 45166
box 0 0 11344 8338
use xres_buf  xres_buf_0
timestamp 1608587411
transform 1 0 608050 0 1 79488
box 414 -400 3522 3800
use user_id_programming  user_id_programming_0
timestamp 1606755340
transform 1 0 635116 0 1 79088
box 0 0 7109 7077
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1636217749
transform 1 0 8367 0 1 212600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1637411465
transform 1 0 7631 0 1 199600
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1636217749
transform -1 0 709467 0 1 177000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1637411465
transform -1 0 710203 0 1 164000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1637411465
transform -1 0 710203 0 1 208400
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1636217749
transform 1 0 8367 0 1 255800
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1637411465
transform 1 0 7631 0 1 242800
box 882 167 34000 13000
use mgmt_protect  mgmt_protect_0
timestamp 1637329592
transform 1 0 206090 0 1 227796
box -400 -400 220400 32400
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1636217749
transform -1 0 709467 0 1 221400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1636217749
transform -1 0 709467 0 1 266600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1637411465
transform -1 0 710203 0 1 253600
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1636217749
transform 1 0 8367 0 1 299000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1637411465
transform 1 0 7631 0 1 286000
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1636217749
transform -1 0 709467 0 1 311800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1637411465
transform -1 0 710203 0 1 298800
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1636217749
transform 1 0 8367 0 1 475400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1636217749
transform 1 0 8367 0 1 428000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1636217749
transform 1 0 8367 0 1 385400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1636217749
transform 1 0 8367 0 1 342200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1637411465
transform 1 0 7631 0 1 372400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1637411465
transform 1 0 7631 0 1 329200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1637411465
transform 1 0 7631 0 1 415000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1637411465
transform 1 0 7631 0 1 462400
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1636217749
transform -1 0 709467 0 1 357600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1636217749
transform -1 0 709467 0 1 402000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1636217749
transform -1 0 709467 0 1 490200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1637411465
transform -1 0 710203 0 1 344600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1637411465
transform -1 0 710203 0 1 389000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1637411465
transform -1 0 710203 0 1 477200
box 882 167 34000 13000
use mgmt_core_wrapper  mgmt_core_wrapper_0
timestamp 1637416673
transform 1 0 56746 0 1 42404
box 382 -400 524400 164400
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1636217749
transform 1 0 8367 0 1 601224
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1637411465
transform 1 0 7631 0 1 588224
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1637411465
transform 1 0 7631 0 1 631400
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1636217749
transform -1 0 709467 0 1 534600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1636217749
transform -1 0 709467 0 1 577800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1636217749
transform -1 0 709467 0 1 624800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1637411465
transform -1 0 710203 0 1 611800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1637411465
transform -1 0 710203 0 1 564800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1637411465
transform -1 0 710203 0 1 521600
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1636217749
transform 1 0 8367 0 1 730800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1636217749
transform 1 0 8367 0 1 687600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1636217749
transform 1 0 8367 0 1 644400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1637411465
transform 1 0 7631 0 1 674600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1637411465
transform 1 0 7631 0 1 717800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1637411465
transform 1 0 7631 0 1 761000
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1636217749
transform -1 0 709467 0 1 670000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1636217749
transform -1 0 709467 0 1 715000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1637411465
transform -1 0 710203 0 1 657000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1637411465
transform -1 0 710203 0 1 702000
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1636217749
transform 1 0 8367 0 1 817200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1636217749
transform 1 0 8367 0 1 774000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1637411465
transform 1 0 7631 0 1 804200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1637411465
transform -1 0 710203 0 1 880800
box 882 167 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1636217749
transform -1 0 709467 0 1 893800
box -38 0 6018 2224
use chip_io_alt  padframe
timestamp 1637517609
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_analog_project_wrapper  user_analog_project_wrapper_0
timestamp 1620244087
transform 1 0 64268 0 1 282662
box -800 -800 584800 704800
use caravan_power_routing  caravan_power_routing_0
timestamp 1637449042
transform 1 0 0 0 1 -2600
box 0 2400 717600 1040000
<< labels >>
flabel metal5 s 187640 6598 200180 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363580 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308780 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418380 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473180 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527980 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030788 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030788 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030788 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158980 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030788 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030788 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030788 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030788 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6811 956610 18975 968778 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203980 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227020 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183820 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249180 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294180 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339180 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384380 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1
port 45 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2
port 46 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda
port 47 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1
port 48 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 49 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2
port 50 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_2
port 51 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1
port 52 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 53 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2
port 54 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1
port 55 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2
port 56 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_2
port 57 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio
port 58 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio
port 59 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa
port 60 nsew signal bidirectional
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd
port 61 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd
port 62 nsew signal bidirectional
flabel metal5 s 698624 953022 710788 965190 0 FreeSans 16000 0 0 0 mprj_io[14]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030788 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030788 0 FreeSans 16000 0 0 0 mprj_io[18]
port 11 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
