magic
tech sky130A
magscale 1 2
timestamp 1649446267
<< checkpaint >>
rect -378 4132 11142 12732
rect -102 372 11142 4132
rect 1738 -220 11142 372
<< isosubstrate >>
rect 1018 1528 2810 4514
<< viali >>
rect 3893 11305 3927 11339
rect 4077 11305 4111 11339
rect 5917 11305 5951 11339
rect 6377 11305 6411 11339
rect 7941 11305 7975 11339
rect 4445 11237 4479 11271
rect 9137 11237 9171 11271
rect 9505 11237 9539 11271
rect 5733 11169 5767 11203
rect 8125 11169 8159 11203
rect 1869 11101 1903 11135
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2697 11101 2731 11135
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 4261 11101 4295 11135
rect 4537 11101 4571 11135
rect 4905 11101 4939 11135
rect 5641 11101 5675 11135
rect 7481 11101 7515 11135
rect 7757 11101 7791 11135
rect 8033 11101 8067 11135
rect 8585 11101 8619 11135
rect 2513 11033 2547 11067
rect 2973 11033 3007 11067
rect 4721 11033 4755 11067
rect 4997 11033 5031 11067
rect 5181 11033 5215 11067
rect 5365 11033 5399 11067
rect 6837 11033 6871 11067
rect 6929 11033 6963 11067
rect 7573 11033 7607 11067
rect 8493 11033 8527 11067
rect 8769 11033 8803 11067
rect 2053 10965 2087 10999
rect 2421 10965 2455 10999
rect 3341 10965 3375 10999
rect 3617 10965 3651 10999
rect 5457 10965 5491 10999
rect 6193 10965 6227 10999
rect 7113 10965 7147 10999
rect 7297 10965 7331 10999
rect 9229 10965 9263 10999
rect 1409 10761 1443 10795
rect 4905 10761 4939 10795
rect 5089 10761 5123 10795
rect 5917 10761 5951 10795
rect 7573 10761 7607 10795
rect 7849 10761 7883 10795
rect 9505 10761 9539 10795
rect 7113 10693 7147 10727
rect 1593 10625 1627 10659
rect 1869 10625 1903 10659
rect 3709 10625 3743 10659
rect 4445 10625 4479 10659
rect 5462 10623 5496 10657
rect 6198 10625 6232 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7665 10625 7699 10659
rect 7941 10625 7975 10659
rect 8309 10625 8343 10659
rect 9321 10625 9355 10659
rect 2237 10557 2271 10591
rect 5273 10557 5307 10591
rect 4273 10489 4307 10523
rect 7389 10489 7423 10523
rect 8125 10489 8159 10523
rect 1685 10421 1719 10455
rect 4721 10421 4755 10455
rect 5733 10421 5767 10455
rect 6285 10421 6319 10455
rect 6653 10421 6687 10455
rect 8493 10421 8527 10455
rect 8677 10421 8711 10455
rect 2697 10217 2731 10251
rect 3249 10217 3283 10251
rect 3893 10217 3927 10251
rect 5549 10149 5583 10183
rect 2881 10081 2915 10115
rect 6469 10081 6503 10115
rect 1317 10013 1351 10047
rect 1961 10013 1995 10047
rect 2053 10013 2087 10047
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 6101 10013 6135 10047
rect 7941 10013 7975 10047
rect 9413 10013 9447 10047
rect 4261 9945 4295 9979
rect 8769 9945 8803 9979
rect 4077 9877 4111 9911
rect 8505 9877 8539 9911
rect 6745 9673 6779 9707
rect 6193 9605 6227 9639
rect 6561 9605 6595 9639
rect 3249 9537 3283 9571
rect 5365 9537 5399 9571
rect 6377 9537 6411 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 8769 9537 8803 9571
rect 1317 9469 1351 9503
rect 3065 9469 3099 9503
rect 3525 9469 3559 9503
rect 3893 9469 3927 9503
rect 7297 9469 7331 9503
rect 5929 9401 5963 9435
rect 2807 9333 2841 9367
rect 3433 9333 3467 9367
rect 9333 9333 9367 9367
rect 3065 9129 3099 9163
rect 3985 9129 4019 9163
rect 4169 9129 4203 9163
rect 4537 9129 4571 9163
rect 4905 9129 4939 9163
rect 5457 9129 5491 9163
rect 9413 9129 9447 9163
rect 5733 9061 5767 9095
rect 7941 8993 7975 9027
rect 1317 8925 1351 8959
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 3433 8925 3467 8959
rect 3801 8925 3835 8959
rect 3893 8925 3927 8959
rect 4353 8925 4387 8959
rect 5089 8925 5123 8959
rect 5825 8925 5859 8959
rect 6193 8925 6227 8959
rect 8309 8925 8343 8959
rect 8769 8925 8803 8959
rect 2789 8857 2823 8891
rect 2973 8857 3007 8891
rect 4629 8857 4663 8891
rect 5181 8857 5215 8891
rect 5365 8857 5399 8891
rect 6009 8857 6043 8891
rect 6469 8857 6503 8891
rect 8125 8857 8159 8891
rect 2697 8789 2731 8823
rect 3341 8789 3375 8823
rect 3617 8789 3651 8823
rect 8493 8789 8527 8823
rect 1409 8585 1443 8619
rect 1593 8585 1627 8619
rect 6469 8585 6503 8619
rect 6929 8585 6963 8619
rect 9505 8585 9539 8619
rect 5365 8517 5399 8551
rect 5825 8517 5859 8551
rect 1869 8449 1903 8483
rect 2237 8449 2271 8483
rect 3709 8449 3743 8483
rect 4445 8449 4479 8483
rect 5181 8449 5215 8483
rect 5641 8449 5675 8483
rect 6193 8449 6227 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7021 8449 7055 8483
rect 7389 8449 7423 8483
rect 9321 8449 9355 8483
rect 1777 8381 1811 8415
rect 7665 8381 7699 8415
rect 4273 8313 4307 8347
rect 5549 8313 5583 8347
rect 9137 8313 9171 8347
rect 5089 8245 5123 8279
rect 5917 8245 5951 8279
rect 6377 8245 6411 8279
rect 7205 8245 7239 8279
rect 4261 8041 4295 8075
rect 4813 8041 4847 8075
rect 5273 8041 5307 8075
rect 6285 8041 6319 8075
rect 6469 8041 6503 8075
rect 9413 8041 9447 8075
rect 5641 7973 5675 8007
rect 3341 7905 3375 7939
rect 1501 7837 1535 7871
rect 1593 7837 1627 7871
rect 3617 7837 3651 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 6009 7837 6043 7871
rect 6653 7837 6687 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 8769 7837 8803 7871
rect 1869 7769 1903 7803
rect 5825 7769 5859 7803
rect 7389 7769 7423 7803
rect 7573 7769 7607 7803
rect 8585 7769 8619 7803
rect 1409 7701 1443 7735
rect 4445 7701 4479 7735
rect 5457 7701 5491 7735
rect 7297 7701 7331 7735
rect 7941 7701 7975 7735
rect 8309 7701 8343 7735
rect 8401 7701 8435 7735
rect 1317 7497 1351 7531
rect 5925 7497 5959 7531
rect 9137 7497 9171 7531
rect 2789 7429 2823 7463
rect 3065 7361 3099 7395
rect 3249 7361 3283 7395
rect 3525 7361 3559 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 8401 7361 8435 7395
rect 9321 7361 9355 7395
rect 3893 7293 3927 7327
rect 6929 7293 6963 7327
rect 6193 7225 6227 7259
rect 9413 7225 9447 7259
rect 3341 7157 3375 7191
rect 8585 7157 8619 7191
rect 8965 7157 8999 7191
rect 1758 6953 1792 6987
rect 7407 6953 7441 6987
rect 9045 6953 9079 6987
rect 9413 6953 9447 6987
rect 1501 6817 1535 6851
rect 4997 6817 5031 6851
rect 5089 6817 5123 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 3617 6749 3651 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 5733 6749 5767 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 1409 6681 1443 6715
rect 3249 6613 3283 6647
rect 5917 6613 5951 6647
rect 9229 6613 9263 6647
rect 1409 6409 1443 6443
rect 1593 6409 1627 6443
rect 3249 6409 3283 6443
rect 9413 6409 9447 6443
rect 7941 6341 7975 6375
rect 8217 6341 8251 6375
rect 2329 6273 2363 6307
rect 2421 6273 2455 6307
rect 3341 6273 3375 6307
rect 5181 6273 5215 6307
rect 8033 6273 8067 6307
rect 8493 6273 8527 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9321 6273 9355 6307
rect 1685 6205 1719 6239
rect 3065 6205 3099 6239
rect 3709 6205 3743 6239
rect 6193 6205 6227 6239
rect 8585 6205 8619 6239
rect 5745 6137 5779 6171
rect 8401 6137 8435 6171
rect 5917 6069 5951 6103
rect 1501 5865 1535 5899
rect 4261 5865 4295 5899
rect 8309 5865 8343 5899
rect 8861 5865 8895 5899
rect 9229 5797 9263 5831
rect 1317 5729 1351 5763
rect 5917 5729 5951 5763
rect 3433 5661 3467 5695
rect 3617 5661 3651 5695
rect 4445 5661 4479 5695
rect 5549 5661 5583 5695
rect 7941 5661 7975 5695
rect 8585 5661 8619 5695
rect 9045 5661 9079 5695
rect 9321 5661 9355 5695
rect 3157 5593 3191 5627
rect 6193 5593 6227 5627
rect 1685 5525 1719 5559
rect 8125 5525 8159 5559
rect 9413 5525 9447 5559
rect 3525 5321 3559 5355
rect 3801 5321 3835 5355
rect 4077 5321 4111 5355
rect 6469 5321 6503 5355
rect 8493 5321 8527 5355
rect 5181 5253 5215 5287
rect 8861 5253 8895 5287
rect 3341 5185 3375 5219
rect 3617 5185 3651 5219
rect 3893 5185 3927 5219
rect 4353 5185 4387 5219
rect 5089 5185 5123 5219
rect 7021 5185 7055 5219
rect 7665 5185 7699 5219
rect 7849 5185 7883 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 4169 5049 4203 5083
rect 7481 5049 7515 5083
rect 4629 4981 4663 5015
rect 4813 4981 4847 5015
rect 7297 4981 7331 5015
rect 7941 4981 7975 5015
rect 8585 4981 8619 5015
rect 9321 4981 9355 5015
rect 3801 4777 3835 4811
rect 4445 4777 4479 4811
rect 4813 4777 4847 4811
rect 8873 4777 8907 4811
rect 5549 4709 5583 4743
rect 6193 4709 6227 4743
rect 6837 4641 6871 4675
rect 3617 4573 3651 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 5917 4573 5951 4607
rect 6377 4573 6411 4607
rect 6469 4573 6503 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 4997 4505 5031 4539
rect 5733 4505 5767 4539
rect 6101 4505 6135 4539
rect 3525 4437 3559 4471
rect 4169 4437 4203 4471
rect 9045 4437 9079 4471
rect 9321 4437 9355 4471
rect 3801 4233 3835 4267
rect 7481 4233 7515 4267
rect 3617 4165 3651 4199
rect 6929 4165 6963 4199
rect 3985 4097 4019 4131
rect 4261 4097 4295 4131
rect 6101 4097 6135 4131
rect 6665 4097 6699 4131
rect 7205 4097 7239 4131
rect 7665 4097 7699 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 9137 4097 9171 4131
rect 9229 4097 9263 4131
rect 9505 4097 9539 4131
rect 3433 4029 3467 4063
rect 4629 4029 4663 4063
rect 7297 4029 7331 4063
rect 7113 3961 7147 3995
rect 9321 3961 9355 3995
rect 4169 3893 4203 3927
rect 7757 3893 7791 3927
rect 7941 3893 7975 3927
rect 8953 3893 8987 3927
rect 3617 3689 3651 3723
rect 6377 3689 6411 3723
rect 9149 3689 9183 3723
rect 3433 3621 3467 3655
rect 4445 3621 4479 3655
rect 4813 3621 4847 3655
rect 5457 3553 5491 3587
rect 6745 3553 6779 3587
rect 3893 3485 3927 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 5181 3485 5215 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6653 3485 6687 3519
rect 7113 3485 7147 3519
rect 8585 3485 8619 3519
rect 9505 3485 9539 3519
rect 4997 3417 5031 3451
rect 3801 3349 3835 3383
rect 4169 3349 4203 3383
rect 4721 3349 4755 3383
rect 6469 3349 6503 3383
rect 9321 3349 9355 3383
rect 3525 3145 3559 3179
rect 8033 3145 8067 3179
rect 6561 3077 6595 3111
rect 8769 3077 8803 3111
rect 8861 3077 8895 3111
rect 3617 3009 3651 3043
rect 5457 3009 5491 3043
rect 3985 2941 4019 2975
rect 6285 2941 6319 2975
rect 8309 2941 8343 2975
rect 8493 2941 8527 2975
rect 9413 2941 9447 2975
rect 6021 2805 6055 2839
rect 3433 2601 3467 2635
rect 8309 2601 8343 2635
rect 9137 2601 9171 2635
rect 5181 2397 5215 2431
rect 5365 2397 5399 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6101 2397 6135 2431
rect 7573 2397 7607 2431
rect 8953 2397 8987 2431
rect 9229 2397 9263 2431
rect 9505 2397 9539 2431
rect 4905 2329 4939 2363
rect 8137 2329 8171 2363
rect 9321 2261 9355 2295
rect 8677 2057 8711 2091
rect 8309 1989 8343 2023
rect 4261 1921 4295 1955
rect 6193 1921 6227 1955
rect 9413 1921 9447 1955
rect 4537 1853 4571 1887
rect 6009 1853 6043 1887
rect 6469 1853 6503 1887
rect 8769 1853 8803 1887
rect 7941 1717 7975 1751
rect 5089 1513 5123 1547
rect 6101 1513 6135 1547
rect 3617 1377 3651 1411
rect 8125 1377 8159 1411
rect 3341 1309 3375 1343
rect 5365 1309 5399 1343
rect 5549 1309 5583 1343
rect 5825 1309 5859 1343
rect 5917 1309 5951 1343
rect 6745 1309 6779 1343
rect 6837 1309 6871 1343
rect 7941 1309 7975 1343
rect 8309 1309 8343 1343
rect 8861 1309 8895 1343
rect 9505 1309 9539 1343
rect 8953 1241 8987 1275
rect 7481 1173 7515 1207
rect 7757 1173 7791 1207
<< metal1 >>
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4890 11540 4896 11552
rect 4212 11512 4896 11540
rect 4212 11500 4218 11512
rect 4890 11500 4896 11512
rect 4948 11540 4954 11552
rect 6362 11540 6368 11552
rect 4948 11512 6368 11540
rect 4948 11500 4954 11512
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 2372 11308 3893 11336
rect 2372 11296 2378 11308
rect 3881 11305 3893 11308
rect 3927 11336 3939 11339
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3927 11308 4077 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 3602 11268 3608 11280
rect 1912 11240 3608 11268
rect 1912 11228 1918 11240
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 3326 11200 3332 11212
rect 2700 11172 3332 11200
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2314 11132 2320 11144
rect 2271 11104 2320 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2700 11141 2728 11172
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 4080 11200 4108 11299
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 5592 11308 5917 11336
rect 5592 11296 5598 11308
rect 5905 11305 5917 11308
rect 5951 11336 5963 11339
rect 5994 11336 6000 11348
rect 5951 11308 6000 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6362 11336 6368 11348
rect 6323 11308 6368 11336
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11336 7987 11339
rect 8202 11336 8208 11348
rect 7975 11308 8208 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 4430 11268 4436 11280
rect 4391 11240 4436 11268
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 4522 11228 4528 11280
rect 4580 11268 4586 11280
rect 9125 11271 9183 11277
rect 4580 11240 8248 11268
rect 4580 11228 4586 11240
rect 4338 11200 4344 11212
rect 4080 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11200 4402 11212
rect 4396 11172 4568 11200
rect 4396 11160 4402 11172
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2915 11104 3157 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 3145 11095 3203 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4540 11141 4568 11172
rect 4982 11160 4988 11212
rect 5040 11200 5046 11212
rect 5534 11200 5540 11212
rect 5040 11172 5540 11200
rect 5040 11160 5046 11172
rect 5534 11160 5540 11172
rect 5592 11200 5598 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5592 11172 5733 11200
rect 5592 11160 5598 11172
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 5721 11163 5779 11169
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7064 11172 8125 11200
rect 7064 11160 7070 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 4939 11104 5641 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7469 11135 7527 11141
rect 7469 11132 7481 11135
rect 7156 11104 7481 11132
rect 7156 11092 7162 11104
rect 7469 11101 7481 11104
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7708 11104 7757 11132
rect 7708 11092 7714 11104
rect 7745 11101 7757 11104
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8220 11132 8248 11240
rect 9125 11237 9137 11271
rect 9171 11268 9183 11271
rect 9493 11271 9551 11277
rect 9493 11268 9505 11271
rect 9171 11240 9505 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9493 11237 9505 11240
rect 9539 11268 9551 11271
rect 13814 11268 13820 11280
rect 9539 11240 13820 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 8067 11104 8248 11132
rect 8573 11135 8631 11141
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 9490 11132 9496 11144
rect 8619 11104 9496 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 1452 11036 2513 11064
rect 1452 11024 1458 11036
rect 2501 11033 2513 11036
rect 2547 11064 2559 11067
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2547 11036 2973 11064
rect 2547 11033 2559 11036
rect 2501 11027 2559 11033
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 4798 11064 4804 11076
rect 4755 11036 4804 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4798 11024 4804 11036
rect 4856 11064 4862 11076
rect 4856 11036 4936 11064
rect 4856 11024 4862 11036
rect 2038 10996 2044 11008
rect 1999 10968 2044 10996
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2409 10999 2467 11005
rect 2409 10965 2421 10999
rect 2455 10996 2467 10999
rect 2590 10996 2596 11008
rect 2455 10968 2596 10996
rect 2455 10965 2467 10968
rect 2409 10959 2467 10965
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 3329 10999 3387 11005
rect 3329 10965 3341 10999
rect 3375 10996 3387 10999
rect 3510 10996 3516 11008
rect 3375 10968 3516 10996
rect 3375 10965 3387 10968
rect 3329 10959 3387 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 4908 10996 4936 11036
rect 4982 11024 4988 11076
rect 5040 11064 5046 11076
rect 5169 11067 5227 11073
rect 5040 11036 5085 11064
rect 5040 11024 5046 11036
rect 5169 11033 5181 11067
rect 5215 11033 5227 11067
rect 5169 11027 5227 11033
rect 5353 11067 5411 11073
rect 5353 11033 5365 11067
rect 5399 11064 5411 11067
rect 6546 11064 6552 11076
rect 5399 11036 6552 11064
rect 5399 11033 5411 11036
rect 5353 11027 5411 11033
rect 5184 10996 5212 11027
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 6822 11064 6828 11076
rect 6783 11036 6828 11064
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 6972 11036 7017 11064
rect 6972 11024 6978 11036
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7248 11036 7573 11064
rect 7248 11024 7254 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 7561 11027 7619 11033
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 8352 11036 8493 11064
rect 8352 11024 8358 11036
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8757 11067 8815 11073
rect 8757 11064 8769 11067
rect 8481 11027 8539 11033
rect 8588 11036 8769 11064
rect 5442 10996 5448 11008
rect 3660 10968 3705 10996
rect 4908 10968 5212 10996
rect 5403 10968 5448 10996
rect 3660 10956 3666 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 6178 10996 6184 11008
rect 5868 10968 6184 10996
rect 5868 10956 5874 10968
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 6932 10996 6960 11024
rect 7101 10999 7159 11005
rect 7101 10996 7113 10999
rect 6696 10968 7113 10996
rect 6696 10956 6702 10968
rect 7101 10965 7113 10968
rect 7147 10996 7159 10999
rect 7285 10999 7343 11005
rect 7285 10996 7297 10999
rect 7147 10968 7297 10996
rect 7147 10965 7159 10968
rect 7101 10959 7159 10965
rect 7285 10965 7297 10968
rect 7331 10996 7343 10999
rect 7650 10996 7656 11008
rect 7331 10968 7656 10996
rect 7331 10965 7343 10968
rect 7285 10959 7343 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8588 10996 8616 11036
rect 8757 11033 8769 11036
rect 8803 11033 8815 11067
rect 8757 11027 8815 11033
rect 9214 10996 9220 11008
rect 8076 10968 8616 10996
rect 9175 10968 9220 10996
rect 8076 10956 8082 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 1394 10792 1400 10804
rect 1355 10764 1400 10792
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4893 10795 4951 10801
rect 4893 10792 4905 10795
rect 4304 10764 4905 10792
rect 4304 10752 4310 10764
rect 4893 10761 4905 10764
rect 4939 10761 4951 10795
rect 4893 10755 4951 10761
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 5040 10764 5089 10792
rect 5040 10752 5046 10764
rect 5077 10761 5089 10764
rect 5123 10761 5135 10795
rect 5810 10792 5816 10804
rect 5077 10755 5135 10761
rect 5276 10764 5816 10792
rect 5276 10736 5304 10764
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 7466 10792 7472 10804
rect 5951 10764 7472 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 7650 10792 7656 10804
rect 7607 10764 7656 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 8110 10792 8116 10804
rect 7883 10764 8116 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9490 10792 9496 10804
rect 9451 10764 9496 10792
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 2590 10684 2596 10736
rect 2648 10684 2654 10736
rect 5258 10684 5264 10736
rect 5316 10684 5322 10736
rect 7098 10724 7104 10736
rect 7059 10696 7104 10724
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7432 10696 8340 10724
rect 7432 10684 7438 10696
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2038 10656 2044 10668
rect 1903 10628 2044 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3568 10628 3709 10656
rect 3568 10616 3574 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4396 10628 4445 10656
rect 4396 10616 4402 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 5450 10657 5508 10663
rect 5450 10623 5462 10657
rect 5496 10654 5508 10657
rect 5626 10656 5632 10668
rect 5552 10654 5632 10656
rect 5496 10628 5632 10654
rect 5496 10626 5580 10628
rect 5496 10623 5508 10626
rect 5450 10617 5508 10623
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6178 10616 6184 10668
rect 6236 10665 6242 10668
rect 6236 10656 6244 10665
rect 6914 10656 6920 10668
rect 6236 10628 6281 10656
rect 6875 10628 6920 10656
rect 6236 10619 6244 10628
rect 6236 10616 6242 10619
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7282 10656 7288 10668
rect 7239 10628 7288 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 8312 10665 8340 10696
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7392 10628 7665 10656
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2406 10588 2412 10600
rect 2271 10560 2412 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5258 10588 5264 10600
rect 4672 10560 5264 10588
rect 4672 10548 4678 10560
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 7392 10588 7420 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 8297 10619 8355 10625
rect 6604 10560 7420 10588
rect 6604 10548 6610 10560
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7944 10588 7972 10619
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 8386 10588 8392 10600
rect 7524 10560 7972 10588
rect 8036 10560 8392 10588
rect 7524 10548 7530 10560
rect 4261 10523 4319 10529
rect 4261 10489 4273 10523
rect 4307 10520 4319 10523
rect 7377 10523 7435 10529
rect 4307 10492 7328 10520
rect 4307 10489 4319 10492
rect 4261 10483 4319 10489
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 2222 10452 2228 10464
rect 1719 10424 2228 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 4706 10452 4712 10464
rect 4619 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10452 4770 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 4764 10424 5733 10452
rect 4764 10412 4770 10424
rect 5721 10421 5733 10424
rect 5767 10452 5779 10455
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5767 10424 6285 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6273 10415 6331 10421
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 6730 10452 6736 10464
rect 6687 10424 6736 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7300 10452 7328 10492
rect 7377 10489 7389 10523
rect 7423 10520 7435 10523
rect 8036 10520 8064 10560
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 7423 10492 8064 10520
rect 8113 10523 8171 10529
rect 7423 10489 7435 10492
rect 7377 10483 7435 10489
rect 8113 10489 8125 10523
rect 8159 10520 8171 10523
rect 13814 10520 13820 10532
rect 8159 10492 13820 10520
rect 8159 10489 8171 10492
rect 8113 10483 8171 10489
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 8018 10452 8024 10464
rect 7300 10424 8024 10452
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8662 10452 8668 10464
rect 8623 10424 8668 10452
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 2464 10220 2697 10248
rect 2464 10208 2470 10220
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 2685 10211 2743 10217
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 3283 10220 3893 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3881 10217 3893 10220
rect 3927 10248 3939 10251
rect 4154 10248 4160 10260
rect 3927 10220 4160 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4154 10208 4160 10220
rect 4212 10248 4218 10260
rect 4706 10248 4712 10260
rect 4212 10220 4712 10248
rect 4212 10208 4218 10220
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 6914 10248 6920 10260
rect 5552 10220 6920 10248
rect 1578 10140 1584 10192
rect 1636 10180 1642 10192
rect 5552 10189 5580 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 13814 10248 13820 10260
rect 8536 10220 13820 10248
rect 8536 10208 8542 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 5537 10183 5595 10189
rect 5537 10180 5549 10183
rect 1636 10152 5549 10180
rect 1636 10140 1642 10152
rect 5537 10149 5549 10152
rect 5583 10149 5595 10183
rect 5537 10143 5595 10149
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 8662 10180 8668 10192
rect 7616 10152 8668 10180
rect 7616 10140 7622 10152
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 1452 10084 2176 10112
rect 1452 10072 1458 10084
rect 1305 10047 1363 10053
rect 1305 10013 1317 10047
rect 1351 10044 1363 10047
rect 1762 10044 1768 10056
rect 1351 10016 1768 10044
rect 1351 10013 1363 10016
rect 1305 10007 1363 10013
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 1995 10016 2053 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 2148 10044 2176 10084
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 2869 10115 2927 10121
rect 2869 10112 2881 10115
rect 2372 10084 2881 10112
rect 2372 10072 2378 10084
rect 2869 10081 2881 10084
rect 2915 10081 2927 10115
rect 2869 10075 2927 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6822 10112 6828 10124
rect 6503 10084 6828 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 8386 10112 8392 10124
rect 7944 10084 8392 10112
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 2148 10016 3341 10044
rect 2041 10007 2099 10013
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3329 10007 3387 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 7944 10053 7972 10084
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 7929 10007 7987 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3620 9976 3648 10004
rect 3016 9948 3648 9976
rect 4249 9979 4307 9985
rect 3016 9936 3022 9948
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 4890 9976 4896 9988
rect 4295 9948 4896 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 8444 9948 8769 9976
rect 8444 9936 8450 9948
rect 8757 9945 8769 9948
rect 8803 9945 8815 9979
rect 8757 9939 8815 9945
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3844 9880 4077 9908
rect 3844 9868 3850 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 7282 9908 7288 9920
rect 6604 9880 7288 9908
rect 6604 9868 6610 9880
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 8493 9911 8551 9917
rect 8493 9877 8505 9911
rect 8539 9908 8551 9911
rect 8662 9908 8668 9920
rect 8539 9880 8668 9908
rect 8539 9877 8551 9880
rect 8493 9871 8551 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6144 9676 6745 9704
rect 6144 9664 6150 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 7098 9704 7104 9716
rect 6733 9667 6791 9673
rect 6932 9676 7104 9704
rect 4430 9596 4436 9648
rect 4488 9596 4494 9648
rect 6178 9636 6184 9648
rect 5276 9608 5672 9636
rect 6139 9608 6184 9636
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5276 9568 5304 9608
rect 4856 9540 5304 9568
rect 5353 9571 5411 9577
rect 4856 9528 4862 9540
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5442 9568 5448 9580
rect 5399 9540 5448 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5644 9568 5672 9608
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6546 9636 6552 9648
rect 6507 9608 6552 9636
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 6932 9636 6960 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8168 9676 8524 9704
rect 8168 9664 8174 9676
rect 6840 9608 6960 9636
rect 6840 9577 6868 9608
rect 8202 9596 8208 9648
rect 8260 9596 8266 9648
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5644 9540 6377 9568
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7190 9568 7196 9580
rect 6963 9540 7196 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8496 9568 8524 9676
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8496 9540 8769 9568
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 1305 9503 1363 9509
rect 1305 9469 1317 9503
rect 1351 9500 1363 9503
rect 1762 9500 1768 9512
rect 1351 9472 1768 9500
rect 1351 9469 1363 9472
rect 1305 9463 1363 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3142 9500 3148 9512
rect 3099 9472 3148 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4062 9500 4068 9512
rect 3927 9472 4068 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9500 7343 9503
rect 7558 9500 7564 9512
rect 7331 9472 7564 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 1394 9392 1400 9444
rect 1452 9432 1458 9444
rect 5917 9435 5975 9441
rect 1452 9404 1808 9432
rect 1452 9392 1458 9404
rect 1780 9364 1808 9404
rect 3252 9404 3556 9432
rect 2795 9367 2853 9373
rect 2795 9364 2807 9367
rect 1780 9336 2807 9364
rect 2795 9333 2807 9336
rect 2841 9364 2853 9367
rect 3252 9364 3280 9404
rect 3418 9364 3424 9376
rect 2841 9336 3280 9364
rect 3379 9336 3424 9364
rect 2841 9333 2853 9336
rect 2795 9327 2853 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3528 9364 3556 9404
rect 5917 9401 5929 9435
rect 5963 9432 5975 9435
rect 5963 9404 7052 9432
rect 5963 9401 5975 9404
rect 5917 9395 5975 9401
rect 5810 9364 5816 9376
rect 3528 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7024 9364 7052 9404
rect 9030 9364 9036 9376
rect 7024 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9321 9367 9379 9373
rect 9321 9333 9333 9367
rect 9367 9364 9379 9367
rect 9582 9364 9588 9376
rect 9367 9336 9588 9364
rect 9367 9333 9379 9336
rect 9321 9327 9379 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 3053 9163 3111 9169
rect 3053 9129 3065 9163
rect 3099 9160 3111 9163
rect 3234 9160 3240 9172
rect 3099 9132 3240 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3973 9163 4031 9169
rect 3973 9160 3985 9163
rect 3568 9132 3985 9160
rect 3568 9120 3574 9132
rect 3973 9129 3985 9132
rect 4019 9129 4031 9163
rect 4154 9160 4160 9172
rect 4115 9132 4160 9160
rect 3973 9123 4031 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4890 9160 4896 9172
rect 4851 9132 4896 9160
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9129 5503 9163
rect 6638 9160 6644 9172
rect 5445 9123 5503 9129
rect 6196 9132 6644 9160
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 1636 9064 2774 9092
rect 1636 9052 1642 9064
rect 2746 9024 2774 9064
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 5460 9092 5488 9123
rect 6196 9104 6224 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7190 9160 7196 9172
rect 6880 9132 7196 9160
rect 6880 9120 6886 9132
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 4764 9064 5488 9092
rect 5721 9095 5779 9101
rect 4764 9052 4770 9064
rect 5721 9061 5733 9095
rect 5767 9092 5779 9095
rect 6178 9092 6184 9104
rect 5767 9064 6184 9092
rect 5767 9061 5779 9064
rect 5721 9055 5779 9061
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 8754 9052 8760 9104
rect 8812 9052 8818 9104
rect 3050 9024 3056 9036
rect 2746 8996 3056 9024
rect 3050 8984 3056 8996
rect 3108 9024 3114 9036
rect 4246 9024 4252 9036
rect 3108 8996 4252 9024
rect 3108 8984 3114 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 5534 9024 5540 9036
rect 4356 8996 5540 9024
rect 1302 8956 1308 8968
rect 1263 8928 1308 8956
rect 1302 8916 1308 8928
rect 1360 8916 1366 8968
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1995 8928 2053 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 2280 8928 3433 8956
rect 2280 8916 2286 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3786 8956 3792 8968
rect 3747 8928 3792 8956
rect 3421 8919 3479 8925
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 2406 8888 2412 8900
rect 1544 8860 2412 8888
rect 1544 8848 1550 8860
rect 2406 8848 2412 8860
rect 2464 8848 2470 8900
rect 2777 8891 2835 8897
rect 2777 8857 2789 8891
rect 2823 8888 2835 8891
rect 2866 8888 2872 8900
rect 2823 8860 2872 8888
rect 2823 8857 2835 8860
rect 2777 8851 2835 8857
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 2961 8891 3019 8897
rect 2961 8857 2973 8891
rect 3007 8888 3019 8891
rect 3234 8888 3240 8900
rect 3007 8860 3240 8888
rect 3007 8857 3019 8860
rect 2961 8851 3019 8857
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 3436 8888 3464 8919
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4356 8965 4384 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 7466 9024 7472 9036
rect 5828 8996 7472 9024
rect 5828 8965 5856 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7708 8996 7941 9024
rect 7708 8984 7714 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 8772 9024 8800 9052
rect 13630 9024 13636 9036
rect 7929 8987 7987 8993
rect 8312 8996 13636 9024
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 4341 8919 4399 8925
rect 4540 8928 5089 8956
rect 3896 8888 3924 8919
rect 3436 8860 3924 8888
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4540 8888 4568 8928
rect 5077 8925 5089 8928
rect 5123 8956 5135 8959
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5123 8928 5825 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 4028 8860 4568 8888
rect 4617 8891 4675 8897
rect 4028 8848 4034 8860
rect 4617 8857 4629 8891
rect 4663 8857 4675 8891
rect 4617 8851 4675 8857
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2280 8792 2697 8820
rect 2280 8780 2286 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3108 8792 3341 8820
rect 3108 8780 3114 8792
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3602 8820 3608 8832
rect 3563 8792 3608 8820
rect 3329 8783 3387 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 4632 8820 4660 8851
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5169 8891 5227 8897
rect 5169 8888 5181 8891
rect 5040 8860 5181 8888
rect 5040 8848 5046 8860
rect 5169 8857 5181 8860
rect 5215 8857 5227 8891
rect 5169 8851 5227 8857
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5534 8888 5540 8900
rect 5399 8860 5540 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 5997 8891 6055 8897
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 6086 8888 6092 8900
rect 6043 8860 6092 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 5442 8820 5448 8832
rect 4632 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 6196 8820 6224 8919
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8312 8965 8340 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 7616 8928 8309 8956
rect 7616 8916 7622 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 8846 8956 8852 8968
rect 8803 8928 8852 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8888 6515 8891
rect 6546 8888 6552 8900
rect 6503 8860 6552 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 7760 8860 8125 8888
rect 7374 8820 7380 8832
rect 5684 8792 7380 8820
rect 5684 8780 5690 8792
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 7760 8820 7788 8860
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 8938 8888 8944 8900
rect 8260 8860 8944 8888
rect 8260 8848 8266 8860
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 7524 8792 7788 8820
rect 8481 8823 8539 8829
rect 7524 8780 7530 8792
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 13722 8820 13728 8832
rect 8527 8792 13728 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 1394 8616 1400 8628
rect 1355 8588 1400 8616
rect 1394 8576 1400 8588
rect 1452 8576 1458 8628
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 3050 8616 3056 8628
rect 1872 8588 3056 8616
rect 1872 8489 1900 8588
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 5828 8588 6469 8616
rect 3602 8548 3608 8560
rect 3358 8520 3608 8548
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4304 8520 4568 8548
rect 4304 8508 4310 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 1857 8443 1915 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3476 8452 3709 8480
rect 3476 8440 3482 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 4430 8480 4436 8492
rect 4391 8452 4436 8480
rect 3697 8443 3755 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4540 8480 4568 8520
rect 4798 8508 4804 8560
rect 4856 8548 4862 8560
rect 5828 8557 5856 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 6917 8619 6975 8625
rect 6917 8616 6929 8619
rect 6880 8588 6929 8616
rect 6880 8576 6886 8588
rect 6917 8585 6929 8588
rect 6963 8585 6975 8619
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 6917 8579 6975 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 13538 8616 13544 8628
rect 12406 8588 13544 8616
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 4856 8520 5365 8548
rect 4856 8508 4862 8520
rect 5353 8517 5365 8520
rect 5399 8548 5411 8551
rect 5813 8551 5871 8557
rect 5813 8548 5825 8551
rect 5399 8520 5825 8548
rect 5399 8517 5411 8520
rect 5353 8511 5411 8517
rect 5813 8517 5825 8520
rect 5859 8517 5871 8551
rect 5813 8511 5871 8517
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4540 8452 5181 8480
rect 4816 8424 4844 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5316 8452 5641 8480
rect 5316 8440 5322 8452
rect 5629 8449 5641 8452
rect 5675 8480 5687 8483
rect 5902 8480 5908 8492
rect 5675 8452 5908 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6178 8480 6184 8492
rect 6139 8452 6184 8480
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6638 8480 6644 8492
rect 6599 8452 6644 8480
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 2866 8412 2872 8424
rect 1811 8384 2872 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 4798 8372 4804 8424
rect 4856 8372 4862 8424
rect 6748 8412 6776 8443
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6880 8452 7021 8480
rect 6880 8440 6886 8452
rect 7009 8449 7021 8452
rect 7055 8480 7067 8483
rect 7098 8480 7104 8492
rect 7055 8452 7104 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7374 8480 7380 8492
rect 7335 8452 7380 8480
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 8996 8452 9321 8480
rect 8996 8440 9002 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 7282 8412 7288 8424
rect 6748 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7650 8412 7656 8424
rect 7611 8384 7656 8412
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 12406 8412 12434 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 8680 8384 12434 8412
rect 4261 8347 4319 8353
rect 4261 8313 4273 8347
rect 4307 8344 4319 8347
rect 4890 8344 4896 8356
rect 4307 8316 4896 8344
rect 4307 8313 4319 8316
rect 4261 8307 4319 8313
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 5534 8344 5540 8356
rect 5495 8316 5540 8344
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 5868 8316 7512 8344
rect 5868 8304 5874 8316
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 5077 8279 5135 8285
rect 5077 8276 5089 8279
rect 4672 8248 5089 8276
rect 4672 8236 4678 8248
rect 5077 8245 5089 8248
rect 5123 8245 5135 8279
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5077 8239 5135 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6365 8279 6423 8285
rect 6365 8245 6377 8279
rect 6411 8276 6423 8279
rect 6546 8276 6552 8288
rect 6411 8248 6552 8276
rect 6411 8245 6423 8248
rect 6365 8239 6423 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6730 8236 6736 8288
rect 6788 8276 6794 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 6788 8248 7205 8276
rect 6788 8236 6794 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 7484 8276 7512 8316
rect 8680 8276 8708 8384
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 8812 8316 9137 8344
rect 8812 8304 8818 8316
rect 9125 8313 9137 8316
rect 9171 8313 9183 8347
rect 9125 8307 9183 8313
rect 7484 8248 8708 8276
rect 7193 8239 7251 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4430 8072 4436 8084
rect 4295 8044 4436 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 5261 8075 5319 8081
rect 5261 8072 5273 8075
rect 4847 8044 5273 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 5261 8041 5273 8044
rect 5307 8072 5319 8075
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 5307 8044 6285 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 8570 8072 8576 8084
rect 6503 8044 8576 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 3050 7964 3056 8016
rect 3108 8004 3114 8016
rect 5626 8004 5632 8016
rect 3108 7976 5632 8004
rect 3108 7964 3114 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 1452 7908 1624 7936
rect 1452 7896 1458 7908
rect 1486 7868 1492 7880
rect 1447 7840 1492 7868
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 1596 7877 1624 7908
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 2924 7908 3341 7936
rect 2924 7896 2930 7908
rect 3329 7905 3341 7908
rect 3375 7905 3387 7939
rect 6178 7936 6184 7948
rect 3329 7899 3387 7905
rect 4080 7908 6184 7936
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 3344 7868 3372 7899
rect 3605 7871 3663 7877
rect 3605 7868 3617 7871
rect 3344 7840 3617 7868
rect 1581 7831 1639 7837
rect 3605 7837 3617 7840
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 1820 7772 1869 7800
rect 1820 7760 1826 7772
rect 1857 7769 1869 7772
rect 1903 7769 1915 7803
rect 3142 7800 3148 7812
rect 3055 7772 3148 7800
rect 1857 7763 1915 7769
rect 3142 7760 3148 7772
rect 3200 7800 3206 7812
rect 4080 7800 4108 7908
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6288 7936 6316 8035
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9364 8044 9413 8072
rect 9364 8032 9370 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 7098 8004 7104 8016
rect 6604 7976 7104 8004
rect 6604 7964 6610 7976
rect 7098 7964 7104 7976
rect 7156 7964 7162 8016
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 8018 8004 8024 8016
rect 7800 7976 8024 8004
rect 7800 7964 7806 7976
rect 8018 7964 8024 7976
rect 8076 8004 8082 8016
rect 8076 7976 8248 8004
rect 8076 7964 8082 7976
rect 6730 7936 6736 7948
rect 6288 7908 6736 7936
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4856 7840 4905 7868
rect 4856 7828 4862 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5258 7868 5264 7880
rect 5040 7840 5264 7868
rect 5040 7828 5046 7840
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5994 7868 6000 7880
rect 5955 7840 6000 7868
rect 5994 7828 6000 7840
rect 6052 7868 6058 7880
rect 6638 7868 6644 7880
rect 6052 7840 6500 7868
rect 6599 7840 6644 7868
rect 6052 7828 6058 7840
rect 3200 7772 4108 7800
rect 5813 7803 5871 7809
rect 3200 7760 3206 7772
rect 5813 7769 5825 7803
rect 5859 7800 5871 7803
rect 6178 7800 6184 7812
rect 5859 7772 6184 7800
rect 5859 7769 5871 7772
rect 5813 7763 5871 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6472 7800 6500 7840
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7524 7840 7757 7868
rect 7524 7828 7530 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8220 7877 8248 7976
rect 8938 7936 8944 7948
rect 8404 7908 8944 7936
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7892 7840 8033 7868
rect 7892 7828 7898 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 6472 7772 7389 7800
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7558 7800 7564 7812
rect 7519 7772 7564 7800
rect 7377 7763 7435 7769
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 3418 7732 3424 7744
rect 1443 7704 3424 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 4396 7704 4445 7732
rect 4396 7692 4402 7704
rect 4433 7701 4445 7704
rect 4479 7701 4491 7735
rect 4433 7695 4491 7701
rect 5445 7735 5503 7741
rect 5445 7701 5457 7735
rect 5491 7732 5503 7735
rect 6362 7732 6368 7744
rect 5491 7704 6368 7732
rect 5491 7701 5503 7704
rect 5445 7695 5503 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7156 7704 7297 7732
rect 7156 7692 7162 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7392 7732 7420 7763
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 8404 7800 8432 7908
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8536 7840 8769 7868
rect 8536 7828 8542 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8312 7772 8432 7800
rect 8573 7803 8631 7809
rect 7834 7732 7840 7744
rect 7392 7704 7840 7732
rect 7285 7695 7343 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8312 7741 8340 7772
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 9214 7800 9220 7812
rect 8619 7772 9220 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 7975 7704 8309 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8297 7695 8355 7701
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7732 8447 7735
rect 8478 7732 8484 7744
rect 8435 7704 8484 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 1302 7528 1308 7540
rect 1263 7500 1308 7528
rect 1302 7488 1308 7500
rect 1360 7488 1366 7540
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1544 7500 3280 7528
rect 1544 7488 1550 7500
rect 2777 7463 2835 7469
rect 2777 7429 2789 7463
rect 2823 7460 2835 7463
rect 2866 7460 2872 7472
rect 2823 7432 2872 7460
rect 2823 7429 2835 7432
rect 2777 7423 2835 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3252 7401 3280 7500
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 4614 7528 4620 7540
rect 3936 7500 4620 7528
rect 3936 7488 3942 7500
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5913 7531 5971 7537
rect 5913 7497 5925 7531
rect 5959 7528 5971 7531
rect 5959 7500 8340 7528
rect 5959 7497 5971 7500
rect 5913 7491 5971 7497
rect 5994 7460 6000 7472
rect 5014 7432 6000 7460
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 7650 7420 7656 7472
rect 7708 7420 7714 7472
rect 8312 7460 8340 7500
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8904 7500 9137 7528
rect 8904 7488 8910 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 8478 7460 8484 7472
rect 8312 7432 8484 7460
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 3237 7395 3295 7401
rect 3108 7364 3153 7392
rect 3108 7352 3114 7364
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 3068 7188 3096 7352
rect 3252 7324 3280 7355
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3476 7364 3525 7392
rect 3476 7352 3482 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 5350 7392 5356 7404
rect 3513 7355 3571 7361
rect 3620 7364 4016 7392
rect 5311 7364 5356 7392
rect 3620 7324 3648 7364
rect 3878 7324 3884 7336
rect 3252 7296 3648 7324
rect 3839 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 3988 7324 4016 7364
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5592 7364 6377 7392
rect 5592 7352 5598 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 7006 7392 7012 7404
rect 6595 7364 7012 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 4522 7324 4528 7336
rect 3988 7296 4528 7324
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7324 6975 7327
rect 7190 7324 7196 7336
rect 6963 7296 7196 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 5592 7228 6193 7256
rect 5592 7216 5598 7228
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 9401 7259 9459 7265
rect 9401 7256 9413 7259
rect 7892 7228 9413 7256
rect 7892 7216 7898 7228
rect 9401 7225 9413 7228
rect 9447 7225 9459 7259
rect 9401 7219 9459 7225
rect 3326 7188 3332 7200
rect 1452 7160 3096 7188
rect 3287 7160 3332 7188
rect 1452 7148 1458 7160
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 8846 7188 8852 7200
rect 8619 7160 8852 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 8953 7191 9011 7197
rect 8953 7157 8965 7191
rect 8999 7188 9011 7191
rect 9122 7188 9128 7200
rect 8999 7160 9128 7188
rect 8999 7157 9011 7160
rect 8953 7151 9011 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1302 6944 1308 6996
rect 1360 6984 1366 6996
rect 1746 6987 1804 6993
rect 1746 6984 1758 6987
rect 1360 6956 1758 6984
rect 1360 6944 1366 6956
rect 1746 6953 1758 6956
rect 1792 6953 1804 6987
rect 1746 6947 1804 6953
rect 7395 6987 7453 6993
rect 7395 6953 7407 6987
rect 7441 6984 7453 6987
rect 8754 6984 8760 6996
rect 7441 6956 8760 6984
rect 7441 6953 7453 6956
rect 7395 6947 7453 6953
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6984 9094 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9088 6956 9413 6984
rect 9088 6944 9094 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9401 6947 9459 6953
rect 8294 6916 8300 6928
rect 8140 6888 8300 6916
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1489 6851 1547 6857
rect 1489 6848 1501 6851
rect 1452 6820 1501 6848
rect 1452 6808 1458 6820
rect 1489 6817 1501 6820
rect 1535 6817 1547 6851
rect 1489 6811 1547 6817
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 1820 6820 3004 6848
rect 1820 6808 1826 6820
rect 1397 6715 1455 6721
rect 1397 6681 1409 6715
rect 1443 6712 1455 6715
rect 1670 6712 1676 6724
rect 1443 6684 1676 6712
rect 1443 6681 1455 6684
rect 1397 6675 1455 6681
rect 1670 6672 1676 6684
rect 1728 6672 1734 6724
rect 2976 6712 3004 6820
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4120 6820 4997 6848
rect 4120 6808 4126 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 6638 6848 6644 6860
rect 5123 6820 6644 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7432 6820 7665 6848
rect 7432 6808 7438 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 3605 6783 3663 6789
rect 3605 6780 3617 6783
rect 3252 6752 3617 6780
rect 3142 6712 3148 6724
rect 2976 6698 3148 6712
rect 2990 6684 3148 6698
rect 3142 6672 3148 6684
rect 3200 6672 3206 6724
rect 3252 6656 3280 6752
rect 3605 6749 3617 6752
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4295 6752 4353 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5767 6752 5948 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 5920 6653 5948 6752
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8140 6780 8168 6888
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 13722 6848 13728 6860
rect 8251 6820 13728 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 8067 6752 8168 6780
rect 8297 6783 8355 6789
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8297 6743 8355 6749
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8312 6712 8340 6743
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 8168 6684 8340 6712
rect 8168 6672 8174 6684
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8772 6712 8800 6743
rect 8536 6684 8800 6712
rect 8536 6672 8542 6684
rect 5905 6647 5963 6653
rect 5905 6613 5917 6647
rect 5951 6644 5963 6647
rect 6546 6644 6552 6656
rect 5951 6616 6552 6644
rect 5951 6613 5963 6616
rect 5905 6607 5963 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 7374 6644 7380 6656
rect 6788 6616 7380 6644
rect 6788 6604 6794 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9306 6644 9312 6656
rect 9263 6616 9312 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1443 6412 1593 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 1581 6409 1593 6412
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 2464 6412 3249 6440
rect 2464 6400 2470 6412
rect 3237 6409 3249 6412
rect 3283 6440 3295 6443
rect 4982 6440 4988 6452
rect 3283 6412 4988 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7834 6440 7840 6452
rect 7248 6412 7840 6440
rect 7248 6400 7254 6412
rect 7834 6400 7840 6412
rect 7892 6440 7898 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 7892 6412 8248 6440
rect 7892 6400 7898 6412
rect 4154 6332 4160 6384
rect 4212 6332 4218 6384
rect 7926 6372 7932 6384
rect 7887 6344 7932 6372
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8220 6381 8248 6412
rect 8404 6412 9413 6440
rect 8205 6375 8263 6381
rect 8205 6341 8217 6375
rect 8251 6341 8263 6375
rect 8205 6335 8263 6341
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6273 2467 6307
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 2409 6267 2467 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2424 6236 2452 6267
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5534 6304 5540 6316
rect 5215 6276 5540 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 5776 6276 8033 6304
rect 5776 6264 5782 6276
rect 8021 6273 8033 6276
rect 8067 6304 8079 6307
rect 8404 6304 8432 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 8067 6276 8432 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8754 6304 8760 6316
rect 8536 6276 8581 6304
rect 8715 6276 8760 6304
rect 8536 6264 8542 6276
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8904 6276 8953 6304
rect 8904 6264 8910 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9582 6304 9588 6316
rect 9355 6276 9588 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 1719 6208 2452 6236
rect 3053 6239 3111 6245
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3099 6208 3709 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 6144 6208 6193 6236
rect 6144 6196 6150 6208
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8168 6208 8585 6236
rect 8168 6196 8174 6208
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 5733 6171 5791 6177
rect 5733 6137 5745 6171
rect 5779 6168 5791 6171
rect 8202 6168 8208 6180
rect 5779 6140 8208 6168
rect 5779 6137 5791 6140
rect 5733 6131 5791 6137
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 8389 6171 8447 6177
rect 8389 6137 8401 6171
rect 8435 6168 8447 6171
rect 9490 6168 9496 6180
rect 8435 6140 9496 6168
rect 8435 6137 8447 6140
rect 8389 6131 8447 6137
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 4856 6072 5917 6100
rect 4856 6060 4862 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 8110 6100 8116 6112
rect 7064 6072 8116 6100
rect 7064 6060 7070 6072
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1489 5899 1547 5905
rect 1489 5865 1501 5899
rect 1535 5896 1547 5899
rect 1670 5896 1676 5908
rect 1535 5868 1676 5896
rect 1535 5865 1547 5868
rect 1489 5859 1547 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 2464 5868 4261 5896
rect 2464 5856 2470 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 7432 5868 8309 5896
rect 7432 5856 7438 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8628 5868 8861 5896
rect 8628 5856 8634 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 8478 5828 8484 5840
rect 5552 5800 8484 5828
rect 1305 5763 1363 5769
rect 1305 5729 1317 5763
rect 1351 5760 1363 5763
rect 1351 5732 5488 5760
rect 1351 5729 1363 5732
rect 1305 5723 1363 5729
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 3421 5695 3479 5701
rect 1728 5664 2070 5692
rect 1728 5652 1734 5664
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 3234 5624 3240 5636
rect 3191 5596 3240 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 3436 5624 3464 5655
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 3844 5664 4445 5692
rect 3844 5652 3850 5664
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 4798 5624 4804 5636
rect 3436 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 5460 5624 5488 5732
rect 5552 5701 5580 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8812 5800 9229 5828
rect 8812 5788 8818 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 13446 5760 13452 5772
rect 5951 5732 13452 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 5537 5655 5595 5661
rect 6012 5664 7941 5692
rect 6012 5624 6040 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 6178 5624 6184 5636
rect 5460 5596 6040 5624
rect 6139 5596 6184 5624
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 7944 5624 7972 5655
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8168 5664 8585 5692
rect 8168 5652 8174 5664
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 8573 5655 8631 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9582 5692 9588 5704
rect 9355 5664 9588 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 13814 5624 13820 5636
rect 7944 5596 13820 5624
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5556 1731 5559
rect 3694 5556 3700 5568
rect 1719 5528 3700 5556
rect 1719 5525 1731 5528
rect 1673 5519 1731 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 7834 5556 7840 5568
rect 4948 5528 7840 5556
rect 4948 5516 4954 5528
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8110 5556 8116 5568
rect 8071 5528 8116 5556
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 8904 5528 9413 5556
rect 8904 5516 8910 5528
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 3476 5324 3525 5352
rect 3476 5312 3482 5324
rect 3513 5321 3525 5324
rect 3559 5321 3571 5355
rect 3513 5315 3571 5321
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4111 5324 5212 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 3804 5284 3832 5315
rect 4154 5284 4160 5296
rect 3804 5256 4160 5284
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 5184 5293 5212 5324
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5500 5324 6469 5352
rect 5500 5312 5506 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8444 5324 8493 5352
rect 8444 5312 8450 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 8812 5324 8892 5352
rect 8812 5312 8818 5324
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5253 5227 5287
rect 7024 5284 7052 5312
rect 7024 5256 7420 5284
rect 5169 5247 5227 5253
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3200 5188 3341 5216
rect 3200 5176 3206 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 3970 5216 3976 5228
rect 3927 5188 3976 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 3620 5148 3648 5179
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4246 5148 4252 5160
rect 3620 5120 4252 5148
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4356 5148 4384 5179
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4488 5188 5089 5216
rect 4488 5176 4494 5188
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 5776 5188 7021 5216
rect 5776 5176 5782 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7392 5216 7420 5256
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 8864 5293 8892 5324
rect 8849 5287 8907 5293
rect 7524 5256 8340 5284
rect 7524 5244 7530 5256
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7392 5188 7665 5216
rect 7009 5179 7067 5185
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5216 7895 5219
rect 7926 5216 7932 5228
rect 7883 5188 7932 5216
rect 7883 5185 7895 5188
rect 7837 5179 7895 5185
rect 6086 5148 6092 5160
rect 4356 5120 6092 5148
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 7852 5148 7880 5179
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8312 5225 8340 5256
rect 8849 5253 8861 5287
rect 8895 5253 8907 5287
rect 8849 5247 8907 5253
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8720 5188 8769 5216
rect 8720 5176 8726 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8938 5216 8944 5228
rect 8899 5188 8944 5216
rect 8757 5179 8815 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9217 5179 9275 5185
rect 6196 5120 7880 5148
rect 9232 5148 9260 5179
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9232 5120 9904 5148
rect 4154 5080 4160 5092
rect 4115 5052 4160 5080
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 5902 5080 5908 5092
rect 5224 5052 5908 5080
rect 5224 5040 5230 5052
rect 5902 5040 5908 5052
rect 5960 5080 5966 5092
rect 6196 5080 6224 5120
rect 5960 5052 6224 5080
rect 7469 5083 7527 5089
rect 5960 5040 5966 5052
rect 7469 5049 7481 5083
rect 7515 5080 7527 5083
rect 9214 5080 9220 5092
rect 7515 5052 9220 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 9214 5040 9220 5052
rect 9272 5040 9278 5092
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4396 4984 4629 5012
rect 4396 4972 4402 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4764 4984 4813 5012
rect 4764 4972 4770 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 4801 4975 4859 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7374 5012 7380 5024
rect 7331 4984 7380 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7926 5012 7932 5024
rect 7887 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 8076 4984 8585 5012
rect 8076 4972 8082 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 8573 4975 8631 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 3418 4768 3424 4820
rect 3476 4808 3482 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3476 4780 3801 4808
rect 3476 4768 3482 4780
rect 3789 4777 3801 4780
rect 3835 4808 3847 4811
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3835 4780 4445 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4433 4777 4445 4780
rect 4479 4808 4491 4811
rect 4706 4808 4712 4820
rect 4479 4780 4712 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 7466 4808 7472 4820
rect 4847 4780 7472 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 8861 4811 8919 4817
rect 8861 4777 8873 4811
rect 8907 4808 8919 4811
rect 9876 4808 9904 5120
rect 13814 4808 13820 4820
rect 8907 4780 13820 4808
rect 8907 4777 8919 4780
rect 8861 4771 8919 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 3602 4700 3608 4752
rect 3660 4740 3666 4752
rect 3660 4712 4384 4740
rect 3660 4700 3666 4712
rect 4154 4672 4160 4684
rect 3620 4644 4160 4672
rect 3510 4564 3516 4616
rect 3568 4564 3574 4616
rect 3620 4613 3648 4644
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4356 4613 4384 4712
rect 4890 4700 4896 4752
rect 4948 4740 4954 4752
rect 5537 4743 5595 4749
rect 4948 4712 5396 4740
rect 4948 4700 4954 4712
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4573 3755 4607
rect 3697 4567 3755 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4387 4576 5120 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 3528 4536 3556 4564
rect 3712 4536 3740 4567
rect 3528 4508 4476 4536
rect 3513 4471 3571 4477
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 4062 4468 4068 4480
rect 3559 4440 4068 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4246 4468 4252 4480
rect 4203 4440 4252 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4448 4468 4476 4508
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 4985 4539 5043 4545
rect 4985 4536 4997 4539
rect 4580 4508 4997 4536
rect 4580 4496 4586 4508
rect 4985 4505 4997 4508
rect 5031 4505 5043 4539
rect 4985 4499 5043 4505
rect 4890 4468 4896 4480
rect 4448 4440 4896 4468
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5092 4468 5120 4576
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5368 4613 5396 4712
rect 5537 4709 5549 4743
rect 5583 4740 5595 4743
rect 5718 4740 5724 4752
rect 5583 4712 5724 4740
rect 5583 4709 5595 4712
rect 5537 4703 5595 4709
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6181 4743 6239 4749
rect 6181 4740 6193 4743
rect 6052 4712 6193 4740
rect 6052 4700 6058 4712
rect 6181 4709 6193 4712
rect 6227 4709 6239 4743
rect 6181 4703 6239 4709
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 7984 4712 9444 4740
rect 7984 4700 7990 4712
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7098 4672 7104 4684
rect 6871 4644 7104 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 9306 4672 9312 4684
rect 8312 4644 9312 4672
rect 5353 4607 5411 4613
rect 5224 4576 5269 4604
rect 5224 4564 5230 4576
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 5353 4567 5411 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6362 4604 6368 4616
rect 6323 4576 6368 4604
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 8312 4613 8340 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 8297 4607 8355 4613
rect 6512 4576 6557 4604
rect 6512 4564 6518 4576
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 8297 4567 8355 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9416 4604 9444 4712
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9416 4576 9505 4604
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4505 5779 4539
rect 5721 4499 5779 4505
rect 5736 4468 5764 4499
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 6052 4508 6101 4536
rect 6052 4496 6058 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 7958 4508 9076 4536
rect 6089 4499 6147 4505
rect 9048 4477 9076 4508
rect 5092 4440 5764 4468
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4437 9091 4471
rect 9306 4468 9312 4480
rect 9267 4440 9312 4468
rect 9033 4431 9091 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3568 4236 3801 4264
rect 3568 4224 3574 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 3789 4227 3847 4233
rect 4246 4224 4252 4276
rect 4304 4224 4310 4276
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 7469 4267 7527 4273
rect 5500 4236 6960 4264
rect 5500 4224 5506 4236
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 3605 4199 3663 4205
rect 3605 4196 3617 4199
rect 3200 4168 3617 4196
rect 3200 4156 3206 4168
rect 3605 4165 3617 4168
rect 3651 4196 3663 4199
rect 3878 4196 3884 4208
rect 3651 4168 3884 4196
rect 3651 4165 3663 4168
rect 3605 4159 3663 4165
rect 3878 4156 3884 4168
rect 3936 4156 3942 4208
rect 4264 4196 4292 4224
rect 6932 4205 6960 4236
rect 7469 4233 7481 4267
rect 7515 4233 7527 4267
rect 7469 4227 7527 4233
rect 6917 4199 6975 4205
rect 3988 4168 4292 4196
rect 5750 4168 6868 4196
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 3786 4128 3792 4140
rect 2740 4100 3792 4128
rect 2740 4088 2746 4100
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3988 4137 4016 4168
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4120 4100 4261 4128
rect 4120 4088 4126 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 6086 4128 6092 4140
rect 6047 4100 6092 4128
rect 4249 4091 4307 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6653 4131 6711 4137
rect 6653 4128 6665 4131
rect 6420 4100 6665 4128
rect 6420 4088 6426 4100
rect 6653 4097 6665 4100
rect 6699 4097 6711 4131
rect 6840 4128 6868 4168
rect 6917 4165 6929 4199
rect 6963 4165 6975 4199
rect 7484 4196 7512 4227
rect 6917 4159 6975 4165
rect 7024 4168 7512 4196
rect 7944 4168 9352 4196
rect 7024 4128 7052 4168
rect 6840 4100 7052 4128
rect 7193 4131 7251 4137
rect 6653 4091 6711 4097
rect 7193 4097 7205 4131
rect 7239 4128 7251 4131
rect 7239 4100 7420 4128
rect 7239 4097 7251 4100
rect 7193 4091 7251 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3602 4060 3608 4072
rect 3467 4032 3608 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6512 4032 7297 4060
rect 6512 4020 6518 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 3568 3964 4384 3992
rect 3568 3952 3574 3964
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4356 3924 4384 3964
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 5592 3964 7113 3992
rect 5592 3952 5598 3964
rect 7101 3961 7113 3964
rect 7147 3992 7159 3995
rect 7392 3992 7420 4100
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7524 4100 7665 4128
rect 7524 4088 7530 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 7944 4128 7972 4168
rect 8110 4128 8116 4140
rect 7800 4100 7972 4128
rect 8071 4100 8116 4128
rect 7800 4088 7806 4100
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8536 4100 9137 4128
rect 8536 4088 8542 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9324 4128 9352 4168
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9324 4100 9505 4128
rect 9217 4091 9275 4097
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 13722 4128 13728 4140
rect 9493 4091 9551 4097
rect 12406 4100 13728 4128
rect 8754 4060 8760 4072
rect 7147 3964 7420 3992
rect 7760 4032 8760 4060
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 7760 3933 7788 4032
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 9232 4060 9260 4091
rect 12406 4060 12434 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 8812 4032 12434 4060
rect 8812 4020 8818 4032
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8444 3964 9321 3992
rect 8444 3952 8450 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 4356 3896 7757 3924
rect 4157 3887 4215 3893
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 7929 3927 7987 3933
rect 7929 3893 7941 3927
rect 7975 3924 7987 3927
rect 8018 3924 8024 3936
rect 7975 3896 8024 3924
rect 7975 3893 7987 3896
rect 7929 3887 7987 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8938 3924 8944 3936
rect 8899 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3602 3720 3608 3732
rect 3563 3692 3608 3720
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 4338 3720 4344 3732
rect 4172 3692 4344 3720
rect 3421 3655 3479 3661
rect 3421 3621 3433 3655
rect 3467 3652 3479 3655
rect 4172 3652 4200 3692
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 4672 3692 6377 3720
rect 4672 3680 4678 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 9137 3723 9195 3729
rect 9137 3689 9149 3723
rect 9183 3720 9195 3723
rect 9490 3720 9496 3732
rect 9183 3692 9496 3720
rect 9183 3689 9195 3692
rect 9137 3683 9195 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 3467 3624 4200 3652
rect 3467 3621 3479 3624
rect 3421 3615 3479 3621
rect 4246 3612 4252 3664
rect 4304 3612 4310 3664
rect 4433 3655 4491 3661
rect 4433 3621 4445 3655
rect 4479 3621 4491 3655
rect 4798 3652 4804 3664
rect 4759 3624 4804 3652
rect 4433 3615 4491 3621
rect 4264 3584 4292 3612
rect 3988 3556 4292 3584
rect 4448 3584 4476 3615
rect 4798 3612 4804 3624
rect 4856 3652 4862 3664
rect 4982 3652 4988 3664
rect 4856 3624 4988 3652
rect 4856 3612 4862 3624
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 6086 3652 6092 3664
rect 5276 3624 6092 3652
rect 5276 3584 5304 3624
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 4448 3556 5304 3584
rect 5445 3587 5503 3593
rect 3988 3525 4016 3556
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 5491 3556 6745 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 3896 3448 3924 3479
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4522 3516 4528 3528
rect 4304 3488 4349 3516
rect 4483 3488 4528 3516
rect 4304 3476 4310 3488
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4890 3476 4896 3528
rect 4948 3516 4954 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 4948 3488 5181 3516
rect 4948 3476 4954 3488
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5169 3479 5227 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5684 3488 5733 3516
rect 5684 3476 5690 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 5721 3479 5779 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9306 3516 9312 3528
rect 8619 3488 9312 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 4172 3448 4200 3476
rect 4798 3448 4804 3460
rect 3896 3420 4804 3448
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 4985 3451 5043 3457
rect 4985 3417 4997 3451
rect 5031 3448 5043 3451
rect 6178 3448 6184 3460
rect 5031 3420 6184 3448
rect 5031 3417 5043 3420
rect 4985 3411 5043 3417
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 8018 3408 8024 3460
rect 8076 3408 8082 3460
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3660 3352 3801 3380
rect 3660 3340 3666 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 3789 3343 3847 3349
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4709 3383 4767 3389
rect 4709 3349 4721 3383
rect 4755 3380 4767 3383
rect 4890 3380 4896 3392
rect 4755 3352 4896 3380
rect 4755 3349 4767 3352
rect 4709 3343 4767 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5902 3340 5908 3392
rect 5960 3380 5966 3392
rect 6457 3383 6515 3389
rect 6457 3380 6469 3383
rect 5960 3352 6469 3380
rect 5960 3340 5966 3352
rect 6457 3349 6469 3352
rect 6503 3349 6515 3383
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 6457 3343 6515 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 3036 3216 9844 3238
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4120 3148 4292 3176
rect 4120 3136 4126 3148
rect 4264 3108 4292 3148
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5994 3176 6000 3188
rect 4488 3148 6000 3176
rect 4488 3136 4494 3148
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 8021 3179 8079 3185
rect 6328 3148 6684 3176
rect 6328 3136 6334 3148
rect 4264 3080 4370 3108
rect 5810 3068 5816 3120
rect 5868 3108 5874 3120
rect 6288 3108 6316 3136
rect 6546 3108 6552 3120
rect 5868 3080 6316 3108
rect 6507 3080 6552 3108
rect 5868 3068 5874 3080
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 6656 3108 6684 3148
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8294 3176 8300 3188
rect 8067 3148 8300 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9306 3136 9312 3188
rect 9364 3136 9370 3188
rect 6822 3108 6828 3120
rect 6656 3080 6828 3108
rect 6822 3068 6828 3080
rect 6880 3108 6886 3120
rect 8754 3108 8760 3120
rect 6880 3080 7038 3108
rect 8715 3080 8760 3108
rect 6880 3068 6886 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3108 8907 3111
rect 9324 3108 9352 3136
rect 8895 3080 9352 3108
rect 8895 3077 8907 3080
rect 8849 3071 8907 3077
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4948 3012 5457 3040
rect 4948 3000 4954 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3712 2944 3985 2972
rect 3712 2836 3740 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2941 6331 2975
rect 6273 2935 6331 2941
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 6288 2904 6316 2935
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7064 2944 8309 2972
rect 7064 2932 7070 2944
rect 8297 2941 8309 2944
rect 8343 2972 8355 2975
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8343 2944 8493 2972
rect 8343 2941 8355 2944
rect 8297 2935 8355 2941
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 8481 2935 8539 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 5040 2876 6316 2904
rect 5040 2864 5046 2876
rect 13814 2864 13820 2916
rect 13872 2904 13878 2916
rect 16666 2904 16672 2916
rect 13872 2876 16672 2904
rect 13872 2864 13878 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 5902 2836 5908 2848
rect 3712 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6009 2839 6067 2845
rect 6009 2805 6021 2839
rect 6055 2836 6067 2839
rect 6362 2836 6368 2848
rect 6055 2808 6368 2836
rect 6055 2805 6067 2808
rect 6009 2799 6067 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 5442 2632 5448 2644
rect 3467 2604 5448 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 7340 2604 8309 2632
rect 7340 2592 7346 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 8297 2595 8355 2601
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 9088 2604 9137 2632
rect 9088 2592 9094 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 4856 2468 5396 2496
rect 4856 2456 4862 2468
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 5368 2437 5396 2468
rect 9232 2468 16574 2496
rect 9232 2440 9260 2468
rect 16546 2440 16574 2468
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5491 2400 5733 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 5721 2391 5779 2397
rect 4798 2320 4804 2372
rect 4856 2360 4862 2372
rect 4893 2363 4951 2369
rect 4893 2360 4905 2363
rect 4856 2332 4905 2360
rect 4856 2320 4862 2332
rect 4893 2329 4905 2332
rect 4939 2329 4951 2363
rect 4893 2323 4951 2329
rect 4982 2320 4988 2372
rect 5040 2360 5046 2372
rect 5184 2360 5212 2391
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8386 2428 8392 2440
rect 7607 2400 8392 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8812 2400 8953 2428
rect 8812 2388 8818 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 9214 2428 9220 2440
rect 9127 2400 9220 2428
rect 8941 2391 8999 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 16546 2400 16580 2440
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 8125 2363 8183 2369
rect 5040 2332 5212 2360
rect 6380 2332 6486 2360
rect 5040 2320 5046 2332
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 6380 2292 6408 2332
rect 8125 2329 8137 2363
rect 8171 2360 8183 2363
rect 8171 2332 16574 2360
rect 8171 2329 8183 2332
rect 8125 2323 8183 2329
rect 9306 2292 9312 2304
rect 4212 2264 6408 2292
rect 9219 2264 9312 2292
rect 4212 2252 4218 2264
rect 9306 2252 9312 2264
rect 9364 2292 9370 2304
rect 13814 2292 13820 2304
rect 9364 2264 13820 2292
rect 9364 2252 9370 2264
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 16546 2292 16574 2332
rect 16666 2292 16672 2304
rect 16546 2264 16672 2292
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 4948 2060 5948 2088
rect 4948 2048 4954 2060
rect 4908 2020 4936 2048
rect 5810 2020 5816 2032
rect 4264 1992 4936 2020
rect 5750 1992 5816 2020
rect 4264 1964 4292 1992
rect 5810 1980 5816 1992
rect 5868 1980 5874 2032
rect 4246 1952 4252 1964
rect 4159 1924 4252 1952
rect 4246 1912 4252 1924
rect 4304 1912 4310 1964
rect 5920 1952 5948 2060
rect 6822 2048 6828 2100
rect 6880 2088 6886 2100
rect 8665 2091 8723 2097
rect 6880 2060 7788 2088
rect 6880 2048 6886 2060
rect 7760 2020 7788 2060
rect 8665 2057 8677 2091
rect 8711 2088 8723 2091
rect 9214 2088 9220 2100
rect 8711 2060 9220 2088
rect 8711 2057 8723 2060
rect 8665 2051 8723 2057
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 8297 2023 8355 2029
rect 8297 2020 8309 2023
rect 7682 1992 8309 2020
rect 8297 1989 8309 1992
rect 8343 1989 8355 2023
rect 8297 1983 8355 1989
rect 6181 1955 6239 1961
rect 6181 1952 6193 1955
rect 5920 1924 6193 1952
rect 6181 1921 6193 1924
rect 6227 1921 6239 1955
rect 6181 1915 6239 1921
rect 8938 1912 8944 1964
rect 8996 1952 9002 1964
rect 9401 1955 9459 1961
rect 9401 1952 9413 1955
rect 8996 1924 9413 1952
rect 8996 1912 9002 1924
rect 9401 1921 9413 1924
rect 9447 1921 9459 1955
rect 9401 1915 9459 1921
rect 4525 1887 4583 1893
rect 4525 1853 4537 1887
rect 4571 1884 4583 1887
rect 5258 1884 5264 1896
rect 4571 1856 5264 1884
rect 4571 1853 4583 1856
rect 4525 1847 4583 1853
rect 5258 1844 5264 1856
rect 5316 1844 5322 1896
rect 5997 1887 6055 1893
rect 5997 1853 6009 1887
rect 6043 1884 6055 1887
rect 6454 1884 6460 1896
rect 6043 1856 6460 1884
rect 6043 1853 6055 1856
rect 5997 1847 6055 1853
rect 6454 1844 6460 1856
rect 6512 1844 6518 1896
rect 7098 1844 7104 1896
rect 7156 1884 7162 1896
rect 8757 1887 8815 1893
rect 8757 1884 8769 1887
rect 7156 1856 8769 1884
rect 7156 1844 7162 1856
rect 8757 1853 8769 1856
rect 8803 1853 8815 1887
rect 8757 1847 8815 1853
rect 6914 1708 6920 1760
rect 6972 1748 6978 1760
rect 7929 1751 7987 1757
rect 7929 1748 7941 1751
rect 6972 1720 7941 1748
rect 6972 1708 6978 1720
rect 7929 1717 7941 1720
rect 7975 1748 7987 1751
rect 8754 1748 8760 1760
rect 7975 1720 8760 1748
rect 7975 1717 7987 1720
rect 7929 1711 7987 1717
rect 8754 1708 8760 1720
rect 8812 1708 8818 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 4798 1504 4804 1556
rect 4856 1544 4862 1556
rect 5074 1544 5080 1556
rect 4856 1516 5080 1544
rect 4856 1504 4862 1516
rect 5074 1504 5080 1516
rect 5132 1504 5138 1556
rect 6086 1544 6092 1556
rect 6047 1516 6092 1544
rect 6086 1504 6092 1516
rect 6144 1504 6150 1556
rect 3605 1411 3663 1417
rect 3605 1377 3617 1411
rect 3651 1408 3663 1411
rect 3694 1408 3700 1420
rect 3651 1380 3700 1408
rect 3651 1377 3663 1380
rect 3605 1371 3663 1377
rect 3694 1368 3700 1380
rect 3752 1368 3758 1420
rect 8113 1411 8171 1417
rect 8113 1377 8125 1411
rect 8159 1408 8171 1411
rect 9306 1408 9312 1420
rect 8159 1380 9312 1408
rect 8159 1377 8171 1380
rect 8113 1371 8171 1377
rect 9306 1368 9312 1380
rect 9364 1368 9370 1420
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1309 3387 1343
rect 5353 1343 5411 1349
rect 5353 1340 5365 1343
rect 4738 1312 5365 1340
rect 3329 1303 3387 1309
rect 5353 1309 5365 1312
rect 5399 1340 5411 1343
rect 5537 1343 5595 1349
rect 5537 1340 5549 1343
rect 5399 1312 5549 1340
rect 5399 1309 5411 1312
rect 5353 1303 5411 1309
rect 5537 1309 5549 1312
rect 5583 1340 5595 1343
rect 5810 1340 5816 1352
rect 5583 1312 5816 1340
rect 5583 1309 5595 1312
rect 5537 1303 5595 1309
rect 3344 1272 3372 1303
rect 5810 1300 5816 1312
rect 5868 1340 5874 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5868 1312 5917 1340
rect 5868 1300 5874 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6454 1300 6460 1352
rect 6512 1340 6518 1352
rect 6733 1343 6791 1349
rect 6733 1340 6745 1343
rect 6512 1312 6745 1340
rect 6512 1300 6518 1312
rect 6733 1309 6745 1312
rect 6779 1309 6791 1343
rect 6733 1303 6791 1309
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1309 6883 1343
rect 6825 1303 6883 1309
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1309 7987 1343
rect 8294 1340 8300 1352
rect 8255 1312 8300 1340
rect 7929 1303 7987 1309
rect 3344 1244 3464 1272
rect 3436 1204 3464 1244
rect 5074 1232 5080 1284
rect 5132 1272 5138 1284
rect 6840 1272 6868 1303
rect 5132 1244 6868 1272
rect 7944 1272 7972 1303
rect 8294 1300 8300 1312
rect 8352 1300 8358 1352
rect 8849 1343 8907 1349
rect 8849 1309 8861 1343
rect 8895 1340 8907 1343
rect 9493 1343 9551 1349
rect 9493 1340 9505 1343
rect 8895 1312 9505 1340
rect 8895 1309 8907 1312
rect 8849 1303 8907 1309
rect 9493 1309 9505 1312
rect 9539 1309 9551 1343
rect 9493 1303 9551 1309
rect 8941 1275 8999 1281
rect 8941 1272 8953 1275
rect 7944 1244 8953 1272
rect 5132 1232 5138 1244
rect 8941 1241 8953 1244
rect 8987 1241 8999 1275
rect 8941 1235 8999 1241
rect 4246 1204 4252 1216
rect 3436 1176 4252 1204
rect 4246 1164 4252 1176
rect 4304 1164 4310 1216
rect 5994 1164 6000 1216
rect 6052 1204 6058 1216
rect 7469 1207 7527 1213
rect 7469 1204 7481 1207
rect 6052 1176 7481 1204
rect 6052 1164 6058 1176
rect 7469 1173 7481 1176
rect 7515 1173 7527 1207
rect 7469 1167 7527 1173
rect 7745 1207 7803 1213
rect 7745 1173 7757 1207
rect 7791 1204 7803 1207
rect 8202 1204 8208 1216
rect 7791 1176 8208 1204
rect 7791 1173 7803 1176
rect 7745 1167 7803 1173
rect 8202 1164 8208 1176
rect 8260 1164 8266 1216
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 4160 11500 4212 11552
rect 4896 11500 4948 11552
rect 6368 11500 6420 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 2320 11296 2372 11348
rect 1860 11228 1912 11280
rect 3608 11228 3660 11280
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2320 11092 2372 11144
rect 3332 11160 3384 11212
rect 5540 11296 5592 11348
rect 6000 11296 6052 11348
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 8208 11296 8260 11348
rect 4436 11271 4488 11280
rect 4436 11237 4445 11271
rect 4445 11237 4479 11271
rect 4479 11237 4488 11271
rect 4436 11228 4488 11237
rect 4528 11228 4580 11280
rect 4344 11160 4396 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4988 11160 5040 11212
rect 5540 11160 5592 11212
rect 7012 11160 7064 11212
rect 7104 11092 7156 11144
rect 7656 11092 7708 11144
rect 13820 11228 13872 11280
rect 9496 11092 9548 11144
rect 1400 11024 1452 11076
rect 4804 11024 4856 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 2596 10956 2648 11008
rect 3516 10956 3568 11008
rect 3608 10999 3660 11008
rect 3608 10965 3617 10999
rect 3617 10965 3651 10999
rect 3651 10965 3660 10999
rect 4988 11067 5040 11076
rect 4988 11033 4997 11067
rect 4997 11033 5031 11067
rect 5031 11033 5040 11067
rect 4988 11024 5040 11033
rect 6552 11024 6604 11076
rect 6828 11067 6880 11076
rect 6828 11033 6837 11067
rect 6837 11033 6871 11067
rect 6871 11033 6880 11067
rect 6828 11024 6880 11033
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 7196 11024 7248 11076
rect 8300 11024 8352 11076
rect 5448 10999 5500 11008
rect 3608 10956 3660 10965
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 5816 10956 5868 11008
rect 6184 10999 6236 11008
rect 6184 10965 6193 10999
rect 6193 10965 6227 10999
rect 6227 10965 6236 10999
rect 6184 10956 6236 10965
rect 6644 10956 6696 11008
rect 7656 10956 7708 11008
rect 8024 10956 8076 11008
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 1400 10795 1452 10804
rect 1400 10761 1409 10795
rect 1409 10761 1443 10795
rect 1443 10761 1452 10795
rect 1400 10752 1452 10761
rect 4252 10752 4304 10804
rect 4988 10752 5040 10804
rect 5816 10752 5868 10804
rect 7472 10752 7524 10804
rect 7656 10752 7708 10804
rect 8116 10752 8168 10804
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 2596 10684 2648 10736
rect 5264 10684 5316 10736
rect 7104 10727 7156 10736
rect 7104 10693 7113 10727
rect 7113 10693 7147 10727
rect 7147 10693 7156 10727
rect 7104 10684 7156 10693
rect 7380 10684 7432 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2044 10616 2096 10668
rect 3516 10616 3568 10668
rect 4344 10616 4396 10668
rect 5632 10616 5684 10668
rect 6184 10659 6236 10668
rect 6184 10625 6198 10659
rect 6198 10625 6232 10659
rect 6232 10625 6236 10659
rect 6920 10659 6972 10668
rect 6184 10616 6236 10625
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7288 10616 7340 10668
rect 2412 10548 2464 10600
rect 4620 10548 4672 10600
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 6552 10548 6604 10600
rect 9312 10659 9364 10668
rect 7472 10548 7524 10600
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 2228 10412 2280 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 6736 10412 6788 10464
rect 8392 10548 8444 10600
rect 13820 10480 13872 10532
rect 8024 10412 8076 10464
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 2412 10208 2464 10260
rect 4160 10208 4212 10260
rect 4712 10208 4764 10260
rect 1584 10140 1636 10192
rect 6920 10208 6972 10260
rect 8484 10208 8536 10260
rect 13820 10208 13872 10260
rect 7564 10140 7616 10192
rect 8668 10140 8720 10192
rect 1400 10072 1452 10124
rect 1768 10004 1820 10056
rect 2320 10072 2372 10124
rect 6828 10072 6880 10124
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 8392 10072 8444 10124
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 2964 9936 3016 9988
rect 4896 9936 4948 9988
rect 6920 9936 6972 9988
rect 8392 9936 8444 9988
rect 3792 9868 3844 9920
rect 6552 9868 6604 9920
rect 7288 9868 7340 9920
rect 8668 9868 8720 9920
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 6092 9664 6144 9716
rect 4436 9596 4488 9648
rect 6184 9639 6236 9648
rect 1676 9528 1728 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 4804 9528 4856 9580
rect 5448 9528 5500 9580
rect 6184 9605 6193 9639
rect 6193 9605 6227 9639
rect 6227 9605 6236 9639
rect 6184 9596 6236 9605
rect 6552 9639 6604 9648
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 7104 9664 7156 9716
rect 8116 9664 8168 9716
rect 8208 9596 8260 9648
rect 7196 9528 7248 9580
rect 1768 9460 1820 9512
rect 3148 9460 3200 9512
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4068 9460 4120 9512
rect 7564 9460 7616 9512
rect 1400 9392 1452 9444
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 5816 9324 5868 9376
rect 9036 9324 9088 9376
rect 9588 9324 9640 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 3240 9120 3292 9172
rect 3516 9120 3568 9172
rect 4160 9163 4212 9172
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 4896 9163 4948 9172
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 1584 9052 1636 9104
rect 4712 9052 4764 9104
rect 6644 9120 6696 9172
rect 6828 9120 6880 9172
rect 7196 9120 7248 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 6184 9052 6236 9104
rect 8760 9052 8812 9104
rect 3056 8984 3108 9036
rect 4252 8984 4304 9036
rect 1308 8959 1360 8968
rect 1308 8925 1317 8959
rect 1317 8925 1351 8959
rect 1351 8925 1360 8959
rect 1308 8916 1360 8925
rect 2228 8916 2280 8968
rect 3792 8959 3844 8968
rect 1492 8848 1544 8900
rect 2412 8848 2464 8900
rect 2872 8848 2924 8900
rect 3240 8848 3292 8900
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 5540 8984 5592 9036
rect 7472 8984 7524 9036
rect 7656 8984 7708 9036
rect 3976 8848 4028 8900
rect 2228 8780 2280 8832
rect 3056 8780 3108 8832
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 4988 8848 5040 8900
rect 5540 8848 5592 8900
rect 6092 8848 6144 8900
rect 5448 8780 5500 8832
rect 5632 8780 5684 8832
rect 7564 8916 7616 8968
rect 13636 8984 13688 9036
rect 8852 8916 8904 8968
rect 6552 8848 6604 8900
rect 7380 8780 7432 8832
rect 7472 8780 7524 8832
rect 8208 8848 8260 8900
rect 8944 8848 8996 8900
rect 13728 8780 13780 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 1400 8619 1452 8628
rect 1400 8585 1409 8619
rect 1409 8585 1443 8619
rect 1443 8585 1452 8619
rect 1400 8576 1452 8585
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3056 8576 3108 8628
rect 3608 8508 3660 8560
rect 4252 8508 4304 8560
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 3424 8440 3476 8492
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4804 8508 4856 8560
rect 6828 8576 6880 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 5264 8440 5316 8492
rect 5908 8440 5960 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 2872 8372 2924 8424
rect 4804 8372 4856 8424
rect 6828 8440 6880 8492
rect 7104 8440 7156 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 8760 8440 8812 8492
rect 8944 8440 8996 8492
rect 7288 8372 7340 8424
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 13544 8576 13596 8628
rect 4896 8304 4948 8356
rect 5540 8347 5592 8356
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 5816 8304 5868 8356
rect 4620 8236 4672 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6552 8236 6604 8288
rect 6736 8236 6788 8288
rect 8760 8304 8812 8356
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 4436 8032 4488 8084
rect 3056 7964 3108 8016
rect 5632 8007 5684 8016
rect 5632 7973 5641 8007
rect 5641 7973 5675 8007
rect 5675 7973 5684 8007
rect 5632 7964 5684 7973
rect 1400 7896 1452 7948
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 2872 7896 2924 7948
rect 1768 7760 1820 7812
rect 3148 7760 3200 7812
rect 6184 7896 6236 7948
rect 8576 8032 8628 8084
rect 9312 8032 9364 8084
rect 6552 7964 6604 8016
rect 7104 7964 7156 8016
rect 7748 7964 7800 8016
rect 8024 7964 8076 8016
rect 6736 7896 6788 7948
rect 4804 7828 4856 7880
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5264 7828 5316 7880
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6644 7871 6696 7880
rect 6000 7828 6052 7837
rect 6184 7760 6236 7812
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7472 7828 7524 7880
rect 7840 7828 7892 7880
rect 7564 7803 7616 7812
rect 3424 7692 3476 7744
rect 4344 7692 4396 7744
rect 6368 7692 6420 7744
rect 7104 7692 7156 7744
rect 7564 7769 7573 7803
rect 7573 7769 7607 7803
rect 7607 7769 7616 7803
rect 7564 7760 7616 7769
rect 8944 7896 8996 7948
rect 8484 7828 8536 7880
rect 7840 7692 7892 7744
rect 9220 7760 9272 7812
rect 8484 7692 8536 7744
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 1308 7531 1360 7540
rect 1308 7497 1317 7531
rect 1317 7497 1351 7531
rect 1351 7497 1360 7531
rect 1308 7488 1360 7497
rect 1492 7488 1544 7540
rect 2872 7420 2924 7472
rect 1676 7352 1728 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3884 7488 3936 7540
rect 4620 7488 4672 7540
rect 6000 7420 6052 7472
rect 7656 7420 7708 7472
rect 8852 7488 8904 7540
rect 8484 7420 8536 7472
rect 3056 7352 3108 7361
rect 1400 7148 1452 7200
rect 3424 7352 3476 7404
rect 5356 7395 5408 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 5540 7352 5592 7404
rect 7012 7352 7064 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 4528 7284 4580 7336
rect 7196 7284 7248 7336
rect 5540 7216 5592 7268
rect 7840 7216 7892 7268
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 8852 7148 8904 7200
rect 9128 7148 9180 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 1308 6944 1360 6996
rect 8760 6944 8812 6996
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 1400 6808 1452 6860
rect 1768 6808 1820 6860
rect 1676 6672 1728 6724
rect 4068 6808 4120 6860
rect 6644 6808 6696 6860
rect 7380 6808 7432 6860
rect 3148 6672 3200 6724
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 6276 6740 6328 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8300 6876 8352 6928
rect 13728 6808 13780 6860
rect 8576 6783 8628 6792
rect 8116 6672 8168 6724
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8484 6672 8536 6724
rect 6552 6604 6604 6656
rect 6736 6604 6788 6656
rect 7380 6604 7432 6656
rect 9312 6604 9364 6656
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 1676 6400 1728 6452
rect 2412 6400 2464 6452
rect 4988 6400 5040 6452
rect 7196 6400 7248 6452
rect 7840 6400 7892 6452
rect 4160 6332 4212 6384
rect 7932 6375 7984 6384
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 7932 6332 7984 6341
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 5540 6264 5592 6316
rect 5724 6264 5776 6316
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8760 6307 8812 6316
rect 8484 6264 8536 6273
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 8852 6264 8904 6316
rect 9588 6264 9640 6316
rect 6092 6196 6144 6248
rect 8116 6196 8168 6248
rect 8208 6128 8260 6180
rect 9496 6128 9548 6180
rect 4804 6060 4856 6112
rect 7012 6060 7064 6112
rect 8116 6060 8168 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1676 5856 1728 5908
rect 2412 5856 2464 5908
rect 7380 5856 7432 5908
rect 8576 5856 8628 5908
rect 1676 5652 1728 5704
rect 3240 5584 3292 5636
rect 3700 5652 3752 5704
rect 3792 5652 3844 5704
rect 4804 5584 4856 5636
rect 8484 5788 8536 5840
rect 8760 5788 8812 5840
rect 13452 5720 13504 5772
rect 6184 5627 6236 5636
rect 6184 5593 6193 5627
rect 6193 5593 6227 5627
rect 6227 5593 6236 5627
rect 6184 5584 6236 5593
rect 8116 5652 8168 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9588 5652 9640 5704
rect 13820 5584 13872 5636
rect 3700 5516 3752 5568
rect 4896 5516 4948 5568
rect 7840 5516 7892 5568
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 8852 5516 8904 5568
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 3424 5312 3476 5364
rect 4160 5244 4212 5296
rect 5448 5312 5500 5364
rect 7012 5312 7064 5364
rect 8392 5312 8444 5364
rect 8760 5312 8812 5364
rect 3148 5176 3200 5228
rect 3976 5176 4028 5228
rect 4252 5108 4304 5160
rect 4436 5176 4488 5228
rect 5724 5176 5776 5228
rect 7472 5244 7524 5296
rect 6092 5108 6144 5160
rect 7932 5176 7984 5228
rect 8668 5176 8720 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 5172 5040 5224 5092
rect 5908 5040 5960 5092
rect 9220 5040 9272 5092
rect 4344 4972 4396 5024
rect 4712 4972 4764 5024
rect 7380 4972 7432 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8024 4972 8076 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 3424 4768 3476 4820
rect 4712 4768 4764 4820
rect 7472 4768 7524 4820
rect 13820 4768 13872 4820
rect 3608 4700 3660 4752
rect 3516 4564 3568 4616
rect 4160 4632 4212 4684
rect 4896 4700 4948 4752
rect 4068 4428 4120 4480
rect 4252 4428 4304 4480
rect 4528 4496 4580 4548
rect 4896 4428 4948 4480
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5724 4700 5776 4752
rect 6000 4700 6052 4752
rect 7932 4700 7984 4752
rect 7104 4632 7156 4684
rect 5172 4564 5224 4573
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 9312 4632 9364 4684
rect 6460 4564 6512 4573
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 6000 4496 6052 4548
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 3516 4224 3568 4276
rect 4252 4224 4304 4276
rect 5448 4224 5500 4276
rect 3148 4156 3200 4208
rect 3884 4156 3936 4208
rect 2688 4088 2740 4140
rect 3792 4088 3844 4140
rect 4068 4088 4120 4140
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 6368 4088 6420 4140
rect 3608 4020 3660 4072
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 6460 4020 6512 4072
rect 3516 3952 3568 4004
rect 4068 3884 4120 3936
rect 5540 3952 5592 4004
rect 7472 4088 7524 4140
rect 7748 4088 7800 4140
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8484 4088 8536 4140
rect 8760 4020 8812 4072
rect 13728 4088 13780 4140
rect 8392 3952 8444 4004
rect 8024 3884 8076 3936
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 4344 3680 4396 3732
rect 4620 3680 4672 3732
rect 9496 3680 9548 3732
rect 4252 3612 4304 3664
rect 4804 3655 4856 3664
rect 4804 3621 4813 3655
rect 4813 3621 4847 3655
rect 4847 3621 4856 3655
rect 4804 3612 4856 3621
rect 4988 3612 5040 3664
rect 6092 3612 6144 3664
rect 4160 3476 4212 3528
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4528 3519 4580 3528
rect 4252 3476 4304 3485
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4896 3476 4948 3528
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 5632 3476 5684 3528
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 9312 3476 9364 3528
rect 9404 3476 9456 3528
rect 4804 3408 4856 3460
rect 6184 3408 6236 3460
rect 8024 3408 8076 3460
rect 3608 3340 3660 3392
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4896 3340 4948 3392
rect 5908 3340 5960 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 4068 3136 4120 3188
rect 4436 3136 4488 3188
rect 6000 3136 6052 3188
rect 6276 3136 6328 3188
rect 5816 3068 5868 3120
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 8300 3136 8352 3188
rect 9312 3136 9364 3188
rect 6828 3068 6880 3120
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4896 3000 4948 3052
rect 4988 2864 5040 2916
rect 7012 2932 7064 2984
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 13820 2864 13872 2916
rect 16672 2864 16724 2916
rect 5908 2796 5960 2848
rect 6368 2796 6420 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 5448 2592 5500 2644
rect 7288 2592 7340 2644
rect 9036 2592 9088 2644
rect 4804 2456 4856 2508
rect 3792 2388 3844 2440
rect 6092 2431 6144 2440
rect 4804 2320 4856 2372
rect 4988 2320 5040 2372
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 8392 2388 8444 2440
rect 8760 2388 8812 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 16580 2388 16632 2440
rect 4160 2252 4212 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 13820 2252 13872 2304
rect 16672 2252 16724 2304
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 4896 2048 4948 2100
rect 5816 1980 5868 2032
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 6828 2048 6880 2100
rect 9220 2048 9272 2100
rect 8944 1912 8996 1964
rect 5264 1844 5316 1896
rect 6460 1887 6512 1896
rect 6460 1853 6469 1887
rect 6469 1853 6503 1887
rect 6503 1853 6512 1887
rect 6460 1844 6512 1853
rect 7104 1844 7156 1896
rect 6920 1708 6972 1760
rect 8760 1708 8812 1760
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 4804 1504 4856 1556
rect 5080 1547 5132 1556
rect 5080 1513 5089 1547
rect 5089 1513 5123 1547
rect 5123 1513 5132 1547
rect 5080 1504 5132 1513
rect 6092 1547 6144 1556
rect 6092 1513 6101 1547
rect 6101 1513 6135 1547
rect 6135 1513 6144 1547
rect 6092 1504 6144 1513
rect 3700 1368 3752 1420
rect 9312 1368 9364 1420
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6460 1300 6512 1352
rect 8300 1343 8352 1352
rect 5080 1232 5132 1284
rect 8300 1309 8309 1343
rect 8309 1309 8343 1343
rect 8343 1309 8352 1343
rect 8300 1300 8352 1309
rect 4252 1164 4304 1216
rect 6000 1164 6052 1216
rect 8208 1164 8260 1216
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
<< metal2 >>
rect 938 12322 994 13000
rect 1398 12322 1454 13000
rect 938 12294 1348 12322
rect 938 12200 994 12294
rect 1320 10962 1348 12294
rect 1398 12294 1532 12322
rect 1398 12200 1454 12294
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10962 1440 11018
rect 1320 10934 1440 10962
rect 1412 10810 1440 10934
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1412 10130 1440 10746
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1400 9444 1452 9450
rect 1400 9386 1452 9392
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1320 7546 1348 8910
rect 1412 8634 1440 9386
rect 1504 8906 1532 12294
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12322 2834 13000
rect 2700 12294 2834 12322
rect 1872 11286 1900 12200
rect 2332 11354 2360 12200
rect 2700 11540 2728 12294
rect 2778 12200 2834 12294
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12322 5134 13000
rect 5000 12294 5134 12322
rect 2700 11512 3096 11540
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1860 11144 1912 11150
rect 1858 11112 1860 11121
rect 2136 11144 2188 11150
rect 1912 11112 1914 11121
rect 2136 11086 2188 11092
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 1858 11047 1914 11056
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10674 2084 10950
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1596 10198 1624 10610
rect 2148 10554 2176 11086
rect 2148 10526 2268 10554
rect 2240 10470 2268 10526
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1596 8634 1624 9046
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1320 7002 1348 7482
rect 1412 7206 1440 7890
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7546 1532 7822
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1688 7410 1716 9522
rect 1780 9518 1808 9998
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1780 7818 1808 9454
rect 2240 8974 2268 10406
rect 2332 10130 2360 11086
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10742 2636 10950
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10266 2452 10542
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2872 8900 2924 8906
rect 2976 8888 3004 9930
rect 3068 9042 3096 11512
rect 3252 11336 3280 12200
rect 3252 11308 3464 11336
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2924 8860 3004 8888
rect 2872 8842 2924 8848
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8498 2268 8774
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1412 6866 1440 7142
rect 1688 6882 1716 7346
rect 1688 6866 1808 6882
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1688 6860 1820 6866
rect 1688 6854 1768 6860
rect 1688 6730 1716 6854
rect 1768 6802 1820 6808
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1688 6458 1716 6666
rect 2424 6458 2452 8842
rect 2884 8430 2912 8842
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8634 3096 8774
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3160 8514 3188 9454
rect 3252 9178 3280 9522
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3240 8900 3292 8906
rect 3344 8888 3372 11154
rect 3436 9674 3464 11308
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3620 11014 3648 11222
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3528 10674 3556 10950
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3620 10062 3648 10950
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3436 9646 3648 9674
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3292 8860 3372 8888
rect 3240 8842 3292 8848
rect 3068 8486 3188 8514
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 3068 8022 3096 8486
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2884 7478 2912 7890
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 3068 7410 3096 7958
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 3160 6730 3188 7754
rect 3344 7290 3372 8860
rect 3436 8498 3464 9318
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 8922 3648 9646
rect 3528 8894 3648 8922
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7410 3464 7686
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3344 7262 3464 7290
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 1688 5914 1716 6394
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5930 2360 6258
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2332 5914 2452 5930
rect 1676 5908 1728 5914
rect 2332 5908 2464 5914
rect 2332 5902 2412 5908
rect 1676 5850 1728 5856
rect 2412 5850 2464 5856
rect 1688 5710 1716 5850
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 3160 5234 3188 6666
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 5642 3280 6598
rect 3344 6322 3372 7142
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3436 5370 3464 7262
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3160 4214 3188 5170
rect 3436 4826 3464 5306
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3528 4622 3556 8894
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8566 3648 8774
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3712 5794 3740 12200
rect 4172 11558 4200 12200
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10810 4292 11086
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4356 10674 4384 11154
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 8974 3832 9862
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3896 7342 3924 7482
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3620 5766 3740 5794
rect 3620 4758 3648 5766
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3712 5574 3740 5646
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3528 4282 3556 4558
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2700 3445 2728 4082
rect 3620 4078 3648 4694
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 2686 3436 2742 3445
rect 2686 3371 2742 3380
rect 3528 3194 3556 3946
rect 3620 3738 3648 4014
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3620 3058 3648 3334
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3712 1426 3740 5510
rect 3804 4146 3832 5646
rect 3988 5234 4016 8842
rect 4080 6866 4108 9454
rect 4172 9178 4200 10202
rect 4448 9654 4476 11222
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4540 9178 4568 11222
rect 4632 10606 4660 12200
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 10266 4752 10406
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4816 9586 4844 11018
rect 4908 10248 4936 11494
rect 5000 11218 5028 12294
rect 5078 12200 5134 12294
rect 5538 12200 5594 13000
rect 5998 12322 6054 13000
rect 5736 12294 6054 12322
rect 5552 11354 5580 12200
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5540 11212 5592 11218
rect 5592 11172 5672 11200
rect 5540 11154 5592 11160
rect 5000 11082 5028 11154
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5000 10810 5028 11018
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5066 10908 5374 10928
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10832 5374 10852
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5276 10606 5304 10678
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 4908 10220 5028 10248
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8566 4292 8978
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 8090 4476 8434
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4434 7984 4490 7993
rect 4434 7919 4490 7928
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4172 5302 4200 6326
rect 4160 5296 4212 5302
rect 4356 5250 4384 7686
rect 4160 5238 4212 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4264 5222 4384 5250
rect 4448 5234 4476 7919
rect 4540 7342 4568 9114
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7546 4660 8230
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 5228 4488 5234
rect 4264 5166 4292 5222
rect 4436 5170 4488 5176
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4690 4200 5034
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3896 2774 3924 4150
rect 4080 4146 4108 4422
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3194 4108 3878
rect 4172 3534 4200 4626
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4282 4292 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4356 4026 4384 4966
rect 4264 3998 4384 4026
rect 4264 3670 4292 3998
rect 4344 3732 4396 3738
rect 4448 3720 4476 5170
rect 4724 5114 4752 9046
rect 4816 8566 4844 9522
rect 4908 9178 4936 9930
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 8906 5028 10220
rect 5066 9820 5374 9840
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9744 5374 9764
rect 5460 9586 5488 10950
rect 5644 10674 5672 11172
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5552 8906 5580 8978
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4816 7886 4844 8366
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 6118 4844 7822
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4632 5086 4752 5114
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4396 3692 4476 3720
rect 4344 3674 4396 3680
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4540 3534 4568 4490
rect 4632 4185 4660 5086
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4826 4752 4966
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4618 4176 4674 4185
rect 4618 4111 4674 4120
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4632 3738 4660 4014
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4816 3670 4844 5578
rect 4908 5574 4936 8298
rect 5000 7993 5028 8842
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5066 8732 5374 8752
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8656 5374 8676
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4986 7984 5042 7993
rect 4986 7919 5042 7928
rect 5276 7886 5304 8434
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5000 6458 5028 7822
rect 5066 7644 5374 7664
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7568 5374 7588
rect 5354 7440 5410 7449
rect 5354 7375 5356 7384
rect 5408 7375 5410 7384
rect 5356 7346 5408 7352
rect 5066 6556 5374 6576
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6480 5374 6500
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 5066 5468 5374 5488
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5392 5374 5412
rect 5460 5370 5488 8774
rect 5552 8673 5580 8842
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5538 8664 5594 8673
rect 5538 8599 5594 8608
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 7410 5580 8298
rect 5644 8022 5672 8774
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6322 5580 7210
rect 5736 6322 5764 12294
rect 5998 12200 6054 12294
rect 6458 12200 6514 13000
rect 9494 12336 9550 12345
rect 9494 12271 9550 12280
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11354 6408 11494
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5828 10810 5856 10950
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 8362 5856 9318
rect 5906 8800 5962 8809
rect 5906 8735 5962 8744
rect 5920 8498 5948 8735
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7993 5948 8230
rect 5906 7984 5962 7993
rect 5906 7919 5962 7928
rect 6012 7886 6040 11290
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6196 10674 6224 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 9722 6132 9998
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6196 9654 6224 10610
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6184 9104 6236 9110
rect 6472 9058 6500 12200
rect 7566 11452 7874 11472
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11376 7874 11396
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6918 11112 6974 11121
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6828 11076 6880 11082
rect 6918 11047 6920 11056
rect 6828 11018 6880 11024
rect 6972 11047 6974 11056
rect 6920 11018 6972 11024
rect 6564 10606 6592 11018
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9654 6592 9862
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6656 9178 6684 10950
rect 6840 10713 6868 11018
rect 6826 10704 6882 10713
rect 6826 10639 6882 10648
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6748 9081 6776 10406
rect 6932 10266 6960 10610
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9178 6868 10066
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6184 9046 6236 9052
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4908 4486 4936 4694
rect 5184 4622 5212 5034
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4908 3534 4936 4422
rect 5066 4380 5374 4400
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4304 5374 4324
rect 5460 4282 5488 5306
rect 5736 5234 5764 6258
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 4758 5764 5170
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5920 4622 5948 5034
rect 6012 4758 6040 7414
rect 6104 6254 6132 8842
rect 6196 8537 6224 9046
rect 6380 9030 6500 9058
rect 6734 9072 6790 9081
rect 6182 8528 6238 8537
rect 6182 8463 6184 8472
rect 6236 8463 6238 8472
rect 6184 8434 6236 8440
rect 6196 7970 6224 8434
rect 6196 7954 6316 7970
rect 6184 7948 6316 7954
rect 6236 7942 6316 7948
rect 6184 7890 6236 7896
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6104 5166 6132 6190
rect 6196 5642 6224 7754
rect 6288 6798 6316 7942
rect 6380 7834 6408 9030
rect 6734 9007 6790 9016
rect 6932 8956 6960 9930
rect 6840 8928 6960 8956
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6564 8378 6592 8842
rect 6734 8664 6790 8673
rect 6840 8634 6868 8928
rect 7024 8888 7052 11154
rect 7104 11144 7156 11150
rect 7656 11144 7708 11150
rect 7104 11086 7156 11092
rect 7484 11104 7656 11132
rect 7116 10742 7144 11086
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7116 9722 7144 10678
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9586 7236 11018
rect 7484 10810 7512 11104
rect 7656 11086 7708 11092
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7668 10810 7696 10950
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7930 10704 7986 10713
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 9926 7328 10610
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6932 8860 7052 8888
rect 6734 8599 6790 8608
rect 6828 8628 6880 8634
rect 6748 8514 6776 8599
rect 6828 8570 6880 8576
rect 6932 8514 6960 8860
rect 6656 8498 6868 8514
rect 6644 8492 6880 8498
rect 6696 8486 6828 8492
rect 6644 8434 6696 8440
rect 6932 8486 7052 8514
rect 6828 8434 6880 8440
rect 6564 8350 6960 8378
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6380 7806 6500 7834
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4264 3346 4292 3470
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3804 2746 3924 2774
rect 3804 2446 3832 2746
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4172 2310 4200 3334
rect 4264 3318 4476 3346
rect 4448 3194 4476 3318
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4816 2514 4844 3402
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5000 2922 5028 3606
rect 5552 3534 5580 3946
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3422 5672 3470
rect 5460 3394 5672 3422
rect 5920 3398 5948 4558
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 5066 3292 5374 3312
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 5066 3216 5374 3236
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5000 2378 5028 2858
rect 5460 2650 5488 3394
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6012 3194 6040 4490
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6104 3670 6132 4082
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6196 3466 6224 5578
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6288 3194 6316 6734
rect 6380 4622 6408 7686
rect 6472 7313 6500 7806
rect 6458 7304 6514 7313
rect 6458 7239 6514 7248
rect 6564 6746 6592 7958
rect 6748 7954 6776 8230
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 6866 6684 7822
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6564 6718 6684 6746
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3369 6408 4082
rect 6472 4078 6500 4558
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6366 3360 6422 3369
rect 6366 3295 6422 3304
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6564 3126 6592 6598
rect 6656 3534 6684 6718
rect 6748 6662 6776 7890
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 3700 1420 3752 1426
rect 3700 1362 3752 1368
rect 4264 1222 4292 1906
rect 4816 1562 4844 2314
rect 5000 2122 5028 2314
rect 5066 2204 5374 2224
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2128 5374 2148
rect 4908 2106 5028 2122
rect 4896 2100 5028 2106
rect 4948 2094 5028 2100
rect 4896 2042 4948 2048
rect 5264 1896 5316 1902
rect 5460 1884 5488 2586
rect 5828 2038 5856 3062
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 5316 1856 5488 1884
rect 5264 1838 5316 1844
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 5080 1556 5132 1562
rect 5080 1498 5132 1504
rect 5092 1290 5120 1498
rect 5828 1358 5856 1974
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 5920 1306 5948 2790
rect 6092 2440 6144 2446
rect 6380 2417 6408 2790
rect 6092 2382 6144 2388
rect 6366 2408 6422 2417
rect 6104 1562 6132 2382
rect 6366 2343 6422 2352
rect 6840 2106 6868 3062
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6472 1358 6500 1838
rect 6932 1766 6960 8350
rect 7024 7410 7052 8486
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 8022 7144 8434
rect 7208 8106 7236 9114
rect 7286 9072 7342 9081
rect 7286 9007 7342 9016
rect 7300 8430 7328 9007
rect 7392 8838 7420 10678
rect 7930 10639 7986 10648
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 9042 7512 10542
rect 7566 10364 7874 10384
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10288 7874 10308
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7576 9518 7604 10134
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7566 9276 7874 9296
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9200 7874 9220
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 8832 7432 8838
rect 7472 8832 7524 8838
rect 7380 8774 7432 8780
rect 7470 8800 7472 8809
rect 7524 8800 7526 8809
rect 7392 8498 7420 8774
rect 7470 8735 7526 8744
rect 7576 8537 7604 8910
rect 7562 8528 7618 8537
rect 7380 8492 7432 8498
rect 7562 8463 7618 8472
rect 7380 8434 7432 8440
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7208 8078 7328 8106
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7194 7712 7250 7721
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 7024 6118 7052 7239
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5370 7052 6054
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7024 2990 7052 5306
rect 7116 4690 7144 7686
rect 7194 7647 7250 7656
rect 7208 7342 7236 7647
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7194 7168 7250 7177
rect 7194 7103 7250 7112
rect 7208 6458 7236 7103
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7116 1902 7144 3470
rect 7300 2650 7328 8078
rect 7392 6866 7420 8434
rect 7668 8430 7696 8978
rect 7656 8424 7708 8430
rect 7654 8392 7656 8401
rect 7708 8392 7710 8401
rect 7654 8327 7710 8336
rect 7566 8188 7874 8208
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8112 7874 8132
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 5914 7420 6598
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7392 5030 7420 5850
rect 7484 5302 7512 7822
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 7449 7604 7754
rect 7656 7472 7708 7478
rect 7562 7440 7618 7449
rect 7760 7449 7788 7958
rect 7840 7880 7892 7886
rect 7838 7848 7840 7857
rect 7892 7848 7894 7857
rect 7838 7783 7894 7792
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7656 7414 7708 7420
rect 7746 7440 7802 7449
rect 7562 7375 7618 7384
rect 7668 7313 7696 7414
rect 7746 7375 7802 7384
rect 7654 7304 7710 7313
rect 7852 7274 7880 7686
rect 7654 7239 7710 7248
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7566 7100 7874 7120
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7024 7874 7044
rect 7838 6896 7894 6905
rect 7838 6831 7894 6840
rect 7852 6798 7880 6831
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7852 6100 7880 6394
rect 7944 6390 7972 10639
rect 8036 10470 8064 10950
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 8022 8064 10406
rect 8128 9722 8156 10746
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9654 8248 11290
rect 9508 11150 9536 12271
rect 13818 11928 13874 11937
rect 13818 11863 13874 11872
rect 13450 11520 13506 11529
rect 13450 11455 13506 11464
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8114 7848 8170 7857
rect 8114 7783 8170 7792
rect 8022 7304 8078 7313
rect 8022 7239 8078 7248
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7852 6072 7972 6100
rect 7566 6012 7874 6032
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5936 7874 5956
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7852 5137 7880 5510
rect 7944 5234 7972 6072
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7838 5128 7894 5137
rect 7838 5063 7894 5072
rect 8036 5030 8064 7239
rect 8128 7041 8156 7783
rect 8114 7032 8170 7041
rect 8114 6967 8170 6976
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8128 6254 8156 6666
rect 8220 6304 8248 8842
rect 8312 6934 8340 11018
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8404 10130 8432 10542
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8496 10266 8524 10406
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8680 10198 8708 10406
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 7721 8432 9930
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8482 8392 8538 8401
rect 8482 8327 8538 8336
rect 8496 7886 8524 8327
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8484 7744 8536 7750
rect 8390 7712 8446 7721
rect 8484 7686 8536 7692
rect 8390 7647 8446 7656
rect 8496 7478 8524 7686
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8220 6276 8340 6304
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5710 8156 6054
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7566 4924 7874 4944
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4848 7874 4868
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4146 7512 4762
rect 7944 4758 7972 4966
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7746 4176 7802 4185
rect 7472 4140 7524 4146
rect 8128 4146 8156 5510
rect 8220 5409 8248 6122
rect 8206 5400 8262 5409
rect 8206 5335 8262 5344
rect 8312 5250 8340 6276
rect 8404 5370 8432 7346
rect 8496 6730 8524 7414
rect 8588 6882 8616 8026
rect 8680 7449 8708 9862
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8772 8498 8800 9046
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8864 8378 8892 8910
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8498 8984 8842
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8772 8362 8892 8378
rect 8760 8356 8892 8362
rect 8812 8350 8892 8356
rect 8760 8298 8812 8304
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8772 7002 8800 8298
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8850 7576 8906 7585
rect 8850 7511 8852 7520
rect 8904 7511 8906 7520
rect 8852 7482 8904 7488
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8588 6854 8708 6882
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8482 6624 8538 6633
rect 8482 6559 8538 6568
rect 8496 6322 8524 6559
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8588 5914 8616 6734
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8220 5222 8340 5250
rect 7746 4111 7748 4120
rect 7472 4082 7524 4088
rect 7800 4111 7802 4120
rect 8116 4140 8168 4146
rect 7748 4082 7800 4088
rect 8116 4082 8168 4088
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7566 3836 7874 3856
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3760 7874 3780
rect 8036 3466 8064 3878
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7566 2748 7874 2768
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2672 7874 2692
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 7566 1660 7874 1680
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1584 7874 1604
rect 6460 1352 6512 1358
rect 5080 1284 5132 1290
rect 5920 1278 6040 1306
rect 6460 1294 6512 1300
rect 5080 1226 5132 1232
rect 6012 1222 6040 1278
rect 8220 1222 8248 5222
rect 8496 4146 8524 5782
rect 8680 5234 8708 6854
rect 8864 6322 8892 7142
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8772 5846 8800 6258
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 5370 8800 5782
rect 8852 5568 8904 5574
rect 8956 5556 8984 7890
rect 9048 7002 9076 9318
rect 9232 7818 9260 10950
rect 9508 10810 9536 11086
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 8090 9352 10610
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9178 9444 9998
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 8634 9536 10231
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9324 7410 9352 7919
rect 9600 7857 9628 9318
rect 9586 7848 9642 7857
rect 9586 7783 9642 7792
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9048 6225 9076 6938
rect 9034 6216 9090 6225
rect 9034 6151 9090 6160
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8904 5528 8984 5556
rect 8852 5510 8904 5516
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8864 5216 8892 5510
rect 8944 5228 8996 5234
rect 8864 5188 8944 5216
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8312 3194 8340 4082
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8312 1358 8340 3130
rect 8404 2446 8432 3946
rect 8772 3126 8800 4014
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8772 1766 8800 2382
rect 8760 1760 8812 1766
rect 8864 1737 8892 5188
rect 8944 5170 8996 5176
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 1970 8984 3878
rect 9048 2650 9076 5646
rect 9140 3777 9168 7142
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5114 9352 6598
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9508 5234 9536 6122
rect 9600 5710 9628 6258
rect 13464 5778 13492 11455
rect 13832 11286 13860 11863
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13832 10538 13860 11047
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13542 9888 13598 9897
rect 13542 9823 13598 9832
rect 13556 8634 13584 9823
rect 13832 9489 13860 10202
rect 13818 9480 13874 9489
rect 13818 9415 13874 9424
rect 13818 9072 13874 9081
rect 13636 9036 13688 9042
rect 13818 9007 13874 9016
rect 13636 8978 13688 8984
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13648 8265 13676 8978
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 8673 13768 8774
rect 13726 8664 13782 8673
rect 13726 8599 13782 8608
rect 13634 8256 13690 8265
rect 13634 8191 13690 8200
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13740 6633 13768 6802
rect 13726 6624 13782 6633
rect 13726 6559 13782 6568
rect 13726 5808 13782 5817
rect 13452 5772 13504 5778
rect 13726 5743 13782 5752
rect 13452 5714 13504 5720
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9220 5092 9272 5098
rect 9324 5086 9444 5114
rect 9220 5034 9272 5040
rect 9232 4622 9260 5034
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4690 9352 4966
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9126 3768 9182 3777
rect 9126 3703 9182 3712
rect 9324 3534 9352 4422
rect 9416 3534 9444 5086
rect 9494 4584 9550 4593
rect 9600 4570 9628 5646
rect 9550 4542 9628 4570
rect 9494 4519 9550 4528
rect 9508 3738 9536 4519
rect 13740 4146 13768 5743
rect 13832 5642 13860 9007
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13832 4185 13860 4762
rect 13818 4176 13874 4185
rect 13728 4140 13780 4146
rect 13818 4111 13874 4120
rect 13728 4082 13780 4088
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3194 9352 3334
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 13818 2952 13874 2961
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9232 2106 9260 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 8760 1702 8812 1708
rect 8850 1728 8906 1737
rect 8850 1663 8906 1672
rect 9324 1426 9352 2246
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 4252 1216 4304 1222
rect 4252 1158 4304 1164
rect 6000 1216 6052 1222
rect 6000 1158 6052 1164
rect 8208 1216 8260 1222
rect 8208 1158 8260 1164
rect 5066 1116 5374 1136
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1040 5374 1060
rect 9416 921 9444 2926
rect 13818 2887 13820 2896
rect 13872 2887 13874 2896
rect 16672 2916 16724 2922
rect 13820 2858 13872 2864
rect 16672 2858 16724 2864
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 9402 912 9458 921
rect 9402 847 9458 856
rect 9508 513 9536 2382
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13832 1329 13860 2246
rect 16592 2145 16620 2382
rect 16684 2310 16712 2858
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 13818 1320 13874 1329
rect 13818 1255 13874 1264
rect 9494 504 9550 513
rect 9494 439 9550 448
<< via2 >>
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 1858 11092 1860 11112
rect 1860 11092 1912 11112
rect 1912 11092 1914 11112
rect 1858 11056 1914 11092
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2686 3380 2742 3436
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 4434 7928 4490 7984
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 4618 4120 4674 4176
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 4986 7928 5042 7984
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5354 7404 5410 7440
rect 5354 7384 5356 7404
rect 5356 7384 5408 7404
rect 5408 7384 5410 7404
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5538 8608 5594 8664
rect 9494 12280 9550 12336
rect 5906 8744 5962 8800
rect 5906 7928 5962 7984
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 6918 11076 6974 11112
rect 6918 11056 6920 11076
rect 6920 11056 6972 11076
rect 6972 11056 6974 11076
rect 6826 10648 6882 10704
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 6182 8492 6238 8528
rect 6182 8472 6184 8492
rect 6184 8472 6236 8492
rect 6236 8472 6238 8492
rect 6734 9016 6790 9072
rect 6734 8608 6790 8664
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 6458 7248 6514 7304
rect 6366 3304 6422 3360
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 6366 2352 6422 2408
rect 7286 9016 7342 9072
rect 7930 10648 7986 10704
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7470 8780 7472 8800
rect 7472 8780 7524 8800
rect 7524 8780 7526 8800
rect 7470 8744 7526 8780
rect 7562 8472 7618 8528
rect 7010 7248 7066 7304
rect 7194 7656 7250 7712
rect 7194 7112 7250 7168
rect 7654 8372 7656 8392
rect 7656 8372 7708 8392
rect 7708 8372 7710 8392
rect 7654 8336 7710 8372
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 7562 7384 7618 7440
rect 7838 7828 7840 7848
rect 7840 7828 7892 7848
rect 7892 7828 7894 7848
rect 7838 7792 7894 7828
rect 7746 7384 7802 7440
rect 7654 7248 7710 7304
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7838 6840 7894 6896
rect 13818 11872 13874 11928
rect 13450 11464 13506 11520
rect 8114 7792 8170 7848
rect 8022 7248 8078 7304
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7838 5072 7894 5128
rect 8114 6976 8170 7032
rect 8482 8336 8538 8392
rect 8390 7656 8446 7712
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7746 4140 7802 4176
rect 8206 5344 8262 5400
rect 8666 7384 8722 7440
rect 8850 7540 8906 7576
rect 8850 7520 8852 7540
rect 8852 7520 8904 7540
rect 8904 7520 8906 7540
rect 8482 6568 8538 6624
rect 7746 4120 7748 4140
rect 7748 4120 7800 4140
rect 7800 4120 7802 4140
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 9494 10240 9550 10296
rect 9310 7928 9366 7984
rect 9586 7792 9642 7848
rect 9034 6160 9090 6216
rect 13818 11056 13874 11112
rect 13542 9832 13598 9888
rect 13818 9424 13874 9480
rect 13818 9016 13874 9072
rect 13726 8608 13782 8664
rect 13634 8200 13690 8256
rect 13726 6568 13782 6624
rect 13726 5752 13782 5808
rect 9126 3712 9182 3768
rect 9494 4528 9550 4584
rect 13818 4120 13874 4176
rect 8850 1672 8906 1728
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 13818 2916 13874 2952
rect 13818 2896 13820 2916
rect 13820 2896 13872 2916
rect 13872 2896 13874 2916
rect 9402 856 9458 912
rect 16578 2080 16634 2136
rect 13818 1264 13874 1320
rect 9494 448 9550 504
<< metal3 >>
rect 9489 12338 9555 12341
rect 14000 12338 34000 12368
rect 9489 12336 34000 12338
rect 9489 12280 9494 12336
rect 9550 12280 34000 12336
rect 9489 12278 34000 12280
rect 9489 12275 9555 12278
rect 14000 12248 34000 12278
rect 13813 11930 13879 11933
rect 14000 11930 34000 11960
rect 13813 11928 34000 11930
rect 13813 11872 13818 11928
rect 13874 11872 34000 11928
rect 13813 11870 34000 11872
rect 13813 11867 13879 11870
rect 14000 11840 34000 11870
rect 13445 11522 13511 11525
rect 14000 11522 34000 11552
rect 13445 11520 34000 11522
rect 13445 11464 13450 11520
rect 13506 11464 34000 11520
rect 13445 11462 34000 11464
rect 13445 11459 13511 11462
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 7560 11456 7880 11457
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 14000 11432 34000 11462
rect 7560 11391 7880 11392
rect 1853 11114 1919 11117
rect 6913 11114 6979 11117
rect 1853 11112 6979 11114
rect 1853 11056 1858 11112
rect 1914 11056 6918 11112
rect 6974 11056 6979 11112
rect 1853 11054 6979 11056
rect 1853 11051 1919 11054
rect 6913 11051 6979 11054
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10847 5380 10848
rect 6821 10706 6887 10709
rect 7925 10706 7991 10709
rect 14000 10706 34000 10736
rect 6821 10704 34000 10706
rect 6821 10648 6826 10704
rect 6882 10648 7930 10704
rect 7986 10648 34000 10704
rect 6821 10646 34000 10648
rect 6821 10643 6887 10646
rect 7925 10643 7991 10646
rect 14000 10616 34000 10646
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 7560 10368 7880 10369
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 10303 7880 10304
rect 9489 10298 9555 10301
rect 14000 10298 34000 10328
rect 9489 10296 34000 10298
rect 9489 10240 9494 10296
rect 9550 10240 34000 10296
rect 9489 10238 34000 10240
rect 9489 10235 9555 10238
rect 14000 10208 34000 10238
rect 13537 9890 13603 9893
rect 14000 9890 34000 9920
rect 13537 9888 34000 9890
rect 13537 9832 13542 9888
rect 13598 9832 34000 9888
rect 13537 9830 34000 9832
rect 13537 9827 13603 9830
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9830
rect 5060 9759 5380 9760
rect 13813 9482 13879 9485
rect 14000 9482 34000 9512
rect 13813 9480 34000 9482
rect 13813 9424 13818 9480
rect 13874 9424 34000 9480
rect 13813 9422 34000 9424
rect 13813 9419 13879 9422
rect 14000 9392 34000 9422
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 7560 9280 7880 9281
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9215 7880 9216
rect 6729 9074 6795 9077
rect 7281 9074 7347 9077
rect 6729 9072 7347 9074
rect 6729 9016 6734 9072
rect 6790 9016 7286 9072
rect 7342 9016 7347 9072
rect 6729 9014 7347 9016
rect 6729 9011 6795 9014
rect 7281 9011 7347 9014
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 14000 8984 34000 9014
rect 5901 8802 5967 8805
rect 7465 8802 7531 8805
rect 5901 8800 7531 8802
rect 5901 8744 5906 8800
rect 5962 8744 7470 8800
rect 7526 8744 7531 8800
rect 5901 8742 7531 8744
rect 5901 8739 5967 8742
rect 7465 8739 7531 8742
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 8671 5380 8672
rect 5533 8666 5599 8669
rect 6729 8666 6795 8669
rect 5533 8664 6795 8666
rect 5533 8608 5538 8664
rect 5594 8608 6734 8664
rect 6790 8608 6795 8664
rect 5533 8606 6795 8608
rect 5533 8603 5599 8606
rect 6729 8603 6795 8606
rect 13721 8666 13787 8669
rect 14000 8666 34000 8696
rect 13721 8664 34000 8666
rect 13721 8608 13726 8664
rect 13782 8608 34000 8664
rect 13721 8606 34000 8608
rect 13721 8603 13787 8606
rect 14000 8576 34000 8606
rect 6177 8530 6243 8533
rect 7557 8530 7623 8533
rect 6177 8528 7623 8530
rect 6177 8472 6182 8528
rect 6238 8472 7562 8528
rect 7618 8472 7623 8528
rect 6177 8470 7623 8472
rect 6177 8467 6243 8470
rect 7557 8467 7623 8470
rect 7649 8394 7715 8397
rect 8477 8394 8543 8397
rect 7649 8392 8543 8394
rect 7649 8336 7654 8392
rect 7710 8336 8482 8392
rect 8538 8336 8543 8392
rect 7649 8334 8543 8336
rect 7649 8331 7715 8334
rect 8477 8331 8543 8334
rect 13629 8258 13695 8261
rect 14000 8258 34000 8288
rect 13629 8256 34000 8258
rect 13629 8200 13634 8256
rect 13690 8200 34000 8256
rect 13629 8198 34000 8200
rect 13629 8195 13695 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 7560 8192 7880 8193
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 14000 8168 34000 8198
rect 7560 8127 7880 8128
rect 4429 7986 4495 7989
rect 4981 7986 5047 7989
rect 4429 7984 5047 7986
rect 4429 7928 4434 7984
rect 4490 7928 4986 7984
rect 5042 7928 5047 7984
rect 4429 7926 5047 7928
rect 4429 7923 4495 7926
rect 4981 7923 5047 7926
rect 5901 7986 5967 7989
rect 9305 7986 9371 7989
rect 5901 7984 9371 7986
rect 5901 7928 5906 7984
rect 5962 7928 9310 7984
rect 9366 7928 9371 7984
rect 5901 7926 9371 7928
rect 5901 7923 5967 7926
rect 9305 7923 9371 7926
rect 7833 7850 7899 7853
rect 8109 7850 8175 7853
rect 7833 7848 8175 7850
rect 7833 7792 7838 7848
rect 7894 7792 8114 7848
rect 8170 7792 8175 7848
rect 7833 7790 8175 7792
rect 7833 7787 7899 7790
rect 8109 7787 8175 7790
rect 9581 7850 9647 7853
rect 14000 7850 34000 7880
rect 9581 7848 34000 7850
rect 9581 7792 9586 7848
rect 9642 7792 34000 7848
rect 9581 7790 34000 7792
rect 9581 7787 9647 7790
rect 14000 7760 34000 7790
rect 7189 7714 7255 7717
rect 8385 7714 8451 7717
rect 7189 7712 8451 7714
rect 7189 7656 7194 7712
rect 7250 7656 8390 7712
rect 8446 7656 8451 7712
rect 7189 7654 8451 7656
rect 7189 7651 7255 7654
rect 8385 7651 8451 7654
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7583 5380 7584
rect 8845 7578 8911 7581
rect 5582 7576 8911 7578
rect 5582 7520 8850 7576
rect 8906 7520 8911 7576
rect 5582 7518 8911 7520
rect 5349 7442 5415 7445
rect 5582 7442 5642 7518
rect 8845 7515 8911 7518
rect 7557 7442 7623 7445
rect 5349 7440 5642 7442
rect 5349 7384 5354 7440
rect 5410 7384 5642 7440
rect 5349 7382 5642 7384
rect 7238 7440 7623 7442
rect 7238 7384 7562 7440
rect 7618 7384 7623 7440
rect 7238 7382 7623 7384
rect 5349 7379 5415 7382
rect 6453 7306 6519 7309
rect 7005 7306 7071 7309
rect 6453 7304 7071 7306
rect 6453 7248 6458 7304
rect 6514 7248 7010 7304
rect 7066 7248 7071 7304
rect 6453 7246 7071 7248
rect 6453 7243 6519 7246
rect 7005 7243 7071 7246
rect 7238 7173 7298 7382
rect 7557 7379 7623 7382
rect 7741 7442 7807 7445
rect 8661 7442 8727 7445
rect 14000 7442 34000 7472
rect 7741 7440 8218 7442
rect 7741 7384 7746 7440
rect 7802 7384 8218 7440
rect 7741 7382 8218 7384
rect 7741 7379 7807 7382
rect 7649 7306 7715 7309
rect 8017 7306 8083 7309
rect 7649 7304 8083 7306
rect 7649 7248 7654 7304
rect 7710 7248 8022 7304
rect 8078 7248 8083 7304
rect 7649 7246 8083 7248
rect 7649 7243 7715 7246
rect 8017 7243 8083 7246
rect 7189 7168 7298 7173
rect 8158 7170 8218 7382
rect 8661 7440 34000 7442
rect 8661 7384 8666 7440
rect 8722 7384 34000 7440
rect 8661 7382 34000 7384
rect 8661 7379 8727 7382
rect 14000 7352 34000 7382
rect 7189 7112 7194 7168
rect 7250 7112 7298 7168
rect 7189 7110 7298 7112
rect 7974 7110 8218 7170
rect 7189 7107 7255 7110
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 7560 7104 7880 7105
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 7039 7880 7040
rect 7833 6898 7899 6901
rect 7974 6898 8034 7110
rect 8109 7034 8175 7037
rect 14000 7034 34000 7064
rect 8109 7032 34000 7034
rect 8109 6976 8114 7032
rect 8170 6976 34000 7032
rect 8109 6974 34000 6976
rect 8109 6971 8175 6974
rect 14000 6944 34000 6974
rect 7833 6896 8034 6898
rect 7833 6840 7838 6896
rect 7894 6840 8034 6896
rect 7833 6838 8034 6840
rect 7833 6835 7899 6838
rect 7974 6626 8034 6838
rect 8477 6626 8543 6629
rect 7974 6624 8543 6626
rect 7974 6568 8482 6624
rect 8538 6568 8543 6624
rect 7974 6566 8543 6568
rect 8477 6563 8543 6566
rect 13721 6626 13787 6629
rect 14000 6626 34000 6656
rect 13721 6624 34000 6626
rect 13721 6568 13726 6624
rect 13782 6568 34000 6624
rect 13721 6566 34000 6568
rect 13721 6563 13787 6566
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6566
rect 5060 6495 5380 6496
rect 9029 6218 9095 6221
rect 14000 6218 34000 6248
rect 9029 6216 34000 6218
rect 9029 6160 9034 6216
rect 9090 6160 34000 6216
rect 9029 6158 34000 6160
rect 9029 6155 9095 6158
rect 14000 6128 34000 6158
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 7560 6016 7880 6017
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5951 7880 5952
rect 13721 5810 13787 5813
rect 14000 5810 34000 5840
rect 13721 5808 34000 5810
rect 13721 5752 13726 5808
rect 13782 5752 34000 5808
rect 13721 5750 34000 5752
rect 13721 5747 13787 5750
rect 14000 5720 34000 5750
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 5407 5380 5408
rect 8201 5402 8267 5405
rect 14000 5402 34000 5432
rect 8201 5400 34000 5402
rect 8201 5344 8206 5400
rect 8262 5344 34000 5400
rect 8201 5342 34000 5344
rect 8201 5339 8267 5342
rect 14000 5312 34000 5342
rect 7833 5130 7899 5133
rect 7833 5128 12450 5130
rect 7833 5072 7838 5128
rect 7894 5072 12450 5128
rect 7833 5070 12450 5072
rect 7833 5067 7899 5070
rect 12390 4994 12450 5070
rect 14000 4994 34000 5024
rect 12390 4934 34000 4994
rect 7560 4928 7880 4929
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 14000 4904 34000 4934
rect 7560 4863 7880 4864
rect 9489 4586 9555 4589
rect 14000 4586 34000 4616
rect 9489 4584 34000 4586
rect 9489 4528 9494 4584
rect 9550 4528 34000 4584
rect 9489 4526 34000 4528
rect 9489 4523 9555 4526
rect 14000 4496 34000 4526
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 4319 5380 4320
rect 4613 4178 4679 4181
rect 7741 4178 7807 4181
rect 4613 4176 7807 4178
rect 4613 4120 4618 4176
rect 4674 4120 7746 4176
rect 7802 4120 7807 4176
rect 4613 4118 7807 4120
rect 4613 4115 4679 4118
rect 7741 4115 7807 4118
rect 13813 4178 13879 4181
rect 14000 4178 34000 4208
rect 13813 4176 34000 4178
rect 13813 4120 13818 4176
rect 13874 4120 34000 4176
rect 13813 4118 34000 4120
rect 13813 4115 13879 4118
rect 14000 4088 34000 4118
rect 7560 3840 7880 3841
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 3775 7880 3776
rect 9121 3770 9187 3773
rect 14000 3770 34000 3800
rect 9121 3768 34000 3770
rect 9121 3712 9126 3768
rect 9182 3712 34000 3768
rect 9121 3710 34000 3712
rect 9121 3707 9187 3710
rect 14000 3680 34000 3710
rect 2681 3438 2747 3441
rect 2484 3436 2747 3438
rect 2484 3380 2686 3436
rect 2742 3380 2747 3436
rect 2484 3378 2747 3380
rect 2681 3375 2747 3378
rect 6361 3362 6427 3365
rect 14000 3362 34000 3392
rect 6361 3360 34000 3362
rect 6361 3304 6366 3360
rect 6422 3304 34000 3360
rect 6361 3302 34000 3304
rect 6361 3299 6427 3302
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3302
rect 5060 3231 5380 3232
rect 13813 2954 13879 2957
rect 14000 2954 34000 2984
rect 13813 2952 34000 2954
rect 13813 2896 13818 2952
rect 13874 2896 34000 2952
rect 13813 2894 34000 2896
rect 13813 2891 13879 2894
rect 14000 2864 34000 2894
rect 7560 2752 7880 2753
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 2687 7880 2688
rect 14000 2546 34000 2576
rect 6870 2486 34000 2546
rect 6361 2410 6427 2413
rect 6870 2410 6930 2486
rect 14000 2456 34000 2486
rect 6361 2408 6930 2410
rect 6361 2352 6366 2408
rect 6422 2352 6930 2408
rect 6361 2350 6930 2352
rect 6361 2347 6427 2350
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 2143 5380 2144
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 8845 1730 8911 1733
rect 14000 1730 34000 1760
rect 8845 1728 34000 1730
rect 8845 1672 8850 1728
rect 8906 1672 34000 1728
rect 8845 1670 34000 1672
rect 8845 1667 8911 1670
rect 7560 1664 7880 1665
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 14000 1640 34000 1670
rect 7560 1599 7880 1600
rect 13813 1322 13879 1325
rect 14000 1322 34000 1352
rect 13813 1320 34000 1322
rect 13813 1264 13818 1320
rect 13874 1264 34000 1320
rect 13813 1262 34000 1264
rect 13813 1259 13879 1262
rect 14000 1232 34000 1262
rect 5060 1120 5380 1121
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1055 5380 1056
rect 9397 914 9463 917
rect 14000 914 34000 944
rect 9397 912 34000 914
rect 9397 856 9402 912
rect 9458 856 34000 912
rect 9397 854 34000 856
rect 9397 851 9463 854
rect 14000 824 34000 854
rect 9489 506 9555 509
rect 14000 506 34000 536
rect 9489 504 34000 506
rect 9489 448 9494 504
rect 9550 448 34000 504
rect 9489 446 34000 448
rect 9489 443 9555 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 5060 10912 5380 11472
rect 7560 11456 7880 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 6060 10956 6380 11424
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1088 6380 3960
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 5060 1040 5380 1056
rect 7560 1040 7880 1222
rect 8560 9266 8880 11424
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1088 8880 2270
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 6102 10956
rect 6338 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 5102 9908
rect 5338 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 6102 7576
rect 6338 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 5102 6528
rect 5338 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 5102 3148
rect 5338 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B
timestamp 1648946573
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A2
timestamp 1648946573
transform -1 0 8004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1648946573
transform -1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1648946573
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1648946573
transform -1 0 8740 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1648946573
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1648946573
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__B
timestamp 1648946573
transform -1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1648946573
transform 1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B_N
timestamp 1648946573
transform 1 0 1288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__B
timestamp 1648946573
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__B_N
timestamp 1648946573
transform -1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__B
timestamp 1648946573
transform -1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B_N
timestamp 1648946573
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B
timestamp 1648946573
transform -1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B_N
timestamp 1648946573
transform -1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B
timestamp 1648946573
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__B_N
timestamp 1648946573
transform 1 0 3864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B
timestamp 1648946573
transform -1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__B_N
timestamp 1648946573
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__B
timestamp 1648946573
transform -1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B_N
timestamp 1648946573
transform -1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__B
timestamp 1648946573
transform -1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__B_N
timestamp 1648946573
transform 1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B
timestamp 1648946573
transform -1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B_N
timestamp 1648946573
transform -1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 1648946573
transform -1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B_N
timestamp 1648946573
transform -1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__B
timestamp 1648946573
transform -1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B_N
timestamp 1648946573
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1648946573
transform -1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__B_N
timestamp 1648946573
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B
timestamp 1648946573
transform -1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B_N
timestamp 1648946573
transform -1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1648946573
transform -1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__RESET_B
timestamp 1648946573
transform -1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__RESET_B
timestamp 1648946573
transform -1 0 1472 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__RESET_B
timestamp 1648946573
transform 1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__RESET_B
timestamp 1648946573
transform -1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__RESET_B
timestamp 1648946573
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__RESET_B
timestamp 1648946573
transform 1 0 5244 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__RESET_B
timestamp 1648946573
transform 1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__RESET_B
timestamp 1648946573
transform 1 0 5888 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__RESET_B
timestamp 1648946573
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__RESET_B
timestamp 1648946573
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__RESET_B
timestamp 1648946573
transform -1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__RESET_B
timestamp 1648946573
transform -1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__RESET_B
timestamp 1648946573
transform 1 0 5704 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1648946573
transform -1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1648946573
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1648946573
transform -1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1648946573
transform -1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 7544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 3312 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 4048 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1648946573
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82
timestamp 1648946573
transform 1 0 8464 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1648946573
transform 1 0 9476 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1648946573
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26
timestamp 1648946573
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1648946573
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1648946573
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1648946573
transform 1 0 3312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1648946573
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1648946573
transform 1 0 8096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1648946573
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1648946573
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1648946573
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1648946573
transform 1 0 3404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1648946573
transform 1 0 3128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1648946573
transform 1 0 6440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1648946573
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1648946573
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1648946573
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_69
timestamp 1648946573
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1648946573
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1648946573
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1648946573
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1648946573
transform 1 0 3128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1648946573
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1648946573
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1648946573
transform 1 0 3404 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1648946573
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1648946573
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 1196 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1648946573
transform 1 0 3404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_31
timestamp 1648946573
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_61
timestamp 1648946573
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_80
timestamp 1648946573
transform 1 0 8280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1648946573
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1648946573
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1648946573
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1648946573
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1648946573
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1648946573
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1648946573
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1648946573
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1648946573
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1648946573
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1648946573
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1648946573
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1648946573
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1648946573
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1648946573
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1648946573
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1648946573
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1648946573
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1648946573
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1648946573
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1648946573
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1648946573
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1648946573
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1648946573
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1648946573
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1648946573
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1648946573
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1648946573
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1648946573
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1648946573
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1648946573
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1648946573
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1648946573
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1648946573
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1648946573
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1648946573
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1648946573
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1648946573
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1648946573
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1648946573
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1648946573
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1648946573
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1648946573
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1648946573
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1648946573
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1648946573
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1648946573
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1648946573
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1648946573
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1648946573
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1648946573
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1648946573
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1648946573
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1648946573
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1648946573
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1648946573
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1648946573
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1648946573
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1648946573
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1648946573
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1648946573
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1648946573
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1648946573
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1648946573
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_2  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8004 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1648946573
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9384 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 8648 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1648946573
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 8188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1648946573
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1648946573
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 2484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _111_
timestamp 1648946573
transform 1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1648946573
transform -1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113__4
timestamp 1648946573
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1648946573
transform 1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _115_
timestamp 1648946573
transform -1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _116_
timestamp 1648946573
transform -1 0 3404 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp 1648946573
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _118_
timestamp 1648946573
transform 1 0 2760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1648946573
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__5
timestamp 1648946573
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _121_
timestamp 1648946573
transform 1 0 3588 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1648946573
transform -1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _123_
timestamp 1648946573
transform -1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _124_
timestamp 1648946573
transform 1 0 6164 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1648946573
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126__6
timestamp 1648946573
transform -1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _127_
timestamp 1648946573
transform 1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1648946573
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _129_
timestamp 1648946573
transform 1 0 4968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1648946573
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131__7
timestamp 1648946573
transform 1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _132_
timestamp 1648946573
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _133_
timestamp 1648946573
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _134_
timestamp 1648946573
transform 1 0 4508 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1648946573
transform -1 0 5704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__8
timestamp 1648946573
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _137_
timestamp 1648946573
transform 1 0 4416 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1648946573
transform 1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _139_
timestamp 1648946573
transform 1 0 5152 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp 1648946573
transform -1 0 6440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1648946573
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142__9
timestamp 1648946573
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1648946573
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _144_
timestamp 1648946573
transform -1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1648946573
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _146_
timestamp 1648946573
transform 1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1648946573
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__10
timestamp 1648946573
transform -1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _149_
timestamp 1648946573
transform 1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1648946573
transform -1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp 1648946573
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _152_
timestamp 1648946573
transform 1 0 7360 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1648946573
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154__11
timestamp 1648946573
transform 1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _155_
timestamp 1648946573
transform 1 0 5980 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1648946573
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _157_
timestamp 1648946573
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1648946573
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159__12
timestamp 1648946573
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _160_
timestamp 1648946573
transform 1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1648946573
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _162_
timestamp 1648946573
transform 1 0 7636 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1648946573
transform -1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164__13
timestamp 1648946573
transform -1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _165_
timestamp 1648946573
transform -1 0 8648 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _166_
timestamp 1648946573
transform -1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _167_
timestamp 1648946573
transform -1 0 5428 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1648946573
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169__1
timestamp 1648946573
transform -1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _170_
timestamp 1648946573
transform 1 0 3680 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1648946573
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _172_
timestamp 1648946573
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1648946573
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__2
timestamp 1648946573
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _175_
timestamp 1648946573
transform 1 0 4324 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1648946573
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _177_
timestamp 1648946573
transform 1 0 5152 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _178_
timestamp 1648946573
transform -1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179__3
timestamp 1648946573
transform 1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _180_
timestamp 1648946573
transform -1 0 5152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1648946573
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 1840 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _183_
timestamp 1648946573
transform 1 0 1840 0 -1 8704
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _184_
timestamp 1648946573
transform 1 0 6072 0 1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _185_
timestamp 1648946573
transform 1 0 6900 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _186_
timestamp 1648946573
transform 1 0 3496 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _187_
timestamp 1648946573
transform 1 0 3312 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _188_
timestamp 1648946573
transform 1 0 3496 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _189_
timestamp 1648946573
transform 1 0 6532 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _190_
timestamp 1648946573
transform 1 0 6440 0 1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _191_
timestamp 1648946573
transform 1 0 6716 0 1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _192_
timestamp 1648946573
transform 1 0 3588 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _193_
timestamp 1648946573
transform 1 0 4232 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _194_
timestamp 1648946573
transform 1 0 5704 0 1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 3128 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _196_
timestamp 1648946573
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _197_
timestamp 1648946573
transform -1 0 3128 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _198_
timestamp 1648946573
transform 1 0 1472 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _199_
timestamp 1648946573
transform -1 0 3496 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _200_
timestamp 1648946573
transform 1 0 3312 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _201_
timestamp 1648946573
transform -1 0 5244 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _202_
timestamp 1648946573
transform 1 0 4232 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _203_
timestamp 1648946573
transform 1 0 6164 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _204_
timestamp 1648946573
transform 1 0 6164 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _205_
timestamp 1648946573
transform 1 0 7360 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _206_
timestamp 1648946573
transform -1 0 7728 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _207_
timestamp 1648946573
transform 1 0 6256 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _209_
timestamp 1648946573
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _210_
timestamp 1648946573
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5152 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__077_
timestamp 1648946573
transform 1 0 4232 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1648946573
transform -1 0 8004 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1648946573
transform -1 0 8004 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__077_
timestamp 1648946573
transform 1 0 1472 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock
timestamp 1648946573
transform -1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_load
timestamp 1648946573
transform -1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__049_
timestamp 1648946573
transform -1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__077_
timestamp 1648946573
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1648946573
transform -1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_load
timestamp 1648946573
transform -1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd2_1  data_delay_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8280 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd2_1  data_delay_2
timestamp 1648946573
transform -1 0 9568 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 4416 0 1 5440
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 1638030917
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1648946573
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1648946573
transform 1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1648946573
transform 1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1648946573
transform 1 0 1288 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1648946573
transform 1 0 1288 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1648946573
transform 1 0 3588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1648946573
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1648946573
transform -1 0 5796 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1648946573
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1648946573
transform 1 0 3588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1648946573
transform -1 0 9476 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1648946573
transform 1 0 4416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1648946573
transform 1 0 2024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1648946573
transform 1 0 2024 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1648946573
transform -1 0 9476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1648946573
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1648946573
transform -1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1648946573
transform 1 0 6624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1648946573
transform -1 0 6808 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1648946573
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1648946573
transform 1 0 6808 0 1 1088
box -38 -48 774 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
