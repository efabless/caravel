* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_363_ _348_/X ext_trim[2] _398_/B _362_/Y VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__a211o_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_294_ _397_/A _325_/A VGND VGND VPWR VPWR _313_/A sky130_fd_sc_hd__xnor2_2
X_432_ _437_/A _433_/B VGND VGND VPWR VPWR _432_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_415_ _376_/A _370_/A _468_/Q VGND VGND VPWR VPWR _416_/B sky130_fd_sc_hd__o21ai_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_346_ _346_/A VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__buf_2
X_277_ _420_/B _302_/A VGND VGND VPWR VPWR _278_/D sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _423_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_329_ _463_/Q _291_/X _328_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__o21a_2
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__392__A2 ext_trim[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__383__A2 ext_trim[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _385_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _383_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_362_ _397_/A _438_/A VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__nor2_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _293_/A VGND VGND VPWR VPWR _328_/B sky130_fd_sc_hd__buf_2
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_431_ _437_/A _433_/B VGND VGND VPWR VPWR _431_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__410__A1 _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_414_ _406_/B _359_/A _371_/Y _403_/B _413_/X VGND VGND VPWR VPWR _414_/X sky130_fd_sc_hd__o2111a_2
X_276_ _465_/Q VGND VGND VPWR VPWR _302_/A sky130_fd_sc_hd__inv_2
X_345_ _455_/Q _456_/Q _345_/S VGND VGND VPWR VPWR _346_/A sky130_fd_sc_hd__mux2_2
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ _463_/Q _328_/B VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_259_ _288_/B _288_/C _258_/X VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__a21o_2
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _421_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _422_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _367_/A dco VGND VGND VPWR VPWR _398_/B sky130_fd_sc_hd__nor2_2
X_292_ _397_/A _325_/A _278_/Y _291_/X VGND VGND VPWR VPWR _293_/A sky130_fd_sc_hd__o31a_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_430_ _437_/A _433_/B VGND VGND VPWR VPWR _430_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_413_ _301_/Y _367_/Y _386_/Y _412_/X VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__o211a_2
X_275_ _466_/Q VGND VGND VPWR VPWR _420_/B sky130_fd_sc_hd__inv_2
X_344_ _344_/A VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__buf_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__410__A2 ext_trim[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _369_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_327_ _327_/A VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__buf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258_ div[1] _258_/B VGND VGND VPWR VPWR _258_/X sky130_fd_sc_hd__and2_2
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _373_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_360_ _352_/X ext_trim[1] _403_/A VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__a21o_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_291_ _285_/X _291_/B _291_/C VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__and3b_2
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__244__A div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_412_ _420_/B _283_/B _381_/A _376_/Y VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__o22a_2
X_274_ _464_/Q _463_/Q VGND VGND VPWR VPWR _324_/B sky130_fd_sc_hd__and2_2
X_343_ _456_/Q _457_/Q _345_/S VGND VGND VPWR VPWR _344_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _409_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_326_ _464_/Q _325_/X _328_/B VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__mux2_2
X_257_ div[0] _257_/B _257_/C VGND VGND VPWR VPWR _288_/C sky130_fd_sc_hd__nand3b_2
X_309_ _309_/A _309_/B VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__and2_2
XANTENNA__252__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__427__A _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _410_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__350__A ext_trim[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ _266_/X _290_/B _290_/C _290_/D VGND VGND VPWR VPWR _291_/C sky130_fd_sc_hd__nand4b_2
XANTENNA__422__A1 _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__404__A1 _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_411_ _379_/X ext_trim[19] _403_/A _403_/B VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__a22o_2
X_273_ _467_/Q VGND VGND VPWR VPWR _376_/A sky130_fd_sc_hd__buf_2
X_342_ _342_/A _347_/B _342_/C VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__nand3_2
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ _325_/A _325_/B VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_256_ _256_/A VGND VGND VPWR VPWR _257_/C sky130_fd_sc_hd__inv_2
X_308_ _420_/A _325_/A VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__xnor2_2
X_239_ _262_/A _239_/B VGND VGND VPWR VPWR _240_/C sky130_fd_sc_hd__nand2b_2
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__348__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__258__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__422__A2 ext_trim[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_410_ _428_/A ext_trim[18] _398_/X VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _360_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XANTENNA__404__A2 ext_trim[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_272_ _302_/B VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__buf_2
X_341_ _342_/C _340_/Y _347_/B VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__a21boi_2
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__266__A div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_255_ _342_/A _473_/Q VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ _324_/A _324_/B VGND VGND VPWR VPWR _325_/B sky130_fd_sc_hd__nor2_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_307_ _313_/A _316_/A _316_/B _398_/A _325_/A VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__a32o_2
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_238_ _461_/Q _476_/Q VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__nand2_2
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__361__B dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _396_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_271_ _260_/X _266_/X _267_/X _290_/C VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__o31a_2
X_340_ _459_/Q _342_/A VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _360_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_469_ _477_/CLK _469_/D _445_/Y VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__389__A2 ext_trim[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_323_ _328_/B _322_/Y _465_/Q _291_/X VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__o2bb2a_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_254_ _342_/A _473_/Q VGND VGND VPWR VPWR _257_/B sky130_fd_sc_hd__nand2_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_306_ _401_/B VGND VGND VPWR VPWR _398_/A sky130_fd_sc_hd__inv_2
X_237_ _461_/Q _476_/Q VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__289__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ div[4] _266_/B _268_/Y _269_/Y VGND VGND VPWR VPWR _290_/C sky130_fd_sc_hd__o211a_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_399_ _379_/X ext_trim[15] _397_/Y _398_/X VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _396_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_468_ _477_/CLK _468_/D _444_/Y VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _322_/A _322_/B VGND VGND VPWR VPWR _322_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_253_ _258_/B _253_/B VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__nand2b_2
X_305_ _301_/Y _322_/A _322_/B _406_/C _325_/A VGND VGND VPWR VPWR _316_/B sky130_fd_sc_hd__a32o_2
X_236_ _251_/A _251_/B _247_/B _235_/X VGND VGND VPWR VPWR _240_/B sky130_fd_sc_hd__a211o_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _461_/Q _476_/Q _345_/S VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _383_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_398_ _398_/A _398_/B VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__and2_2
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_467_ _477_/CLK _467_/D _442_/Y VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_321_ _420_/B _321_/B VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__xnor2_2
X_252_ div[1] VGND VGND VPWR VPWR _253_/B sky130_fd_sc_hd__inv_2
X_304_ _302_/B _303_/Y _324_/B VGND VGND VPWR VPWR _322_/B sky130_fd_sc_hd__a21o_2
X_235_ _459_/Q _474_/Q VGND VGND VPWR VPWR _235_/X sky130_fd_sc_hd__and2_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ _218_/A VGND VGND VPWR VPWR _477_/D sky130_fd_sc_hd__buf_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _421_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__270__A1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_397_ _397_/A _397_/B VGND VGND VPWR VPWR _397_/Y sky130_fd_sc_hd__nand2_2
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_466_ _477_/CLK _466_/D _441_/Y VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfrtp_2
X_320_ _302_/A _322_/B _319_/X _293_/A VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__o211a_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_251_ _251_/A _251_/B VGND VGND VPWR VPWR _258_/B sky130_fd_sc_hd__xnor2_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_449_ _454_/A _451_/B VGND VGND VPWR VPWR _449_/Y sky130_fd_sc_hd__nor2_2
X_303_ _324_/A VGND VGND VPWR VPWR _303_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_234_ _460_/Q _475_/Q VGND VGND VPWR VPWR _247_/B sky130_fd_sc_hd__and2_2
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _433_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__470__D osc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_217_ _462_/Q _477_/Q _347_/B VGND VGND VPWR VPWR _218_/A sky130_fd_sc_hd__mux2_2
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__419__A1 _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _380_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_396_ _379_/X ext_trim[14] _372_/X _395_/X VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__a22o_2
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_465_ _477_/CLK _465_/D _440_/Y VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_250_ _250_/A _250_/B VGND VGND VPWR VPWR _250_/Y sky130_fd_sc_hd__nand2_2
X_379_ dco VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__buf_2
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_448_ _454_/A _451_/B VGND VGND VPWR VPWR _448_/Y sky130_fd_sc_hd__nor2_2
X_302_ _302_/A _302_/B VGND VGND VPWR VPWR _322_/A sky130_fd_sc_hd__xnor2_2
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_233_ _459_/Q _474_/Q VGND VGND VPWR VPWR _251_/B sky130_fd_sc_hd__xor2_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ _345_/S VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__buf_2
XANTENNA__419__A2 ext_trim[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_464_ _477_/CLK _464_/D _439_/Y VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _419_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_395_ _376_/B _395_/B _395_/C VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__and3b_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_378_ _352_/X ext_trim[7] _377_/X VGND VGND VPWR VPWR _378_/X sky130_fd_sc_hd__a21o_2
X_447_ dco VGND VGND VPWR VPWR _454_/A sky130_fd_sc_hd__buf_2
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_301_ _406_/C _381_/A VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__nand2_2
X_232_ _458_/Q _473_/Q VGND VGND VPWR VPWR _251_/A sky130_fd_sc_hd__and2_2
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _375_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__373__A2 ext_trim[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_215_ _215_/A VGND VGND VPWR VPWR _345_/S sky130_fd_sc_hd__buf_2
XANTENNA__364__A2 ext_trim[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _420_/A _278_/D _420_/C VGND VGND VPWR VPWR _395_/C sky130_fd_sc_hd__o21ai_2
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_463_ _477_/CLK _463_/D _437_/Y VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_2
X_377_ _406_/C _376_/Y _403_/A VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__o21a_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_446_ _446_/A _451_/B VGND VGND VPWR VPWR _446_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _369_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_300_ _370_/A _465_/Q VGND VGND VPWR VPWR _381_/A sky130_fd_sc_hd__nand2_2
X_231_ _460_/Q _231_/B VGND VGND VPWR VPWR _240_/A sky130_fd_sc_hd__nand2b_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_429_ _438_/A VGND VGND VPWR VPWR _437_/A sky130_fd_sc_hd__buf_2
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _385_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _411_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_214_ _472_/D _472_/Q VGND VGND VPWR VPWR _215_/A sky130_fd_sc_hd__xnor2_2
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_393_ _468_/Q _406_/C _376_/A _367_/A VGND VGND VPWR VPWR _395_/B sky130_fd_sc_hd__a211o_2
X_462_ _477_/CLK _462_/D _436_/Y VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _409_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_376_ _376_/A _376_/B VGND VGND VPWR VPWR _376_/Y sky130_fd_sc_hd__nand2_2
X_445_ _446_/A _451_/B VGND VGND VPWR VPWR _445_/Y sky130_fd_sc_hd__nor2_2
X_230_ _475_/Q VGND VGND VPWR VPWR _231_/B sky130_fd_sc_hd__inv_2
X_359_ _359_/A _359_/B VGND VGND VPWR VPWR _403_/A sky130_fd_sc_hd__and2_2
X_428_ _428_/A _433_/B VGND VGND VPWR VPWR _428_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _422_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__421__B1 ext_trim[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_392_ _428_/A ext_trim[13] _391_/X VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__a21o_2
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_461_ _477_/CLK _461_/D _435_/Y VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ _352_/X ext_trim[6] _374_/Y VGND VGND VPWR VPWR _375_/X sky130_fd_sc_hd__a21o_2
X_444_ _446_/A _451_/B VGND VGND VPWR VPWR _444_/Y sky130_fd_sc_hd__nor2_2
X_358_ dco _358_/B VGND VGND VPWR VPWR _359_/B sky130_fd_sc_hd__nor2_2
X_427_ _428_/A _433_/B VGND VGND VPWR VPWR _427_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ div[3] _242_/Y _249_/X _250_/Y VGND VGND VPWR VPWR _290_/D sky130_fd_sc_hd__o211a_2
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _351_/Y VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__267__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__425__A enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_391_ _370_/A _376_/Y _403_/A VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__o21a_2
X_460_ _477_/CLK _460_/D _433_/Y VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_374_ _420_/B _358_/B dco VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_443_ _454_/B VGND VGND VPWR VPWR _451_/B sky130_fd_sc_hd__buf_2
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _364_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_357_ _469_/Q _398_/A VGND VGND VPWR VPWR _358_/B sky130_fd_sc_hd__nor2_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _258_/X _288_/B _288_/C _288_/D VGND VGND VPWR VPWR _290_/B sky130_fd_sc_hd__and4b_2
X_426_ _454_/B VGND VGND VPWR VPWR _433_/B sky130_fd_sc_hd__buf_2
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _392_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_409_ _405_/Y _407_/X _408_/X ext_trim[17] _348_/X VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__a32o_2
XANTENNA__428__A _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_8
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ringosc.dstage\[0\].id.delaybuf0_A ringosc.ibufp00/A VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__425__B resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ _438_/A VGND VGND VPWR VPWR _428_/A sky130_fd_sc_hd__buf_2
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_373_ _352_/X ext_trim[5] _372_/X VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__a21o_2
X_442_ _446_/A _442_/B VGND VGND VPWR VPWR _442_/Y sky130_fd_sc_hd__nor2_2
X_356_ _386_/B _371_/B VGND VGND VPWR VPWR _359_/A sky130_fd_sc_hd__nor2_2
X_287_ _251_/A _256_/A div[0] VGND VGND VPWR VPWR _288_/D sky130_fd_sc_hd__o21ai_2
X_425_ enable resetb VGND VGND VPWR VPWR _454_/B sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _404_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _420_/B _365_/Y _401_/Y _406_/B _403_/B VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__o221a_2
X_339_ _339_/A VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__buf_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _424_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__349__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_372_ _301_/Y _367_/Y _359_/B _371_/Y VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__o211a_2
X_441_ _446_/A _442_/B VGND VGND VPWR VPWR _441_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__447__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_355_ _367_/A _397_/A _467_/Q VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__and3_2
X_424_ _379_/X ext_trim[25] _403_/X _407_/C VGND VGND VPWR VPWR _424_/X sky130_fd_sc_hd__a22o_2
X_286_ _215_/A _455_/Q _457_/Q _456_/Q VGND VGND VPWR VPWR _291_/B sky130_fd_sc_hd__and4b_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _407_/A _407_/B _407_/C VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__and3_2
X_269_ _462_/Q _477_/Q VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__nand2_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_338_ _347_/B _338_/B VGND VGND VPWR VPWR _339_/A sky130_fd_sc_hd__and2_2
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_371_ _397_/B _371_/B VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__nand2_2
X_440_ _446_/A _442_/B VGND VGND VPWR VPWR _440_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ _467_/Q _376_/B VGND VGND VPWR VPWR _386_/B sky130_fd_sc_hd__and2b_2
X_423_ _379_/X ext_trim[24] _362_/Y _420_/A VGND VGND VPWR VPWR _423_/X sky130_fd_sc_hd__a22o_2
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_285_ _302_/B _285_/B _324_/A VGND VGND VPWR VPWR _285_/X sky130_fd_sc_hd__and3_2
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_406_ _401_/Y _406_/B _406_/C VGND VGND VPWR VPWR _407_/C sky130_fd_sc_hd__nand3b_2
X_268_ _268_/A _268_/B VGND VGND VPWR VPWR _268_/Y sky130_fd_sc_hd__nand2_2
X_337_ _331_/B _335_/Y _342_/C VGND VGND VPWR VPWR _338_/B sky130_fd_sc_hd__o21ai_2
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__424__A2 ext_trim[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_370_ _370_/A _465_/Q VGND VGND VPWR VPWR _397_/B sky130_fd_sc_hd__nor2_2
X_353_ _469_/Q _397_/A VGND VGND VPWR VPWR _376_/B sky130_fd_sc_hd__nor2_2
X_422_ _428_/A ext_trim[23] _398_/B VGND VGND VPWR VPWR _422_/X sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _351_/Y VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_284_ _464_/Q _463_/Q VGND VGND VPWR VPWR _324_/A sky130_fd_sc_hd__nor2_2
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _378_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_405_ _420_/A _406_/B _420_/C VGND VGND VPWR VPWR _405_/Y sky130_fd_sc_hd__nand3_2
X_267_ div[3] _242_/Y _249_/X VGND VGND VPWR VPWR _267_/X sky130_fd_sc_hd__o21ba_2
X_336_ _462_/Q _336_/B VGND VGND VPWR VPWR _342_/C sky130_fd_sc_hd__nand2_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__379__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__409__B1 ext_trim[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__360__A2 ext_trim[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ _465_/Q _324_/A _325_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__260__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_421_ _407_/X _408_/X _420_/Y ext_trim[22] _348_/X VGND VGND VPWR VPWR _421_/X sky130_fd_sc_hd__a32o_2
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _392_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _438_/A VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__buf_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_283_ _298_/A _283_/B VGND VGND VPWR VPWR _285_/B sky130_fd_sc_hd__nor2_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _417_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_404_ _428_/A ext_trim[16] _403_/X VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__a21o_2
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_266_ div[4] _266_/B VGND VGND VPWR VPWR _266_/X sky130_fd_sc_hd__and2_2
X_335_ _459_/Q _342_/A _460_/Q VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_318_ _318_/A VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__buf_2
X_249_ _243_/Y _242_/A _242_/B _250_/A _250_/B VGND VGND VPWR VPWR _249_/X sky130_fd_sc_hd__o32a_2
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _380_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclockp_buffer_0 _477_/CLK VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_16
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ringosc.ibufp00_A ringosc.ibufp00/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_420_ _420_/A _420_/B _420_/C VGND VGND VPWR VPWR _420_/Y sky130_fd_sc_hd__nand3_2
X_282_ _367_/A _401_/B VGND VGND VPWR VPWR _283_/B sky130_fd_sc_hd__nand2_2
X_351_ _348_/X _285_/B _350_/Y VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _403_/A _403_/B _407_/B VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__and3_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_334_ _461_/Q _331_/B _333_/Y _347_/B VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__o211a_2
X_265_ _268_/A _268_/B VGND VGND VPWR VPWR _266_/B sky130_fd_sc_hd__xnor2_2
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_317_ _376_/A _316_/X _328_/B VGND VGND VPWR VPWR _318_/A sky130_fd_sc_hd__mux2_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_248_ _248_/A _248_/B VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _364_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _419_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
Xclockp_buffer_1 ringosc.ibufp11/Y VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_16
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__384__A_N ext_trim[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_281_ _468_/Q _467_/Q VGND VGND VPWR VPWR _401_/B sky130_fd_sc_hd__nor2_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_350_ ext_trim[0] _438_/A VGND VGND VPWR VPWR _350_/Y sky130_fd_sc_hd__nand2_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__257__A_N div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ _381_/A _376_/Y _401_/Y _406_/C VGND VGND VPWR VPWR _407_/B sky130_fd_sc_hd__o22a_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ _462_/Q _336_/B VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__nand2b_2
X_264_ _262_/Y _240_/A _240_/B _263_/X VGND VGND VPWR VPWR _268_/B sky130_fd_sc_hd__a31o_2
XANTENNA__363__A2 ext_trim[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_316_ _316_/A _316_/B VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__xor2_2
X_247_ _247_/A _247_/B VGND VGND VPWR VPWR _248_/B sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _404_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ _469_/Q VGND VGND VPWR VPWR _367_/A sky130_fd_sc_hd__inv_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_401_ _469_/Q _401_/B VGND VGND VPWR VPWR _401_/Y sky130_fd_sc_hd__nand2_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _462_/Q _336_/B _347_/B VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__o21a_2
X_263_ _461_/Q _476_/Q VGND VGND VPWR VPWR _263_/X sky130_fd_sc_hd__and2_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_246_ _460_/Q _475_/Q VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__nor2_2
X_315_ _315_/A VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__buf_2
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _468_/Q VGND VGND VPWR VPWR _397_/A sky130_fd_sc_hd__inv_2
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__clkinv_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_477_ _477_/CLK _477_/D _454_/Y VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _376_/Y _406_/B VGND VGND VPWR VPWR _403_/B sky130_fd_sc_hd__nand2b_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _262_/A VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_331_ _461_/Q _331_/B VGND VGND VPWR VPWR _336_/B sky130_fd_sc_hd__and2_2
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _468_/Q _313_/Y _328_/B VGND VGND VPWR VPWR _315_/A sky130_fd_sc_hd__mux2_2
X_245_ _251_/A _251_/B _235_/X VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _373_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_228_ _469_/Q VGND VGND VPWR VPWR _420_/A sky130_fd_sc_hd__buf_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__375__A2 ext_trim[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR ringosc.ibufp11/Y sky130_fd_sc_hd__clkinv_8
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ _477_/CLK _476_/D _453_/Y VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _462_/Q _477_/Q VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__xor2_2
X_330_ _460_/Q _459_/Q _342_/A VGND VGND VPWR VPWR _331_/B sky130_fd_sc_hd__and3_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_459_ _477_/CLK _459_/D _432_/Y VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_313_ _313_/A _313_/B VGND VGND VPWR VPWR _313_/Y sky130_fd_sc_hd__xnor2_2
X_244_ div[2] VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _410_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_227_ _227_/A VGND VGND VPWR VPWR _473_/D sky130_fd_sc_hd__buf_2
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__387__B1 ext_trim[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _477_/CLK sky130_fd_sc_hd__clkinv_8
X_475_ _477_/CLK _475_/D _452_/Y VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ div[3] _242_/Y _249_/X _250_/Y _259_/X VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__o2111a_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_389_ _352_/X ext_trim[12] _388_/X VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__a21o_2
XANTENNA__243__A div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_458_ _477_/CLK _458_/D _431_/Y VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_312_ _316_/A _316_/B _297_/B VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__a21oi_2
X_243_ div[3] VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _387_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_8
X_226_ _342_/A _473_/Q _345_/S VGND VGND VPWR VPWR _227_/A sky130_fd_sc_hd__mux2_2
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__411__A2 ext_trim[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_474_ _477_/CLK _474_/D _451_/Y VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__287__B1 div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ _370_/A _367_/Y _359_/B VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__o21a_2
X_457_ _477_/CLK _457_/D _430_/Y VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfrtp_2
X_311_ _420_/A _328_/B _309_/X _310_/Y VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__o22a_2
X_242_ _242_/A _242_/B VGND VGND VPWR VPWR _242_/Y sky130_fd_sc_hd__nor2_2
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _423_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_225_ _458_/Q VGND VGND VPWR VPWR _342_/A sky130_fd_sc_hd__buf_2
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__396__A2 ext_trim[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__378__A2 ext_trim[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__369__A2 ext_trim[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_473_ _477_/CLK _473_/D _450_/Y VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_387_ _367_/Y _359_/B _386_/Y ext_trim[11] _348_/X VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__a32o_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_456_ _477_/CLK _456_/D _428_/Y VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ _309_/A _309_/B _328_/B VGND VGND VPWR VPWR _310_/Y sky130_fd_sc_hd__o21ai_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _363_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_241_ _240_/A _240_/B _240_/C VGND VGND VPWR VPWR _242_/B sky130_fd_sc_hd__a21oi_2
X_439_ _446_/A _442_/B VGND VGND VPWR VPWR _439_/Y sky130_fd_sc_hd__nor2_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_224_ _224_/A VGND VGND VPWR VPWR _474_/D sky130_fd_sc_hd__buf_2
XFILLER_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _375_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_472_ _477_/CLK _472_/D _449_/Y VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__358__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_386_ _406_/B _386_/B VGND VGND VPWR VPWR _386_/Y sky130_fd_sc_hd__nand2_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_455_ _477_/CLK _455_/D _427_/Y VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _399_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__423__A2 ext_trim[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _240_/A _240_/B _240_/C VGND VGND VPWR VPWR _242_/A sky130_fd_sc_hd__and3_2
X_369_ _352_/X ext_trim[4] _407_/A VGND VGND VPWR VPWR _369_/X sky130_fd_sc_hd__a21o_2
X_438_ _438_/A VGND VGND VPWR VPWR _446_/A sky130_fd_sc_hd__buf_2
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_223_ _459_/Q _474_/Q _345_/S VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__mux2_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _411_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_471_ _477_/CLK _471_/D _448_/Y VGND VGND VPWR VPWR _472_/D sky130_fd_sc_hd__dfrtp_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_385_ _348_/X _283_/B _278_/D _384_/Y VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__o31a_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _389_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_2
X_454_ _454_/A _454_/B VGND VGND VPWR VPWR _454_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__417__B1 ext_trim[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_368_ _370_/A _365_/Y _367_/Y _359_/B VGND VGND VPWR VPWR _407_/A sky130_fd_sc_hd__o211a_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ _466_/Q VGND VGND VPWR VPWR _370_/A sky130_fd_sc_hd__buf_2
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_437_ _437_/A _442_/B VGND VGND VPWR VPWR _437_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_222_ _222_/A VGND VGND VPWR VPWR _475_/D sky130_fd_sc_hd__buf_2
XANTENNA__399__A2 ext_trim[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _363_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_470_ _477_/CLK osc _446_/Y VGND VGND VPWR VPWR _471_/D sky130_fd_sc_hd__dfrtp_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ ext_trim[10] _438_/A VGND VGND VPWR VPWR _384_/Y sky130_fd_sc_hd__nand2b_2
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _424_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_2
X_453_ _454_/A _454_/B VGND VGND VPWR VPWR _453_/Y sky130_fd_sc_hd__nor2_2
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ _367_/A _420_/C VGND VGND VPWR VPWR _367_/Y sky130_fd_sc_hd__nand2_2
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_298_ _298_/A VGND VGND VPWR VPWR _406_/C sky130_fd_sc_hd__buf_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_436_ _437_/A _442_/B VGND VGND VPWR VPWR _436_/Y sky130_fd_sc_hd__nor2_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_221_ _460_/Q _475_/Q _345_/S VGND VGND VPWR VPWR _222_/A sky130_fd_sc_hd__mux2_2
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_419_ _428_/A ext_trim[21] _418_/X VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__a21o_2
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _399_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _379_/X ext_trim[9] _372_/X _382_/X VGND VGND VPWR VPWR _383_/X sky130_fd_sc_hd__a22o_2
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_452_ _454_/A _454_/B VGND VGND VPWR VPWR _452_/Y sky130_fd_sc_hd__nor2_2
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_366_ _397_/A _376_/A VGND VGND VPWR VPWR _420_/C sky130_fd_sc_hd__and2_2
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_297_ _297_/A _297_/B VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__nor2_2
X_435_ _437_/A _442_/B VGND VGND VPWR VPWR _435_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_220_ _220_/A VGND VGND VPWR VPWR _476_/D sky130_fd_sc_hd__buf_2
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_418_ _370_/A _302_/A _401_/Y _403_/X VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__o31a_2
X_349_ dco VGND VGND VPWR VPWR _438_/A sky130_fd_sc_hd__buf_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.ctrlen0 _433_/B _389_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__380__A2 ext_trim[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_382_ _406_/C _365_/Y _367_/Y _406_/B VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__o22a_2
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_451_ _454_/A _451_/B VGND VGND VPWR VPWR _451_/Y sky130_fd_sc_hd__nor2_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_365_ _386_/B VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__inv_2
X_296_ _467_/Q _302_/B VGND VGND VPWR VPWR _297_/B sky130_fd_sc_hd__and2_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_434_ _454_/B VGND VGND VPWR VPWR _442_/B sky130_fd_sc_hd__buf_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_417_ _374_/Y _414_/X _416_/Y ext_trim[20] _348_/X VGND VGND VPWR VPWR _417_/X sky130_fd_sc_hd__a32o_2
X_348_ dco VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__buf_2
X_279_ _420_/B _302_/A VGND VGND VPWR VPWR _298_/A sky130_fd_sc_hd__nand2_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _378_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__374__B1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_381_ _381_/A VGND VGND VPWR VPWR _406_/B sky130_fd_sc_hd__buf_2
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_450_ _454_/A _451_/B VGND VGND VPWR VPWR _450_/Y sky130_fd_sc_hd__nor2_2
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_433_ _437_/A _433_/B VGND VGND VPWR VPWR _433_/Y sky130_fd_sc_hd__nor2_2
X_364_ _352_/X ext_trim[3] _359_/B VGND VGND VPWR VPWR _364_/X sky130_fd_sc_hd__a21o_2
X_295_ _376_/A _302_/B VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__nor2_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_416_ _420_/A _416_/B VGND VGND VPWR VPWR _416_/Y sky130_fd_sc_hd__nand2_2
X_278_ _469_/Q _376_/A _324_/B _278_/D VGND VGND VPWR VPWR _278_/Y sky130_fd_sc_hd__nand4_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_347_ _455_/Q _347_/B VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__nand2b_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _387_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _417_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__392__A1 _428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_380_ _379_/X ext_trim[8] _359_/B _371_/Y VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__a22o_2
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

