module sky130_fd_sc_hd__conb_1 (
   output HI,
   output LO,
   input VPWR,
   input VGND,
   input VPB,
   input VNB
);
endmodule
