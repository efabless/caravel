* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 porb resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_432_ clknet_1_1__leaf_pll_clk _097_ net27 VGND VGND VPWR VPWR divider.odd_0.initial_begin\[2\]
+ sky130_fd_sc_hd__dfrtn_1
X_294_ _007_ _143_ _145_ net24 VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ divider.odd_0.initial_begin\[2\] _014_ _003_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__mux2_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__428__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_346_ _167_ divider2.odd_0.out_counter net23 VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__a21oi_1
X_415_ net40 net47 net31 VGND VGND VPWR VPWR reset_delay\[1\] sky130_fd_sc_hd__dfstp_1
X_277_ _130_ divider2.odd_0.counter2\[1\] VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__nand2_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_329_ divider2.odd_0.initial_begin\[1\] divider2.odd_0.initial_begin\[0\] VGND VGND
+ VPWR VPWR _061_ sky130_fd_sc_hd__xnor2_1
XANTENNA__312__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__037_ clknet_0__037_ VGND VGND VPWR VPWR clknet_1_1__leaf__037_ sky130_fd_sc_hd__clkbuf_16
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_362_ divider.odd_0.initial_begin\[0\] _012_ _003_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__mux2_1
X_431_ net38 _096_ net27 VGND VGND VPWR VPWR divider.odd_0.initial_begin\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ _140_ divider.odd_0.counter2\[1\] VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__nand2_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_345_ net14 net15 net16 divider2.odd_0.counter\[0\] _148_ VGND VGND VPWR VPWR _167_
+ sky130_fd_sc_hd__o2111ai_2
X_276_ net22 _130_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__nand2b_1
X_414_ net39 net44 net28 VGND VGND VPWR VPWR reset_delay\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__405__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__238__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_328_ net15 net16 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_292_ _143_ _144_ _122_ _141_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__o2bb2ai_1
X_361_ _124_ _142_ _178_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_430_ clknet_1_1__leaf_pll_clk _095_ net27 VGND VGND VPWR VPWR divider.odd_0.initial_begin\[0\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_275_ _127_ _128_ net22 VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a21oi_1
X_344_ net2 net3 net4 VGND VGND VPWR VPWR divider.even_0.resetb sky130_fd_sc_hd__and3b_1
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_258_ _006_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__inv_2
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ divider.even_0.counter\[1\] divider.even_0.counter\[0\] VGND VGND VPWR VPWR
+ _058_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__B1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_408__8 clknet_1_1__leaf_net11 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__inv_4
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_360_ net24 _140_ divider.odd_0.counter2\[2\] VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__nand3b_1
X_291_ _136_ _122_ divider.odd_0.counter2\[0\] net25 VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__a31o_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ divider2.even_0.counter\[1\] divider2.even_0.counter\[0\] VGND VGND VPWR VPWR
+ _078_ sky130_fd_sc_hd__xnor2_1
X_274_ _131_ _132_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__nand2_1
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_326_ _159_ _160_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_309_ divider2.odd_0.out_counter2 divider2.odd_0.out_counter VGND VGND VPWR VPWR
+ _153_ sky130_fd_sc_hd__and2_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_divider.out divider.out VGND VGND VPWR VPWR clknet_0_divider.out sky130_fd_sc_hd__clkbuf_1
XFILLER_19_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput12 net12 VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_12
XFILLER_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input8_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ net24 _140_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clknet_0_pll_clk sky130_fd_sc_hd__clkbuf_16
X_342_ _165_ _166_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nand2b_1
X_273_ _034_ _127_ _128_ _121_ net22 VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__a41oi_1
XANTENNA__331__B1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_325_ divider.odd_0.counter\[1\] divider.odd_0.counter\[0\] divider.odd_0.counter\[2\]
+ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_256_ reset_delay\[0\] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkinv_4
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_239_ _073_ net15 _035_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__mux2_1
X_308_ net17 _038_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand2b_2
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__286__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__A2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_pll_clk90 clknet_0_pll_clk90 VGND VGND VPWR VPWR clknet_1_0__leaf_pll_clk90
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_341_ divider2.odd_0.counter\[1\] divider2.odd_0.counter\[0\] divider2.odd_0.counter\[2\]
+ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__o21ai_1
X_272_ _034_ _127_ _128_ _121_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__a31o_1
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ divider.odd_0.counter\[1\] divider.odd_0.counter\[0\] divider.odd_0.counter\[2\]
+ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__nor3_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_255_ net1 VGND VGND VPWR VPWR pll_clk_sel sky130_fd_sc_hd__clkinv_4
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_238_ _072_ net16 net23 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__mux2_1
X_307_ _151_ _139_ _150_ _149_ VGND VGND VPWR VPWR divider.out sky130_fd_sc_hd__o31ai_1
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_340_ divider2.odd_0.counter\[1\] divider2.odd_0.counter\[0\] divider2.odd_0.counter\[2\]
+ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__nor3_1
X_271_ _130_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_469_ clknet_1_0__leaf_divider2.out net42 net30 VGND VGND VPWR VPWR divider2.even_0.N\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_254_ divider2.odd_0.counter\[0\] VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__clkinv_4
X_323_ divider.odd_0.counter\[1\] divider.odd_0.counter\[0\] VGND VGND VPWR VPWR _053_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__240__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__434__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_306_ divider.odd_0.out_counter2 divider.odd_0.out_counter VGND VGND VPWR VPWR _151_
+ sky130_fd_sc_hd__nor2_1
X_237_ _071_ net16 _035_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__222__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__404__S net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input6_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ divider2.even_0.N\[2\] net15 net17 _127_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__o211ai_4
X_468_ clknet_1_1__leaf_divider2.out net43 net30 VGND VGND VPWR VPWR divider2.even_0.N\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_399_ net23 divider2.odd_0.counter\[2\] _128_ _198_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__o31a_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _157_ _158_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2b_1
X_253_ divider2.odd_0.counter2\[0\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__inv_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ divider.odd_0.out_counter2 divider.odd_0.out_counter VGND VGND VPWR VPWR _150_
+ sky130_fd_sc_hd__and2_1
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_236_ _070_ divider2.even_0.N\[2\] net22 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__mux2_1
XFILLER_1_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout27_A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _050_ net18 net24 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__mux2_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_398_ net23 _128_ _022_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__o21bai_1
XANTENNA__446__D net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_467_ clknet_1_0__leaf_divider2.out net7 net30 VGND VGND VPWR VPWR divider2.syncNp\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ divider.odd_0.counter2\[1\] divider.odd_0.counter2\[0\] divider.odd_0.counter2\[2\]
+ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_252_ divider2.odd_0.initial_begin\[0\] VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_net11 clknet_0_net11 VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_16
X_304_ net21 _036_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__nand2b_2
X_235_ _069_ net14 _034_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _049_ net18 _030_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_clk_out_buffer user_clk_buffered VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_397_ net23 divider2.odd_0.counter\[1\] _128_ _197_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__o31a_1
X_466_ clknet_1_1__leaf_divider2.out net6 net30 VGND VGND VPWR VPWR divider2.syncNp\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__433__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__243__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ divider2.even_0.counter\[0\] VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__inv_2
X_320_ divider.odd_0.counter2\[1\] divider.odd_0.counter2\[0\] divider.odd_0.counter2\[2\]
+ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nor3_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_449_ clknet_1_0__leaf_pll_clk90 _105_ net29 VGND VGND VPWR VPWR divider2.even_0.out_counter
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__216__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider.out clknet_0_divider.out VGND VGND VPWR VPWR clknet_1_1__leaf_divider.out
+ sky130_fd_sc_hd__clkbuf_1
X_303_ divider2.odd_0.counter\[1\] divider2.odd_0.counter\[2\] _071_ VGND VGND VPWR
+ VPWR _035_ sky130_fd_sc_hd__nor3_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_234_ _068_ divider2.even_0.N\[1\] net22 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__mux2_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_217_ _048_ net19 net25 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__270__A2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_465_ clknet_1_1__leaf_divider2.out net5 net31 VGND VGND VPWR VPWR divider2.syncNp\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_396_ net23 _128_ _021_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__o21bai_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout20 divider.even_0.N\[0\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_4
X_250_ divider.odd_0.counter\[0\] VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkinv_4
Xfanout31 divider.even_0.resetb VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_448_ clknet_1_0__leaf_pll_clk90 net14 VGND VGND VPWR VPWR divider2.odd_0.old_N\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_379_ divider2.even_0.counter\[0\] _185_ divider2.even_0.out_counter VGND VGND VPWR
+ VPWR _187_ sky130_fd_sc_hd__a21bo_1
X_302_ divider2.odd_0.counter\[1\] divider2.odd_0.counter\[2\] VGND VGND VPWR VPWR
+ _148_ sky130_fd_sc_hd__nor2_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_233_ _067_ divider2.even_0.N\[1\] _034_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__mux2_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_216_ _047_ net19 _030_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_464_ clknet_1_0__leaf_pll_clk90 _120_ net29 VGND VGND VPWR VPWR divider2.even_0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_395_ _071_ _000_ _196_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 divider.even_0.N\[0\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_378_ divider2.even_0.out_counter _185_ divider2.even_0.counter\[0\] VGND VGND VPWR
+ VPWR _186_ sky130_fd_sc_hd__nand3b_1
X_447_ clknet_1_0__leaf_pll_clk90 net15 VGND VGND VPWR VPWR divider2.odd_0.old_N\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_232_ _066_ net17 divider2.odd_0.rst_pulse VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__mux2_1
X_301_ net23 _129_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__nand2b_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__037_ clknet_0__037_ VGND VGND VPWR VPWR clknet_1_0__leaf__037_ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ _046_ net20 net24 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__mux2_1
XANTENNA__429__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_463_ clknet_1_0__leaf_pll_clk90 _119_ net29 VGND VGND VPWR VPWR divider2.even_0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_394_ net23 _128_ _020_ VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__o21ai_1
XANTENNA__237__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_411__6 clknet_1_1__leaf_pll_clk VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__inv_4
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_pll_clk90 clknet_0_pll_clk90 VGND VGND VPWR VPWR clknet_1_1__leaf_pll_clk90
+ sky130_fd_sc_hd__clkbuf_16
X_377_ net16 divider2.even_0.counter\[2\] divider2.even_0.counter\[1\] VGND VGND VPWR
+ VPWR _185_ sky130_fd_sc_hd__nor3_1
X_446_ clknet_1_0__leaf_pll_clk90 net16 VGND VGND VPWR VPWR divider2.odd_0.old_N\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_300_ divider2.even_0.counter\[2\] divider2.even_0.counter\[1\] _077_ VGND VGND VPWR
+ VPWR _032_ sky130_fd_sc_hd__nor3_1
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_231_ _065_ net17 _034_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clknet_0_ext_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_429_ net37 _094_ net28 VGND VGND VPWR VPWR divider.odd_0.out_counter2 sky130_fd_sc_hd__dfstp_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_214_ _045_ net20 _030_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__mux2_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_462_ clknet_1_0__leaf_pll_clk90 _118_ net29 VGND VGND VPWR VPWR divider2.even_0.counter\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_393_ divider2.odd_0.initial_begin\[2\] _025_ _002_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__mux2_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__400__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout23 divider2.odd_0.rst_pulse VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input10_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_445_ clknet_1_1__leaf_pll_clk _104_ VGND VGND VPWR VPWR ext_clk_syncd_pre sky130_fd_sc_hd__dfxtp_1
X_376_ ext_clk_syncd_pre net27 _184_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__o21ba_2
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _063_ _064_ net22 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__mux2_1
X_428_ clknet_1_0__leaf_pll_clk _093_ net28 VGND VGND VPWR VPWR divider.odd_0.counter2\[2\]
+ sky130_fd_sc_hd__dfrtn_1
X_359_ _123_ _142_ _177_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__o21ai_1
Xinput2 ext_reset VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_213_ _043_ _044_ net26 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__mux2_1
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259__4 clknet_1_0__leaf_pll_clk VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__inv_4
X_461_ clknet_1_0__leaf_pll_clk _117_ net28 VGND VGND VPWR VPWR divider.odd_0.out_counter
+ sky130_fd_sc_hd__dfstp_1
X_392_ divider2.odd_0.initial_begin\[0\] _023_ _002_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__mux2_1
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout24 net26 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_444_ clknet_1_1__leaf_divider.out divider.syncNp\[2\] net28 VGND VGND VPWR VPWR
+ divider.even_0.N\[2\] sky130_fd_sc_hd__dfrtp_1
X_375_ net2 clknet_1_0__leaf_ext_clk net4 net3 VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__and4bb_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_358_ net24 _140_ divider.odd_0.counter2\[0\] VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__nand3b_1
X_427_ net36 _092_ net28 VGND VGND VPWR VPWR divider.odd_0.counter2\[1\] sky130_fd_sc_hd__dfstp_2
X_289_ _137_ _138_ net24 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__a21oi_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 porb VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_212_ _041_ _042_ net26 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__mux2_1
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_net11 net11 VGND VGND VPWR VPWR clknet_0_net11 sky130_fd_sc_hd__clkbuf_16
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_460_ clknet_1_0__leaf_pll_clk90 _116_ net29 VGND VGND VPWR VPWR divider2.odd_0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_391_ _126_ _133_ _195_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout25 net26 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout14 divider2.even_0.N\[2\] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
X_443_ clknet_1_0__leaf_divider.out divider.syncNp\[1\] net28 VGND VGND VPWR VPWR
+ divider.even_0.N\[1\] sky130_fd_sc_hd__dfstp_2
X_374_ _182_ _183_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__nand2b_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_426_ clknet_1_0__leaf_pll_clk _091_ net28 VGND VGND VPWR VPWR divider.odd_0.counter2\[0\]
+ sky130_fd_sc_hd__dfrtn_1
X_357_ net26 _138_ _173_ _176_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__o22a_1
X_288_ net18 net19 net20 _030_ _137_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__o2111a_1
Xinput4 resetb VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_211_ _039_ _040_ net26 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__mux2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__285__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_409__9 core_clk VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__inv_4
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_390_ net22 _130_ divider2.odd_0.counter2\[2\] VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__nand3b_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout26 divider.odd_0.rst_pulse VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xfanout15 divider2.even_0.N\[1\] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_pll_clk clknet_0_pll_clk VGND VGND VPWR VPWR clknet_1_1__leaf_pll_clk
+ sky130_fd_sc_hd__clkbuf_16
X_442_ clknet_1_0__leaf_divider.out divider.syncNp\[0\] net29 VGND VGND VPWR VPWR
+ divider.even_0.N\[0\] sky130_fd_sc_hd__dfrtp_1
X_373_ net21 divider.even_0.counter\[1\] divider.even_0.counter\[0\] divider.even_0.counter\[2\]
+ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_287_ _140_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_356_ _174_ _175_ _138_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__o21ai_1
X_425_ clknet_1_0__leaf_pll_clk _090_ net27 VGND VGND VPWR VPWR divider.odd_0.rst_pulse
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 sel2[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ clknet_1_1__leaf__037_ clknet_1_0__leaf_divider2.out use_pll_second VGND VGND
+ VPWR VPWR user_clk_buffered sky130_fd_sc_hd__mux2_1
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_339_ divider2.odd_0.counter\[1\] divider2.odd_0.counter\[0\] VGND VGND VPWR VPWR
+ _073_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_divider2.out clknet_0_divider2.out VGND VGND VPWR VPWR clknet_1_0__leaf_divider2.out
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout16 divider2.even_0.N\[0\] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_4
Xfanout27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_441_ clknet_1_0__leaf_divider.out net10 net29 VGND VGND VPWR VPWR divider.syncNp\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_372_ net21 divider.even_0.counter\[1\] divider.even_0.counter\[0\] divider.even_0.counter\[2\]
+ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__nor4_1
XANTENNA__422__D net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__267__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_424_ clknet_1_1__leaf_pll_clk _089_ net27 VGND VGND VPWR VPWR divider.even_0.out_counter
+ sky130_fd_sc_hd__dfstp_1
X_286_ net18 net19 net20 _137_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__o211ai_4
X_355_ divider.even_0.N\[2\] divider.odd_0.old_N\[2\] VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__and2_1
Xinput6 sel2[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_407_ _201_ _202_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__nand2b_1
X_338_ _163_ _164_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nand2b_1
X_269_ divider2.even_0.N\[2\] divider2.even_0.N\[1\] net17 VGND VGND VPWR VPWR _129_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__406__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__037_ _037_ VGND VGND VPWR VPWR clknet_0__037_ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout17 divider2.even_0.N\[0\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout28 net31 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_440_ clknet_1_0__leaf_divider.out net9 net29 VGND VGND VPWR VPWR divider.syncNp\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_371_ _005_ divider.even_0.counter\[1\] net21 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ divider.even_0.N\[2\] divider.odd_0.old_N\[2\] VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__nor2_1
X_423_ clknet_1_1__leaf_pll_clk net18 VGND VGND VPWR VPWR divider.odd_0.old_N\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__267__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ net18 net19 net20 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__o21ai_2
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel2[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__288__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_406_ net16 divider2.even_0.counter\[1\] divider2.even_0.counter\[0\] divider2.even_0.counter\[2\]
+ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__o31ai_1
X_337_ divider2.odd_0.counter2\[1\] divider2.odd_0.counter2\[0\] divider2.odd_0.counter2\[2\]
+ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__o21ai_1
X_268_ net14 net15 net16 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__o21a_4
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 sel[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_divider.out clknet_0_divider.out VGND VGND VPWR VPWR clknet_1_0__leaf_divider.out
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout29 net30 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
Xfanout18 divider.even_0.N\[2\] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ _004_ divider.even_0.counter\[0\] net21 VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__mux2_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ net18 net19 net20 VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__o21a_1
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__283__B net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_353_ _171_ _172_ divider.odd_0.old_N\[0\] VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__nand3_1
X_422_ clknet_1_1__leaf_pll_clk net19 VGND VGND VPWR VPWR divider.odd_0.old_N\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 sel[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_pll_clk clknet_0_pll_clk VGND VGND VPWR VPWR clknet_1_0__leaf_pll_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__384__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_405_ net16 divider2.even_0.counter\[2\] divider2.even_0.counter\[1\] divider2.even_0.counter\[0\]
+ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__nor4_1
X_267_ net14 net15 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__nor2_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_336_ divider2.odd_0.counter2\[1\] divider2.odd_0.counter2\[0\] divider2.odd_0.counter2\[2\]
+ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nor3_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__381__A_N net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ divider.odd_0.counter2\[1\] divider.odd_0.counter2\[0\] VGND VGND VPWR VPWR
+ _047_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout19 divider.even_0.N\[1\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_4
XANTENNA_input9_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__242__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__447__D net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_412__2 clknet_1_1__leaf_pll_clk90 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__inv_4
X_421_ clknet_1_1__leaf_pll_clk net21 VGND VGND VPWR VPWR divider.odd_0.old_N\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_283_ net18 net19 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
X_352_ divider.odd_0.old_N\[1\] divider.even_0.N\[1\] VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__nand2b_1
Xinput9 sel[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_404_ _016_ divider2.even_0.counter\[1\] net16 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__mux2_1
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ divider2.odd_0.initial_begin\[1\] divider2.odd_0.initial_begin\[2\] VGND VGND
+ VPWR VPWR _127_ sky130_fd_sc_hd__nor2_2
X_335_ divider2.odd_0.counter2\[1\] divider2.odd_0.counter2\[0\] VGND VGND VPWR VPWR
+ _067_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ divider.odd_0.counter2\[0\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_1
XANTENNA__345__B1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_318_ _039_ _137_ _156_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a21o_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 divider2.syncNp\[2\] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_divider2.out divider2.out VGND VGND VPWR VPWR clknet_0_divider2.out sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ divider.even_0.N\[1\] divider.odd_0.old_N\[1\] VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__nand2b_1
X_420_ clknet_1_1__leaf_pll_clk net45 net27 VGND VGND VPWR VPWR ext_clk_syncd sky130_fd_sc_hd__dfrtp_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_282_ divider.odd_0.initial_begin\[1\] divider.odd_0.initial_begin\[2\] VGND VGND
+ VPWR VPWR _137_ sky130_fd_sc_hd__nor2_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__426__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_403_ _015_ divider2.even_0.counter\[0\] net16 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__mux2_1
X_334_ _059_ _127_ _162_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21o_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ divider2.odd_0.counter2\[1\] divider2.odd_0.counter2\[2\] divider2.odd_0.counter2\[0\]
+ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nor3b_4
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__345__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_317_ divider.odd_0.initial_begin\[1\] divider.odd_0.initial_begin\[0\] divider.odd_0.initial_begin\[2\]
+ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__o21a_1
X_248_ divider.odd_0.initial_begin\[0\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__inv_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 divider2.syncNp\[1\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_262__1 clknet_1_1__leaf_pll_clk90 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__inv_4
X_350_ _169_ _170_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand2_1
X_281_ divider.odd_0.counter2\[1\] divider.odd_0.counter2\[2\] divider.odd_0.counter2\[0\]
+ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nor3b_2
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ divider.odd_0.out_counter _199_ _200_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__o21ai_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ divider2.odd_0.initial_begin\[1\] _024_ _002_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__mux2_1
X_333_ divider2.odd_0.initial_begin\[1\] divider2.odd_0.initial_begin\[0\] divider2.odd_0.initial_begin\[2\]
+ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__o21a_1
XFILLER_25_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__345__A2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_316_ _155_ _044_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__nor2_1
X_247_ divider.even_0.counter\[0\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 divider2.syncNp\[0\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input7_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_280_ divider.odd_0.counter2\[1\] divider.odd_0.counter2\[2\] VGND VGND VPWR VPWR
+ _136_ sky130_fd_sc_hd__nor2_1
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_divider2.out clknet_0_divider2.out VGND VGND VPWR VPWR clknet_1_1__leaf_divider2.out
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__435__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_401_ _199_ divider.odd_0.out_counter net24 VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__a21oi_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_332_ _161_ _064_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nor2_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _019_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__inv_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ divider.odd_0.out_counter2 VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__clkinv_4
X_315_ divider.even_0.N\[1\] net20 net18 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__o21a_1
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_229_ _061_ _062_ net22 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__mux2_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 reset_delay\[1\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_400_ net18 net19 net20 divider.odd_0.counter\[0\] _147_ VGND VGND VPWR VPWR _199_
+ sky130_fd_sc_hd__o2111ai_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ divider2.even_0.N\[1\] net17 net14 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__o21a_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_ext_clk clknet_0_ext_clk VGND VGND VPWR VPWR clknet_1_1__leaf_ext_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__414__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ divider.even_0.N\[2\] divider.even_0.N\[1\] net20 VGND VGND VPWR VPWR _155_
+ sky130_fd_sc_hd__nor3_1
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ divider2.odd_0.out_counter2 VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__clkinv_4
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_228_ _059_ _060_ net22 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__mux2_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 ext_clk_syncd_pre VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__444__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_330_ net14 net15 net16 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__nor3_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_261_ _017_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__inv_2
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ clknet_1_0__leaf_pll_clk90 _115_ net29 VGND VGND VPWR VPWR divider2.odd_0.counter\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_23_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_244_ _078_ net14 _032_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__mux2_1
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ divider.odd_0.initial_begin\[1\] divider.odd_0.initial_begin\[0\] VGND VGND
+ VPWR VPWR _041_ sky130_fd_sc_hd__xnor2_1
XANTENNA__330__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_227_ divider.even_0.N\[2\] _058_ _028_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__mux2_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__239__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 use_pll_first VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _008_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__inv_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_458_ clknet_1_0__leaf_pll_clk90 _114_ net30 VGND VGND VPWR VPWR divider2.odd_0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_389_ _125_ _133_ _194_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21ai_1
XANTENNA__284__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__443__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__328__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_243_ _077_ net15 _032_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__mux2_1
X_312_ net19 net20 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__330__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ divider.even_0.N\[1\] _057_ _028_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 reset_delay\[2\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
X_209_ divider2.even_0.out_counter clknet_1_1__leaf_pll_clk90 _027_ VGND VGND VPWR
+ VPWR _038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_457_ clknet_1_1__leaf_pll_clk90 _113_ net30 VGND VGND VPWR VPWR divider2.odd_0.initial_begin\[2\]
+ sky130_fd_sc_hd__dfrtn_1
X_388_ net22 _130_ divider2.odd_0.counter2\[0\] VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__nand3b_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__328__B net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_242_ _076_ net14 net23 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__mux2_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_311_ _154_ _129_ _153_ _152_ VGND VGND VPWR VPWR divider2.out sky130_fd_sc_hd__o31ai_2
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__330__C net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_ext_clk clknet_0_ext_clk VGND VGND VPWR VPWR clknet_1_0__leaf_ext_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_225_ _056_ net18 net25 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__mux2_1
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_208_ clknet_1_0__leaf__037_ clknet_1_1__leaf_divider.out use_pll_second VGND VGND
+ VPWR VPWR net11 sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257__7 clknet_1_1__leaf_net11 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__inv_4
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_456_ net35 _112_ net27 VGND VGND VPWR VPWR divider2.odd_0.initial_begin\[1\] sky130_fd_sc_hd__dfstp_1
X_387_ net23 _128_ _190_ _193_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__o22a_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_310_ divider2.odd_0.out_counter2 divider2.odd_0.out_counter VGND VGND VPWR VPWR
+ _154_ sky130_fd_sc_hd__nor2_1
X_241_ _075_ net14 _035_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__mux2_1
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_439_ clknet_1_0__leaf_divider.out net8 net29 VGND VGND VPWR VPWR divider.syncNp\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_224_ _055_ net18 _031_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__mux2_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_207_ clknet_1_1__leaf_ext_clk ext_clk_syncd use_pll_first VGND VGND VPWR VPWR _037_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ _191_ _192_ _128_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_455_ clknet_1_1__leaf_pll_clk90 _111_ net30 VGND VGND VPWR VPWR divider2.odd_0.initial_begin\[0\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _074_ net15 net23 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__mux2_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_369_ net25 _181_ _001_ _011_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_438_ clknet_1_1__leaf_pll_clk _103_ net27 VGND VGND VPWR VPWR divider.even_0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_223_ _054_ net19 net25 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__mux2_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ divider.even_0.out_counter clknet_1_0__leaf_pll_clk _026_ VGND VGND VPWR VPWR
+ _036_ sky130_fd_sc_hd__mux2_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__403__S net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_385_ net14 divider2.odd_0.old_N\[2\] VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__and2_1
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_454_ net34 _110_ net30 VGND VGND VPWR VPWR divider2.odd_0.out_counter2 sky130_fd_sc_hd__dfstp_1
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ _139_ divider.odd_0.counter\[2\] VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__nand2_1
X_299_ divider.odd_0.counter\[1\] divider.odd_0.counter\[2\] _051_ VGND VGND VPWR
+ VPWR _031_ sky130_fd_sc_hd__nor3_2
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_437_ clknet_1_1__leaf_pll_clk _102_ net27 VGND VGND VPWR VPWR divider.even_0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_222_ _053_ net19 _031_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__mux2_1
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _000_ net22 _033_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__mux2_1
XFILLER_2_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clknet_0_pll_clk90 sky130_fd_sc_hd__clkbuf_16
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__377__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__241__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__223__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__461__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_470_ clknet_1_1__leaf_divider2.out net13 net31 VGND VGND VPWR VPWR divider2.even_0.N\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_453_ clknet_1_1__leaf_pll_clk90 _109_ net30 VGND VGND VPWR VPWR divider2.odd_0.counter2\[2\]
+ sky130_fd_sc_hd__dfrtn_1
X_384_ net14 divider2.odd_0.old_N\[2\] VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__nor2_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__385__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_436_ clknet_1_1__leaf_pll_clk _101_ net27 VGND VGND VPWR VPWR divider.even_0.counter\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ divider.odd_0.counter\[1\] divider.odd_0.counter\[2\] VGND VGND VPWR VPWR _147_
+ sky130_fd_sc_hd__nor2_1
X_367_ net24 _180_ _001_ _010_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ _052_ net20 net24 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__mux2_1
XFILLER_8_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_419_ clknet_1_1__leaf_pll_clk90 _088_ net29 VGND VGND VPWR VPWR divider2.odd_0.out_counter
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__382__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_204_ _001_ net24 _029_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__mux2_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__448__D net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_383_ _188_ _189_ divider2.odd_0.old_N\[0\] VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__nand3_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_452_ net33 _108_ net30 VGND VGND VPWR VPWR divider2.odd_0.counter2\[1\] sky130_fd_sc_hd__dfstp_2
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_366_ _139_ divider.odd_0.counter\[1\] VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__nand2_1
X_435_ clknet_1_0__leaf_pll_clk _100_ net28 VGND VGND VPWR VPWR divider.odd_0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_297_ net25 _139_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nand2b_1
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_220_ _051_ net20 _031_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__mux2_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_349_ net21 _028_ divider.even_0.out_counter VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__o21ai_1
X_418_ clknet_1_1__leaf_pll_clk net46 net31 VGND VGND VPWR VPWR use_pll_second sky130_fd_sc_hd__dfrtp_1
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_net11 clknet_0_net11 VGND VGND VPWR VPWR clknet_1_1__leaf_net11 sky130_fd_sc_hd__clkbuf_16
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_413__3 clknet_1_1__leaf_pll_clk90 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__inv_4
X_416__32 VGND VGND VPWR VPWR _416__32/HI net32 sky130_fd_sc_hd__conb_1
XFILLER_17_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_382_ divider2.odd_0.old_N\[1\] net15 VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__nand2b_1
X_451_ clknet_1_1__leaf_pll_clk90 _107_ net30 VGND VGND VPWR VPWR divider2.odd_0.counter2\[0\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ _051_ _001_ _179_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_434_ clknet_1_0__leaf_pll_clk _099_ net28 VGND VGND VPWR VPWR divider.odd_0.counter\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_296_ divider.even_0.counter\[0\] _146_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nand2_1
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_279_ divider.odd_0.initial_begin\[1\] _013_ _003_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__mux2_1
X_417_ clknet_1_1__leaf_pll_clk pll_clk_sel net27 VGND VGND VPWR VPWR use_pll_first
+ sky130_fd_sc_hd__dfrtp_1
X_348_ net21 divider.even_0.out_counter _146_ divider.even_0.counter\[0\] VGND VGND
+ VPWR VPWR _169_ sky130_fd_sc_hd__nand4bb_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__244__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__235__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__217__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_450_ clknet_1_0__leaf_pll_clk90 _106_ net29 VGND VGND VPWR VPWR divider2.odd_0.rst_pulse
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_381_ net15 divider2.odd_0.old_N\[1\] VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__nand2b_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__427__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_433_ clknet_1_0__leaf_pll_clk _098_ net28 VGND VGND VPWR VPWR divider.odd_0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_364_ net24 _138_ _009_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ divider.even_0.counter\[1\] divider.even_0.counter\[2\] VGND VGND VPWR VPWR
+ _146_ sky130_fd_sc_hd__nor2_1
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_410__5 clknet_1_0__leaf_pll_clk VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__inv_4
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_416_ net41 net32 net31 VGND VGND VPWR VPWR reset_delay\[2\] sky130_fd_sc_hd__dfstp_1
X_347_ divider2.odd_0.out_counter _167_ _168_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__o21ai_1
X_278_ _018_ _134_ _135_ net22 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_380_ _186_ _187_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

