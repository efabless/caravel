* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rst_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
X_05903_ _10163_/Q _05897_/X _09547_/A1 _05899_/X VGND VGND VPWR VPWR _10163_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06883_ _09965_/Q VGND VGND VPWR VPWR _06883_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09671_ _09803_/Q _09802_/Q _09773_/Q VGND VGND VPWR VPWR _09671_/X sky130_fd_sc_hd__mux2_1
X_08622_ _09233_/A _09247_/B _09247_/C _08774_/A VGND VGND VPWR VPWR _08766_/B sky130_fd_sc_hd__or4_4
X_05834_ _10204_/Q _05831_/X _09658_/A1 _05832_/Y VGND VGND VPWR VPWR _10204_/D sky130_fd_sc_hd__a22o_1
X_05765_ _05765_/A VGND VGND VPWR VPWR _05765_/X sky130_fd_sc_hd__clkbuf_2
X_08553_ _09278_/A _08553_/B _08546_/B _08552_/X VGND VGND VPWR VPWR _08553_/X sky130_fd_sc_hd__or4bb_1
XFILLER_82_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08484_ _09029_/A VGND VGND VPWR VPWR _08484_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07504_ _10058_/Q VGND VGND VPWR VPWR _07504_/Y sky130_fd_sc_hd__inv_6
X_05696_ _10285_/Q _05690_/X _09576_/X _05692_/X VGND VGND VPWR VPWR _10285_/D sky130_fd_sc_hd__a22o_1
X_07435_ _07421_/X _07427_/A _09751_/Q _07428_/A VGND VGND VPWR VPWR _09751_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07366_ _07364_/Y _05821_/B _07365_/Y _06304_/B VGND VGND VPWR VPWR _07366_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09105_ _09105_/A _09105_/B VGND VGND VPWR VPWR _09105_/Y sky130_fd_sc_hd__nor2_1
X_07297_ _10124_/Q _05073_/Y input47/X _09679_/S _07296_/X VGND VGND VPWR VPWR _07303_/C
+ sky130_fd_sc_hd__a221o_1
X_06317_ _09954_/Q _06314_/X _09581_/X _06316_/X VGND VGND VPWR VPWR _09954_/D sky130_fd_sc_hd__a22o_1
X_09036_ _09036_/A _09036_/B VGND VGND VPWR VPWR _09036_/X sky130_fd_sc_hd__or2_1
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06248_ _06248_/A VGND VGND VPWR VPWR _09989_/D sky130_fd_sc_hd__inv_2
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06179_ _10003_/Q _10002_/Q VGND VGND VPWR VPWR _08027_/A sky130_fd_sc_hd__or2_1
X_09938_ _10313_/CLK _09938_/D repeater404/X VGND VGND VPWR VPWR _09938_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09869_ _10490_/CLK _09869_/D repeater404/X VGND VGND VPWR VPWR _09869_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_85_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10009_ _10500_/CLK _10009_/D repeater407/X VGND VGND VPWR VPWR _10009_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05550_ _05603_/A _05550_/B VGND VGND VPWR VPWR _05552_/A sky130_fd_sc_hd__or2_2
XFILLER_189_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05481_ _10386_/Q _05475_/X _09536_/A3 _05476_/Y VGND VGND VPWR VPWR _10386_/D sky130_fd_sc_hd__a22o_1
X_07220_ _10247_/Q VGND VGND VPWR VPWR _07220_/Y sky130_fd_sc_hd__clkinv_4
X_07151_ _09879_/Q VGND VGND VPWR VPWR _07151_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_185_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06102_ _10042_/Q _06097_/X _09579_/X _06099_/X VGND VGND VPWR VPWR _10042_/D sky130_fd_sc_hd__a22o_1
X_07082_ _09463_/A _06515_/A _09475_/A _06338_/A _07081_/X VGND VGND VPWR VPWR _07089_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_133_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06033_ _10083_/Q _06026_/A _06683_/B1 _06027_/A VGND VGND VPWR VPWR _10083_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07984_ _07011_/Y _06232_/A _06945_/Y _07519_/A _07983_/X VGND VGND VPWR VPWR _07987_/C
+ sky130_fd_sc_hd__o221a_1
X_09723_ _10289_/Q _09499_/A VGND VGND VPWR VPWR _09723_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06935_ _06935_/A _06935_/B _06931_/X _06934_/X VGND VGND VPWR VPWR _07029_/B sky130_fd_sc_hd__or4bb_2
X_06866_ _06864_/Y _06402_/B _06865_/Y _06503_/B VGND VGND VPWR VPWR _06866_/X sky130_fd_sc_hd__o22a_1
X_09654_ _08350_/X _09812_/Q _09770_/Q VGND VGND VPWR VPWR _09654_/X sky130_fd_sc_hd__mux2_1
X_05817_ _10213_/Q _05810_/A _09660_/A1 _05811_/A VGND VGND VPWR VPWR _10213_/D sky130_fd_sc_hd__a22o_1
X_08605_ _08784_/A _08605_/B VGND VGND VPWR VPWR _08605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09585_ _10309_/Q _09661_/A1 _09699_/S VGND VGND VPWR VPWR _09585_/X sky130_fd_sc_hd__mux2_1
X_06797_ _09900_/Q VGND VGND VPWR VPWR _06797_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05748_ _05748_/A VGND VGND VPWR VPWR _05749_/B sky130_fd_sc_hd__clkbuf_4
X_08536_ _08936_/A VGND VGND VPWR VPWR _09020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05679_ _05679_/A VGND VGND VPWR VPWR _05680_/A sky130_fd_sc_hd__inv_2
X_08467_ _08467_/A _08787_/B VGND VGND VPWR VPWR _08784_/A sky130_fd_sc_hd__or2_1
XFILLER_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08398_ _08505_/A _08472_/B _08398_/C VGND VGND VPWR VPWR _08430_/B sky130_fd_sc_hd__or3_2
X_07418_ _07418_/A _07418_/B _07418_/C _07418_/D VGND VGND VPWR VPWR _07419_/D sky130_fd_sc_hd__and4_1
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07349_ _07349_/A _07349_/B _07349_/C _07349_/D VGND VGND VPWR VPWR _07419_/A sky130_fd_sc_hd__and4_1
XFILLER_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10360_ _10364_/CLK _10360_/D repeater410/X VGND VGND VPWR VPWR _10360_/Q sky130_fd_sc_hd__dfrtp_1
X_10291_ _10296_/CLK _10291_/D repeater402/X VGND VGND VPWR VPWR _10291_/Q sky130_fd_sc_hd__dfrtp_1
X_09019_ _08934_/A _09023_/A _09004_/Y _09017_/X _09018_/X VGND VGND VPWR VPWR _09022_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_163_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10489_ _10490_/CLK _10489_/D repeater404/X VGND VGND VPWR VPWR _10489_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04981_ _04981_/A VGND VGND VPWR VPWR _04982_/A sky130_fd_sc_hd__inv_2
X_06720_ _06718_/Y _05138_/A _06719_/Y _05762_/B VGND VGND VPWR VPWR _06720_/X sky130_fd_sc_hd__o22a_1
X_06651_ _06655_/A VGND VGND VPWR VPWR _06652_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05602_ _10337_/Q _05596_/X _09536_/A3 _05597_/Y VGND VGND VPWR VPWR _10337_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09370_ _09388_/B _09370_/B VGND VGND VPWR VPWR _09371_/B sky130_fd_sc_hd__or2_1
X_06582_ _06582_/A VGND VGND VPWR VPWR _09811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08321_ _06992_/Y _08201_/A _07974_/Y _08202_/A VGND VGND VPWR VPWR _08321_/X sky130_fd_sc_hd__o22a_1
X_05533_ _10376_/Q _05529_/X _09580_/X _05531_/X VGND VGND VPWR VPWR _10376_/D sky130_fd_sc_hd__a22o_1
XFILLER_177_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ _05350_/Y _08205_/X _05260_/Y _08206_/X _08251_/X VGND VGND VPWR VPWR _08255_/C
+ sky130_fd_sc_hd__o221a_1
X_05464_ _05497_/A VGND VGND VPWR VPWR _05465_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ _09943_/Q VGND VGND VPWR VPWR _07203_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08183_ _08183_/A VGND VGND VPWR VPWR _08183_/X sky130_fd_sc_hd__buf_2
X_05395_ _05395_/A _09773_/Q _09770_/Q VGND VGND VPWR VPWR _05397_/A sky130_fd_sc_hd__or3_4
XFILLER_192_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07134_ _10152_/Q VGND VGND VPWR VPWR _07134_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_145_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07065_ _10079_/Q VGND VGND VPWR VPWR _07065_/Y sky130_fd_sc_hd__inv_2
Xoutput231 _09514_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput220 _09494_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput253 _09716_/Z VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_2
X_06016_ _10095_/Q _06012_/X _09580_/X _06014_/X VGND VGND VPWR VPWR _10095_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput242 _09466_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_2
Xoutput264 _09726_/Z VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_2
Xoutput275 _09565_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput286 _07491_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_2
XFILLER_181_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput297 _10431_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_2
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07967_ _06990_/Y _07527_/A _06999_/Y _07629_/A VGND VGND VPWR VPWR _07967_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09706_ _10282_/Q _09465_/A VGND VGND VPWR VPWR _09706_/Z sky130_fd_sc_hd__ebufn_1
X_06918_ _10101_/Q _05070_/Y _10137_/Q _06705_/Y _06917_/X VGND VGND VPWR VPWR _06925_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07898_ _10338_/Q VGND VGND VPWR VPWR _07898_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09637_ _09636_/X _09892_/Q _09776_/Q VGND VGND VPWR VPWR _09637_/X sky130_fd_sc_hd__mux2_1
X_06849_ _10086_/Q _06692_/Y _10448_/Q _06688_/X VGND VGND VPWR VPWR _06849_/X sky130_fd_sc_hd__a22o_1
X_09568_ _07050_/Y input82/X input79/X VGND VGND VPWR VPWR _09568_/X sky130_fd_sc_hd__mux2_8
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08519_ _08620_/A _08520_/B VGND VGND VPWR VPWR _09327_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09499_ _09499_/A VGND VGND VPWR VPWR _09500_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10412_ _04807_/A1 _10412_/D _05417_/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfrtp_2
XFILLER_139_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10343_ _10349_/CLK _10343_/D repeater405/X VGND VGND VPWR VPWR _10343_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10274_ _10406_/CLK _10274_/D _05712_/X VGND VGND VPWR VPWR _10274_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05180_ _10482_/Q VGND VGND VPWR VPWR _05180_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08870_ _09229_/A _08757_/A _08869_/Y VGND VGND VPWR VPWR _08871_/C sky130_fd_sc_hd__o21bai_1
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07821_ _06786_/Y _07816_/X _06784_/Y _07817_/X _07820_/X VGND VGND VPWR VPWR _07832_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07752_ _06894_/Y _07634_/X _06899_/Y _07635_/X VGND VGND VPWR VPWR _07752_/X sky130_fd_sc_hd__o22a_1
X_04964_ _04992_/A _05338_/A VGND VGND VPWR VPWR _05085_/A sky130_fd_sc_hd__or2_2
X_04895_ _10490_/Q _04888_/A _09660_/A1 _04889_/A VGND VGND VPWR VPWR _10490_/D sky130_fd_sc_hd__a22o_1
X_07683_ _07252_/Y _07645_/X _07247_/Y _07533_/B _07682_/X VGND VGND VPWR VPWR _07684_/D
+ sky130_fd_sc_hd__o221a_1
X_06703_ input60/X _05114_/X _10062_/Q _05162_/X _06702_/X VGND VGND VPWR VPWR _06715_/A
+ sky130_fd_sc_hd__a221o_1
X_09422_ _09422_/A VGND VGND VPWR VPWR _09422_/Y sky130_fd_sc_hd__inv_2
X_06634_ _09797_/Q _06633_/X _09536_/A3 _05124_/A _09678_/X VGND VGND VPWR VPWR _09797_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09353_ _09353_/A _09353_/B _09353_/C _09049_/Y VGND VGND VPWR VPWR _09431_/C sky130_fd_sc_hd__or4b_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08304_ _07122_/Y _08199_/A _07098_/Y _08200_/A _08303_/X VGND VGND VPWR VPWR _08309_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06565_ _06565_/A _09680_/X VGND VGND VPWR VPWR _06575_/S sky130_fd_sc_hd__or2b_1
XFILLER_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05516_ _09686_/X _10380_/Q _05525_/S VGND VGND VPWR VPWR _05517_/A sky130_fd_sc_hd__mux2_1
X_06496_ _06496_/A VGND VGND VPWR VPWR _06496_/Y sky130_fd_sc_hd__inv_2
X_09284_ _09353_/B _09431_/A _09284_/C _09389_/C VGND VGND VPWR VPWR _09288_/A sky130_fd_sc_hd__or4_2
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08235_ _06729_/Y _08213_/X _06709_/Y _08214_/X VGND VGND VPWR VPWR _08235_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05447_ _05447_/A VGND VGND VPWR VPWR _05447_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08166_ _06882_/Y _08080_/X _06871_/Y _08081_/X _08165_/X VGND VGND VPWR VPWR _08171_/B
+ sky130_fd_sc_hd__o221a_1
X_05378_ _05378_/A VGND VGND VPWR VPWR _05379_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_180_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07117_ _10144_/Q VGND VGND VPWR VPWR _09495_/A sky130_fd_sc_hd__inv_6
XFILLER_146_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08097_ _07357_/Y _08092_/X _07663_/A _08093_/X _08096_/X VGND VGND VPWR VPWR _08098_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07048_ _10410_/Q VGND VGND VPWR VPWR _07048_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08999_ _08999_/A _08999_/B VGND VGND VPWR VPWR _09000_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10326_ _10483_/CLK _10326_/D _05034_/A VGND VGND VPWR VPWR _10326_/Q sky130_fd_sc_hd__dfrtp_4
X_10257_ _10257_/CLK _10257_/D repeater407/X VGND VGND VPWR VPWR _10257_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10188_ _10364_/CLK _10188_/D repeater410/X VGND VGND VPWR VPWR _10188_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06350_ _09933_/Q _06341_/A _09659_/A1 _06342_/A VGND VGND VPWR VPWR _09933_/D sky130_fd_sc_hd__a22o_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06281_ _06282_/A VGND VGND VPWR VPWR _06281_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05301_ _05291_/Y _05952_/B _05294_/Y _05838_/A _05300_/X VGND VGND VPWR VPWR _05321_/B
+ sky130_fd_sc_hd__o221a_1
X_05232_ _09955_/Q VGND VGND VPWR VPWR _05232_/Y sky130_fd_sc_hd__inv_2
X_08020_ _08027_/A _08045_/C _08040_/C VGND VGND VPWR VPWR _08188_/A sky130_fd_sc_hd__or3_4
XFILLER_190_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05163_ _05357_/A _05163_/B VGND VGND VPWR VPWR _06704_/A sky130_fd_sc_hd__nor2_2
X_09971_ _10283_/CLK _09971_/D repeater406/X VGND VGND VPWR VPWR _09971_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05094_ _05980_/B VGND VGND VPWR VPWR _05094_/Y sky130_fd_sc_hd__clkinv_2
X_08922_ _09307_/B _08922_/B _09283_/B _09207_/B VGND VGND VPWR VPWR _08926_/A sky130_fd_sc_hd__or4_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08853_ _08855_/A _08853_/B VGND VGND VPWR VPWR _09357_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05996_ _10106_/Q _05994_/X _09578_/X _05995_/Y VGND VGND VPWR VPWR _10106_/D sky130_fd_sc_hd__a22o_1
X_08784_ _08784_/A VGND VGND VPWR VPWR _08996_/A sky130_fd_sc_hd__inv_2
X_07804_ _07798_/Y _07799_/X _07800_/Y _07801_/X _07803_/X VGND VGND VPWR VPWR _07810_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04947_ _04948_/B VGND VGND VPWR VPWR _04947_/Y sky130_fd_sc_hd__inv_2
X_07735_ _10111_/Q VGND VGND VPWR VPWR _07735_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04878_ _10496_/Q _04872_/X _09536_/A3 _04873_/Y VGND VGND VPWR VPWR _10496_/D sky130_fd_sc_hd__a22o_1
X_09405_ _09405_/A _09405_/B _09405_/C _08596_/A VGND VGND VPWR VPWR _09408_/B sky130_fd_sc_hd__or4b_1
X_07666_ _07827_/A VGND VGND VPWR VPWR _07666_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07597_ _09989_/Q _09988_/Q _07597_/C _07602_/D VGND VGND VPWR VPWR _07812_/A sky130_fd_sc_hd__or4_4
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06617_ _06668_/A VGND VGND VPWR VPWR _06666_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09336_ _09344_/A _09336_/B VGND VGND VPWR VPWR _09336_/X sky130_fd_sc_hd__and2_1
X_06548_ _09821_/Q _06540_/A _09661_/A1 _06541_/A VGND VGND VPWR VPWR _09821_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09267_ _09313_/D VGND VGND VPWR VPWR _09267_/Y sky130_fd_sc_hd__inv_2
X_06479_ _09862_/Q _06473_/X _09574_/X _06474_/Y VGND VGND VPWR VPWR _09862_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08218_ _08218_/A _08218_/B _08218_/C _08218_/D VGND VGND VPWR VPWR _08218_/Y sky130_fd_sc_hd__nand4_4
XFILLER_181_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09198_ _09446_/A _09198_/B _09198_/C VGND VGND VPWR VPWR _09309_/D sky130_fd_sc_hd__or3_1
XFILLER_181_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_134_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08149_ _06973_/Y _08086_/X _06948_/Y _08087_/X _08148_/X VGND VGND VPWR VPWR _08152_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10111_ _10135_/CLK _10111_/D repeater405/X VGND VGND VPWR VPWR _10111_/Q sky130_fd_sc_hd__dfrtp_2
X_10042_ _10404_/CLK _10042_/D repeater410/X VGND VGND VPWR VPWR _10042_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__buf_12
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold30 hold30/A VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 _05261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10309_ _10310_/CLK _10309_/D repeater404/X VGND VGND VPWR VPWR _10309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05850_ _10193_/Q _05841_/A _09574_/X _05842_/A VGND VGND VPWR VPWR _10193_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05781_ _10233_/Q _05776_/X _09661_/A1 _05777_/Y VGND VGND VPWR VPWR _10233_/D sky130_fd_sc_hd__a22o_1
X_07520_ _07546_/C _07597_/C VGND VGND VPWR VPWR _07596_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10257_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07451_ _07452_/A VGND VGND VPWR VPWR _07451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06402_ _06481_/A _06402_/B VGND VGND VPWR VPWR _06404_/A sky130_fd_sc_hd__or2_2
X_07382_ _10366_/Q VGND VGND VPWR VPWR _07382_/Y sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06333_ _09944_/Q _06330_/X _09577_/X _06331_/Y VGND VGND VPWR VPWR _09944_/D sky130_fd_sc_hd__a22o_1
X_09121_ _09326_/B _09287_/A VGND VGND VPWR VPWR _09339_/C sky130_fd_sc_hd__or2_1
XFILLER_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09052_ _09052_/A _09052_/B _08891_/X VGND VGND VPWR VPWR _09056_/C sky130_fd_sc_hd__or3b_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06264_ _06264_/A VGND VGND VPWR VPWR _06264_/Y sky130_fd_sc_hd__inv_2
X_05215_ _05286_/A _05357_/B VGND VGND VPWR VPWR _06515_/A sky130_fd_sc_hd__or2_4
X_06195_ _08000_/B _06193_/Y _09777_/Q _06194_/X VGND VGND VPWR VPWR _10004_/D sky130_fd_sc_hd__a31o_1
X_08003_ _08010_/C _08019_/B _10006_/Q VGND VGND VPWR VPWR _08174_/A sky130_fd_sc_hd__or3_4
X_05146_ _06679_/C VGND VGND VPWR VPWR _05146_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05077_ _10097_/Q _05070_/Y _10123_/Q _05073_/Y _05076_/X VGND VGND VPWR VPWR _05108_/A
+ sky130_fd_sc_hd__a221o_1
X_09954_ _10062_/CLK _09954_/D repeater405/X VGND VGND VPWR VPWR _09954_/Q sky130_fd_sc_hd__dfrtp_1
X_08905_ _08965_/A _08905_/B VGND VGND VPWR VPWR _08933_/A sky130_fd_sc_hd__or2_2
XFILLER_106_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09885_ _09919_/CLK _09885_/D repeater409/X VGND VGND VPWR VPWR _09885_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08836_/A _08836_/B VGND VGND VPWR VPWR _09287_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05979_ _10115_/Q _05970_/A _09574_/X _05971_/A VGND VGND VPWR VPWR _10115_/D sky130_fd_sc_hd__a22o_1
X_08767_ _08767_/A _09384_/B VGND VGND VPWR VPWR _08772_/A sky130_fd_sc_hd__nor2_1
Xrepeater394 _09577_/X VGND VGND VPWR VPWR _09658_/A1 sky130_fd_sc_hd__buf_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08698_ _08701_/A _09048_/A _08697_/X VGND VGND VPWR VPWR _08700_/C sky130_fd_sc_hd__o21ai_1
X_07718_ _10085_/Q VGND VGND VPWR VPWR _07718_/Y sky130_fd_sc_hd__inv_2
X_07649_ _07381_/Y _07645_/X _07406_/Y _07533_/B _07648_/X VGND VGND VPWR VPWR _07650_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09319_ _09319_/A _09319_/B _09319_/C _08577_/X VGND VGND VPWR VPWR _09447_/A sky130_fd_sc_hd__or4b_1
XFILLER_178_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput120 sram_ro_data[5] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__buf_2
Xinput153 wb_adr_i[29] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_adr_i[19] VGND VGND VPWR VPWR _08399_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 usr2_vdd_pwrgood VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__buf_6
X_10025_ _10411_/CLK _10025_/D repeater407/X VGND VGND VPWR VPWR _10025_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput164 wb_cyc_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput186 wb_dat_i[29] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[19] VGND VGND VPWR VPWR _08363_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput197 wb_rst_i VGND VGND VPWR VPWR _07450_/A sky130_fd_sc_hd__buf_8
XFILLER_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05000_ _10447_/Q _04994_/X _09545_/A1 _04996_/X VGND VGND VPWR VPWR _10447_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06951_ _10390_/Q VGND VGND VPWR VPWR _06951_/Y sky130_fd_sc_hd__clkinv_2
X_05902_ _10164_/Q _05897_/X _09579_/X _05899_/X VGND VGND VPWR VPWR _10164_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _09669_/X _10394_/Q _10299_/Q VGND VGND VPWR VPWR _09670_/X sky130_fd_sc_hd__mux2_4
X_08621_ _09102_/D _09223_/B _08621_/C VGND VGND VPWR VPWR _08882_/A sky130_fd_sc_hd__or3_1
X_06882_ _09873_/Q VGND VGND VPWR VPWR _06882_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05833_ _10205_/Q _05831_/X _09545_/A1 _05832_/Y VGND VGND VPWR VPWR _10205_/D sky130_fd_sc_hd__a22o_1
X_05764_ _05764_/A VGND VGND VPWR VPWR _05765_/A sky130_fd_sc_hd__inv_2
X_08552_ _08552_/A _08552_/B VGND VGND VPWR VPWR _08552_/X sky130_fd_sc_hd__or2_1
X_08483_ _08571_/C _09236_/A _09295_/A _08483_/D VGND VGND VPWR VPWR _09029_/A sky130_fd_sc_hd__or4_4
X_07503_ _10032_/Q VGND VGND VPWR VPWR _07503_/Y sky130_fd_sc_hd__inv_6
X_05695_ _10286_/Q _05690_/X _09550_/A0 _05692_/X VGND VGND VPWR VPWR _10286_/D sky130_fd_sc_hd__a22o_1
X_07434_ _07290_/X _07427_/A _09752_/Q _07428_/A VGND VGND VPWR VPWR _09752_/D sky130_fd_sc_hd__o22a_1
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07365_ _09956_/Q VGND VGND VPWR VPWR _07365_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09104_ _09104_/A VGND VGND VPWR VPWR _09104_/Y sky130_fd_sc_hd__inv_2
X_07296_ input62/X _06844_/X input12/X _06698_/X VGND VGND VPWR VPWR _07296_/X sky130_fd_sc_hd__a22o_1
X_06316_ _06316_/A VGND VGND VPWR VPWR _06316_/X sky130_fd_sc_hd__clkbuf_2
X_09035_ _09082_/A _09035_/B VGND VGND VPWR VPWR _09036_/B sky130_fd_sc_hd__or2_1
XFILLER_108_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06247_ _09777_/Q _07611_/A _07612_/A _06243_/A _06203_/Y VGND VGND VPWR VPWR _06248_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06178_ _06227_/B VGND VGND VPWR VPWR _06184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05129_ _05129_/A VGND VGND VPWR VPWR _05129_/X sky130_fd_sc_hd__buf_2
X_09937_ _10310_/CLK _09937_/D repeater404/X VGND VGND VPWR VPWR _09937_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09868_ _10490_/CLK _09868_/D repeater404/X VGND VGND VPWR VPWR _09868_/Q sky130_fd_sc_hd__dfstp_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _08836_/A _08819_/B VGND VGND VPWR VPWR _09283_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09799_ _10406_/CLK _09799_/D _06628_/X VGND VGND VPWR VPWR _09799_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10008_ _10411_/CLK _10008_/D repeater407/X VGND VGND VPWR VPWR _10008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05480_ _10387_/Q _05475_/X _06684_/B1 _05476_/Y VGND VGND VPWR VPWR _10387_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07150_ _10256_/Q VGND VGND VPWR VPWR _07150_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07081_ _09497_/A _05882_/A _07080_/Y _06079_/B VGND VGND VPWR VPWR _07081_/X sky130_fd_sc_hd__o22a_1
X_06101_ _10043_/Q _06097_/X _09580_/X _06099_/X VGND VGND VPWR VPWR _10043_/D sky130_fd_sc_hd__a22o_1
X_06032_ _10084_/Q _06025_/X _09658_/A1 _06027_/X VGND VGND VPWR VPWR _10084_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_24_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10313_/CLK sky130_fd_sc_hd__clkbuf_16
X_09722_ _10508_/Q _09497_/A VGND VGND VPWR VPWR _09722_/Z sky130_fd_sc_hd__ebufn_1
X_07983_ _07983_/A _07983_/B VGND VGND VPWR VPWR _07983_/X sky130_fd_sc_hd__or2_1
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_39_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10371_/CLK sky130_fd_sc_hd__clkbuf_16
X_06934_ _06932_/Y _06291_/B _05139_/X _06780_/X _06933_/Y VGND VGND VPWR VPWR _06934_/X
+ sky130_fd_sc_hd__o2111a_1
X_06865_ _09846_/Q VGND VGND VPWR VPWR _06865_/Y sky130_fd_sc_hd__clkinv_2
X_09653_ _08348_/Y input58/X _09770_/Q VGND VGND VPWR VPWR _09653_/X sky130_fd_sc_hd__mux2_1
X_09584_ _09581_/X _10307_/Q _09677_/S VGND VGND VPWR VPWR _09584_/X sky130_fd_sc_hd__mux2_1
X_05816_ _10214_/Q _05809_/X _09550_/A0 _05811_/X VGND VGND VPWR VPWR _10214_/D sky130_fd_sc_hd__a22o_1
X_08604_ _08385_/B _08491_/C _08980_/B _09415_/A _08603_/X VGND VGND VPWR VPWR _08605_/B
+ sky130_fd_sc_hd__a311oi_1
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08535_ _08585_/A _08581_/B VGND VGND VPWR VPWR _09446_/A sky130_fd_sc_hd__nor2_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06796_ _09953_/Q VGND VGND VPWR VPWR _06796_/Y sky130_fd_sc_hd__inv_2
X_05747_ _10253_/Q _05741_/X _09574_/X _05742_/Y VGND VGND VPWR VPWR _10253_/D sky130_fd_sc_hd__a22o_1
X_05678_ _05679_/A VGND VGND VPWR VPWR _05678_/X sky130_fd_sc_hd__clkbuf_2
X_08466_ _08466_/A VGND VGND VPWR VPWR _08787_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08397_ _08493_/B VGND VGND VPWR VPWR _08398_/C sky130_fd_sc_hd__inv_2
X_07417_ _07412_/Y _05527_/A _07413_/Y _06480_/A _07416_/X VGND VGND VPWR VPWR _07418_/D
+ sky130_fd_sc_hd__o221a_1
X_07348_ _07343_/Y _06635_/B _07344_/Y _06010_/A _07347_/X VGND VGND VPWR VPWR _07349_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07279_ _07277_/Y _06037_/B _07278_/Y _06494_/B VGND VGND VPWR VPWR _07279_/X sky130_fd_sc_hd__o22a_1
X_10290_ _10290_/CLK _10290_/D repeater402/X VGND VGND VPWR VPWR _10290_/Q sky130_fd_sc_hd__dfrtp_1
X_09018_ _09020_/A _08961_/B _09162_/A VGND VGND VPWR VPWR _09018_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10488_ _10495_/CLK _10488_/D repeater404/X VGND VGND VPWR VPWR _10488_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04980_ _04981_/A VGND VGND VPWR VPWR _04980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06650_ _06650_/A VGND VGND VPWR VPWR _06650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05601_ _10338_/Q _05596_/X _06684_/B1 _05597_/Y VGND VGND VPWR VPWR _10338_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06581_ input58/X _09811_/Q _06581_/S VGND VGND VPWR VPWR _06582_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08320_ _07004_/Y _08193_/A _06938_/Y _08194_/A _08319_/X VGND VGND VPWR VPWR _08327_/A
+ sky130_fd_sc_hd__o221a_1
X_05532_ _10377_/Q _05529_/X _09581_/X _05531_/X VGND VGND VPWR VPWR _10377_/D sky130_fd_sc_hd__a22o_1
XFILLER_177_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05463_ _06663_/A VGND VGND VPWR VPWR _05497_/A sky130_fd_sc_hd__buf_2
X_08251_ _05204_/Y _08207_/X _05312_/Y _08208_/X VGND VGND VPWR VPWR _08251_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07202_ _10372_/Q VGND VGND VPWR VPWR _07202_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05394_ _05394_/A VGND VGND VPWR VPWR _05394_/X sky130_fd_sc_hd__clkbuf_1
X_08182_ _06829_/Y _08177_/X _06783_/Y _08178_/X _08181_/X VGND VGND VPWR VPWR _08218_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_145_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07133_ _10040_/Q VGND VGND VPWR VPWR _09487_/A sky130_fd_sc_hd__clkinv_8
XFILLER_173_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput210 _09476_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07064_ _07048_/Y _05419_/B _07051_/X _07057_/X _07063_/X VGND VGND VPWR VPWR _07064_/X
+ sky130_fd_sc_hd__o2111a_1
Xoutput232 _09516_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput221 _09496_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_06015_ _10096_/Q _06012_/X _09581_/X _06014_/X VGND VGND VPWR VPWR _10096_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput243 _09468_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_2
Xoutput265 _09727_/Z VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput254 _09717_/Z VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput276 _09702_/Z VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput298 _10432_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_2
Xoutput287 _09573_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_2
X_07966_ _06928_/Y _07777_/A _06938_/Y _07778_/A _07965_/X VGND VGND VPWR VPWR _07988_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09705_ _09705_/A _09463_/A VGND VGND VPWR VPWR _09705_/Z sky130_fd_sc_hd__ebufn_1
X_06917_ input56/X _05114_/A input16/X _06698_/A VGND VGND VPWR VPWR _06917_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07897_ _07895_/Y _07799_/X _07320_/Y _07801_/X _07896_/X VGND VGND VPWR VPWR _07901_/C
+ sky130_fd_sc_hd__o221a_1
X_09636_ _07988_/Y _10328_/Q _09682_/S VGND VGND VPWR VPWR _09636_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06848_ input68/X _09679_/S _10334_/Q _05151_/X _06847_/X VGND VGND VPWR VPWR _06855_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06779_ _10113_/Q VGND VGND VPWR VPWR _06779_/Y sky130_fd_sc_hd__inv_2
X_09567_ _09780_/Q _07049_/Y hold1/A VGND VGND VPWR VPWR _09567_/X sky130_fd_sc_hd__mux2_4
X_09498_ _09498_/A VGND VGND VPWR VPWR _09498_/X sky130_fd_sc_hd__clkbuf_1
X_08518_ _08746_/A _08520_/B VGND VGND VPWR VPWR _09030_/A sky130_fd_sc_hd__or2_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08449_ _09085_/C _08631_/B _09085_/B VGND VGND VPWR VPWR _09344_/A sky130_fd_sc_hd__or3_4
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10411_ _10411_/CLK _10411_/D repeater407/X VGND VGND VPWR VPWR _10411_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10342_ _09572_/A1 _10342_/D _05589_/X VGND VGND VPWR VPWR _10342_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10273_ _10504_/CLK _10273_/D repeater403/X VGND VGND VPWR VPWR _10273_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07820_ _06828_/Y _07818_/X _06779_/Y _07819_/X VGND VGND VPWR VPWR _07820_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07751_ _06882_/Y _07627_/X _06877_/Y _07628_/X _07750_/X VGND VGND VPWR VPWR _07761_/A
+ sky130_fd_sc_hd__o221a_1
X_06702_ input99/X _05101_/X input117/X _05112_/A VGND VGND VPWR VPWR _06702_/X sky130_fd_sc_hd__a22o_2
X_04963_ _05005_/C _04963_/B _05027_/A _04991_/B VGND VGND VPWR VPWR _05338_/A sky130_fd_sc_hd__or4_2
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_04894_ _10491_/Q _04887_/X _09550_/A0 _04889_/X VGND VGND VPWR VPWR _10491_/D sky130_fd_sc_hd__a22o_1
X_07682_ _07207_/Y _07646_/X _07208_/Y _07647_/X VGND VGND VPWR VPWR _07682_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _09421_/A _09421_/B _09421_/C _09421_/D VGND VGND VPWR VPWR _09450_/A sky130_fd_sc_hd__or4_1
X_06633_ _06633_/A VGND VGND VPWR VPWR _06633_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09352_ _09352_/A _09352_/B _09352_/C VGND VGND VPWR VPWR _09353_/C sky130_fd_sc_hd__nor3_1
X_06564_ _07489_/A _06601_/B _05397_/A _06579_/D _06563_/X VGND VGND VPWR VPWR _06565_/A
+ sky130_fd_sc_hd__o32a_1
X_05515_ _05515_/A VGND VGND VPWR VPWR _05515_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08303_ _07146_/Y _08201_/A _07948_/Y _08202_/A VGND VGND VPWR VPWR _08303_/X sky130_fd_sc_hd__o22a_1
X_06495_ _06496_/A VGND VGND VPWR VPWR _06495_/X sky130_fd_sc_hd__clkbuf_2
X_09283_ _09283_/A _09283_/B _09283_/C VGND VGND VPWR VPWR _09389_/C sky130_fd_sc_hd__or3_1
X_08234_ _06710_/Y _08205_/X _06753_/Y _08206_/X _08233_/X VGND VGND VPWR VPWR _08237_/C
+ sky130_fd_sc_hd__o221a_1
X_05446_ _05459_/A VGND VGND VPWR VPWR _05447_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08165_ _06895_/Y _08082_/X _06874_/Y _08083_/X VGND VGND VPWR VPWR _08165_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05377_ _10421_/Q _09810_/Q _09772_/Q _05376_/X VGND VGND VPWR VPWR _10421_/D sky130_fd_sc_hd__o211a_1
X_07116_ _10118_/Q VGND VGND VPWR VPWR _09493_/A sky130_fd_sc_hd__clkinv_4
XFILLER_180_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08096_ _07346_/Y _08094_/X _07363_/Y _08095_/X VGND VGND VPWR VPWR _08096_/X sky130_fd_sc_hd__o22a_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07047_ _07047_/A _07047_/B _07047_/C VGND VGND VPWR VPWR _07158_/B sky130_fd_sc_hd__or3_2
XFILLER_133_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08998_ _08998_/A VGND VGND VPWR VPWR _09312_/A sky130_fd_sc_hd__inv_2
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07949_ _07121_/Y _07646_/A _07153_/Y _07807_/A VGND VGND VPWR VPWR _07949_/X sky130_fd_sc_hd__o22a_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09619_ _09618_/X _09883_/Q _09776_/Q VGND VGND VPWR VPWR _09619_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10325_ _10510_/CLK _10325_/D _05034_/A VGND VGND VPWR VPWR _10325_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10256_ _10411_/CLK _10256_/D repeater407/X VGND VGND VPWR VPWR _10256_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ _10191_/CLK _10187_/D repeater410/X VGND VGND VPWR VPWR _10187_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06280_ _06304_/A _06280_/B VGND VGND VPWR VPWR _06282_/A sky130_fd_sc_hd__or2_2
X_05300_ _05296_/Y _05992_/A _05298_/Y _05820_/A VGND VGND VPWR VPWR _05300_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05231_ _05346_/A _05349_/B VGND VGND VPWR VPWR _06279_/A sky130_fd_sc_hd__or2_1
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05162_ _05162_/A VGND VGND VPWR VPWR _05162_/X sky130_fd_sc_hd__clkbuf_2
X_09970_ _10283_/CLK _09970_/D repeater406/X VGND VGND VPWR VPWR _09970_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05093_ _06630_/A _05198_/A VGND VGND VPWR VPWR _05980_/B sky130_fd_sc_hd__or2_2
XFILLER_170_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08921_ _08927_/A _08921_/B _08921_/C VGND VGND VPWR VPWR _09207_/B sky130_fd_sc_hd__nor3_1
XFILLER_130_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08852_ _08852_/A _09342_/B VGND VGND VPWR VPWR _08854_/A sky130_fd_sc_hd__or2_1
X_07803_ _06824_/Y _07755_/X _06802_/Y _07802_/X VGND VGND VPWR VPWR _07803_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05995_ _05995_/A VGND VGND VPWR VPWR _05995_/Y sky130_fd_sc_hd__inv_2
X_08783_ _08783_/A _08783_/B VGND VGND VPWR VPWR _09139_/A sky130_fd_sc_hd__nor2_1
X_07734_ _06973_/Y _07533_/D _07021_/Y _07651_/X _07733_/X VGND VGND VPWR VPWR _07743_/A
+ sky130_fd_sc_hd__o221a_1
X_04946_ _05118_/A _05173_/B VGND VGND VPWR VPWR _04948_/B sky130_fd_sc_hd__or2_1
X_07665_ _07825_/A VGND VGND VPWR VPWR _07665_/X sky130_fd_sc_hd__clkbuf_2
X_09404_ _09383_/Y _09385_/X _09392_/Y _09394_/X _09403_/Y VGND VGND VPWR VPWR _09404_/Y
+ sky130_fd_sc_hd__o221ai_1
X_04877_ _10497_/Q _04872_/X _06684_/B1 _04873_/Y VGND VGND VPWR VPWR _10497_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06616_ _09803_/Q _06604_/X _09648_/X _06606_/X VGND VGND VPWR VPWR _09803_/D sky130_fd_sc_hd__a22o_1
X_07596_ _07601_/A _07596_/B VGND VGND VPWR VPWR _07811_/A sky130_fd_sc_hd__or2_4
X_09335_ _08788_/A _09334_/X _09257_/X VGND VGND VPWR VPWR _09422_/A sky130_fd_sc_hd__o21ai_1
X_06547_ _09822_/Q _06540_/A _09660_/A1 _06541_/A VGND VGND VPWR VPWR _09822_/D sky130_fd_sc_hd__a22o_1
X_06478_ _09863_/Q _06473_/X hold46/X _06474_/Y VGND VGND VPWR VPWR _09863_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09266_ _08812_/A _09105_/B _08860_/A _09099_/X _08863_/A VGND VGND VPWR VPWR _09343_/B
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08217_ _08217_/A _08217_/B _08217_/C _08217_/D VGND VGND VPWR VPWR _08218_/D sky130_fd_sc_hd__and4_2
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05429_ _05429_/A _06579_/D _06593_/A _05429_/D VGND VGND VPWR VPWR _05430_/A sky130_fd_sc_hd__or4_2
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09197_ _09432_/A _09425_/A _09415_/A VGND VGND VPWR VPWR _09315_/A sky130_fd_sc_hd__or3_1
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08148_ _06976_/Y _08088_/X _06943_/Y _08089_/X VGND VGND VPWR VPWR _08148_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08079_ _07325_/Y _08074_/X _07395_/Y _08075_/X _08078_/X VGND VGND VPWR VPWR _08098_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10110_ _10110_/CLK _10110_/D repeater405/X VGND VGND VPWR VPWR _10110_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10041_ _10404_/CLK _10041_/D repeater410/X VGND VGND VPWR VPWR _10041_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 hold20/A VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 porb VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _05261_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10308_ _10313_/CLK _10308_/D repeater404/X VGND VGND VPWR VPWR _10308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10239_ _10491_/CLK _10239_/D repeater403/X VGND VGND VPWR VPWR _10239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05780_ _10234_/Q _05776_/X _09576_/X _05777_/Y VGND VGND VPWR VPWR _10234_/D sky130_fd_sc_hd__a22o_1
X_07450_ _07450_/A _07450_/B VGND VGND VPWR VPWR _07452_/A sky130_fd_sc_hd__or2_2
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07381_ _09895_/Q VGND VGND VPWR VPWR _07381_/Y sky130_fd_sc_hd__inv_2
X_06401_ _06401_/A VGND VGND VPWR VPWR _06402_/B sky130_fd_sc_hd__buf_2
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06332_ _09945_/Q _06330_/X _09545_/A1 _06331_/Y VGND VGND VPWR VPWR _09945_/D sky130_fd_sc_hd__a22o_1
X_09120_ _09260_/A _09109_/B _09117_/X _09119_/Y VGND VGND VPWR VPWR _09120_/X sky130_fd_sc_hd__o211a_1
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09051_ _09051_/A _09051_/B VGND VGND VPWR VPWR _09083_/B sky130_fd_sc_hd__or2_1
XFILLER_190_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06263_ _07477_/A _06133_/Y _06203_/Y _06262_/X VGND VGND VPWR VPWR _06264_/A sky130_fd_sc_hd__a31o_1
X_08002_ _08026_/A _10002_/Q _08032_/B _08019_/C VGND VGND VPWR VPWR _08173_/A sky130_fd_sc_hd__or4_4
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05214_ _05277_/A VGND VGND VPWR VPWR _05357_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06194_ _06184_/A _07989_/B _06177_/A _10004_/Q VGND VGND VPWR VPWR _06194_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05145_ _05167_/A _05148_/A VGND VGND VPWR VPWR _06679_/C sky130_fd_sc_hd__or2_1
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05076_ _10511_/Q _04835_/Y input71/X _06770_/A VGND VGND VPWR VPWR _05076_/X sky130_fd_sc_hd__a22o_1
X_09953_ _10191_/CLK _09953_/D repeater405/X VGND VGND VPWR VPWR _09953_/Q sky130_fd_sc_hd__dfrtp_1
X_08904_ _08921_/B _08943_/A VGND VGND VPWR VPWR _09307_/C sky130_fd_sc_hd__nor2_2
XFILLER_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09884_ _10023_/CLK _09884_/D repeater409/X VGND VGND VPWR VPWR _09884_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08835_ _08835_/A _08847_/B VGND VGND VPWR VPWR _09068_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08766_/A _08766_/B VGND VGND VPWR VPWR _09384_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05978_ _10116_/Q _05970_/A hold46/X _05971_/A VGND VGND VPWR VPWR _10116_/D sky130_fd_sc_hd__a22o_1
Xrepeater395 _09577_/X VGND VGND VPWR VPWR _09550_/A0 sky130_fd_sc_hd__buf_12
XFILLER_122_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07717_ _07717_/A _07717_/B _07717_/C VGND VGND VPWR VPWR _07717_/Y sky130_fd_sc_hd__nand3_2
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08697_ _08697_/A _08697_/B VGND VGND VPWR VPWR _08697_/X sky130_fd_sc_hd__or2_1
X_04929_ _04929_/A VGND VGND VPWR VPWR _10480_/D sky130_fd_sc_hd__clkbuf_1
X_07648_ _07407_/Y _07646_/X _07338_/Y _07647_/X VGND VGND VPWR VPWR _07648_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07579_ _07579_/A VGND VGND VPWR VPWR _07788_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09318_ _09384_/B _09318_/B VGND VGND VPWR VPWR _09417_/B sky130_fd_sc_hd__or2_1
XFILLER_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09249_ _09249_/A _09416_/B VGND VGND VPWR VPWR _09331_/D sky130_fd_sc_hd__or2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 sram_ro_data[25] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__buf_2
Xinput143 wb_adr_i[1] VGND VGND VPWR VPWR _09102_/C sky130_fd_sc_hd__clkbuf_4
Xinput132 wb_adr_i[0] VGND VGND VPWR VPWR _08494_/A sky130_fd_sc_hd__clkbuf_4
Xinput154 wb_adr_i[2] VGND VGND VPWR VPWR _09085_/B sky130_fd_sc_hd__buf_4
X_10024_ _10411_/CLK _10024_/D repeater407/X VGND VGND VPWR VPWR _10024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput121 sram_ro_data[6] VGND VGND VPWR VPWR input121/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput187 wb_dat_i[2] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[1] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_dat_i[0] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput198 wb_sel_i[0] VGND VGND VPWR VPWR _05490_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06950_ _10189_/Q VGND VGND VPWR VPWR _06950_/Y sky130_fd_sc_hd__inv_2
X_05901_ _10165_/Q _05897_/X _09580_/X _05899_/X VGND VGND VPWR VPWR _10165_/D sky130_fd_sc_hd__a22o_1
X_06881_ _09859_/Q VGND VGND VPWR VPWR _06881_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08620_ _08620_/A VGND VGND VPWR VPWR _09223_/B sky130_fd_sc_hd__buf_2
XFILLER_94_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05832_ _05832_/A VGND VGND VPWR VPWR _05832_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08551_ _08571_/C _08556_/D _08695_/A VGND VGND VPWR VPWR _08552_/B sky130_fd_sc_hd__or3_4
X_05763_ _05764_/A VGND VGND VPWR VPWR _05763_/X sky130_fd_sc_hd__clkbuf_2
X_05694_ _10287_/Q _05690_/X _09578_/X _05692_/X VGND VGND VPWR VPWR _10287_/D sky130_fd_sc_hd__a22o_1
X_08482_ _08482_/A VGND VGND VPWR VPWR _09082_/A sky130_fd_sc_hd__inv_2
X_07502_ _07502_/A VGND VGND VPWR VPWR _07502_/X sky130_fd_sc_hd__buf_4
X_07433_ _07159_/X _07426_/X _09753_/Q _07428_/X VGND VGND VPWR VPWR _09753_/D sky130_fd_sc_hd__o22a_1
XFILLER_167_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07364_ _10207_/Q VGND VGND VPWR VPWR _07364_/Y sky130_fd_sc_hd__clkinv_2
X_09103_ _09103_/A _09103_/B VGND VGND VPWR VPWR _09103_/X sky130_fd_sc_hd__or2_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07295_ input53/X _05114_/X _10452_/Q _05089_/X _07294_/X VGND VGND VPWR VPWR _07303_/B
+ sky130_fd_sc_hd__a221o_1
X_06315_ _06315_/A VGND VGND VPWR VPWR _06316_/A sky130_fd_sc_hd__inv_2
XFILLER_175_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09034_ _09374_/A _09312_/A _09034_/C VGND VGND VPWR VPWR _09036_/A sky130_fd_sc_hd__or3_1
X_06246_ _07546_/C VGND VGND VPWR VPWR _07612_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06177_ _06177_/A VGND VGND VPWR VPWR _06177_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05128_ _05163_/B _05349_/A VGND VGND VPWR VPWR _05129_/A sky130_fd_sc_hd__nor2_2
X_09936_ _10310_/CLK _09936_/D repeater404/X VGND VGND VPWR VPWR _09936_/Q sky130_fd_sc_hd__dfrtp_1
X_05059_ _05059_/A VGND VGND VPWR VPWR _05059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09867_ _10382_/CLK _09867_/D _06452_/X VGND VGND VPWR VPWR _09867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08806_/Y _08808_/X _08808_/A _08804_/A _08817_/X VGND VGND VPWR VPWR _08821_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09798_ _10512_/CLK _09798_/D _07492_/B VGND VGND VPWR VPWR _09798_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _08749_/A VGND VGND VPWR VPWR _08750_/C sky130_fd_sc_hd__inv_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_5_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10411_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10007_ _10500_/CLK _10007_/D repeater407/X VGND VGND VPWR VPWR _10007_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06100_ _10044_/Q _06097_/X _09581_/X _06099_/X VGND VGND VPWR VPWR _10044_/D sky130_fd_sc_hd__a22o_1
X_07080_ _10053_/Q VGND VGND VPWR VPWR _07080_/Y sky130_fd_sc_hd__inv_4
X_06031_ _10085_/Q _06025_/X _09545_/A1 _06027_/X VGND VGND VPWR VPWR _10085_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07982_ _06951_/Y _07816_/A _06939_/Y _07817_/A _07981_/X VGND VGND VPWR VPWR _07987_/B
+ sky130_fd_sc_hd__o221a_1
X_09721_ _10507_/Q _09495_/A VGND VGND VPWR VPWR _09721_/Z sky130_fd_sc_hd__ebufn_1
X_06933_ _10476_/Q _06933_/B VGND VGND VPWR VPWR _06933_/Y sky130_fd_sc_hd__nand2_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06864_ _09899_/Q VGND VGND VPWR VPWR _06864_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09652_ _08347_/X _09805_/Q _09773_/Q VGND VGND VPWR VPWR _09652_/X sky130_fd_sc_hd__mux2_1
X_09583_ _09580_/X _10306_/Q _09677_/S VGND VGND VPWR VPWR _09583_/X sky130_fd_sc_hd__mux2_1
X_05815_ _10215_/Q _05809_/X _09547_/A1 _05811_/X VGND VGND VPWR VPWR _10215_/D sky130_fd_sc_hd__a22o_1
X_08603_ _09184_/A _08603_/B VGND VGND VPWR VPWR _08603_/X sky130_fd_sc_hd__or2_1
X_06795_ _06790_/Y _06439_/B _06791_/Y _06481_/B _06794_/X VGND VGND VPWR VPWR _06814_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05746_ _10254_/Q _05741_/X _09661_/A1 _05742_/Y VGND VGND VPWR VPWR _10254_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08534_ _08942_/B VGND VGND VPWR VPWR _08581_/B sky130_fd_sc_hd__buf_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05677_ _05794_/A _05677_/B VGND VGND VPWR VPWR _05679_/A sky130_fd_sc_hd__or2_4
X_08465_ _08661_/A VGND VGND VPWR VPWR _08466_/A sky130_fd_sc_hd__buf_2
X_08396_ _08884_/A VGND VGND VPWR VPWR _08556_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_168_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07416_ _07414_/Y _04870_/A _07415_/Y _05433_/A VGND VGND VPWR VPWR _07416_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07347_ _07345_/Y _05474_/B _07346_/Y _05748_/A VGND VGND VPWR VPWR _07347_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07278_ _09851_/Q VGND VGND VPWR VPWR _07278_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ _09204_/A _09007_/X _08925_/A _09023_/A _09016_/X VGND VGND VPWR VPWR _09017_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06229_ _07602_/D VGND VGND VPWR VPWR _07612_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09919_ _09919_/CLK _09919_/D repeater409/X VGND VGND VPWR VPWR _09919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10487_ _10487_/CLK _10487_/D _05034_/A VGND VGND VPWR VPWR _10487_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05600_ _10339_/Q _05596_/X _06683_/B1 _05597_/Y VGND VGND VPWR VPWR _10339_/D sky130_fd_sc_hd__a22o_1
X_06580_ _06580_/A VGND VGND VPWR VPWR _06581_/S sky130_fd_sc_hd__clkbuf_1
X_05531_ _05531_/A VGND VGND VPWR VPWR _05531_/X sky130_fd_sc_hd__clkbuf_2
X_05462_ _06646_/A VGND VGND VPWR VPWR _06663_/A sky130_fd_sc_hd__clkbuf_2
X_08250_ _05360_/Y _08199_/X _05296_/Y _08200_/X _08249_/X VGND VGND VPWR VPWR _08255_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07201_ _10195_/Q VGND VGND VPWR VPWR _07201_/Y sky130_fd_sc_hd__clkinv_4
X_08181_ _06809_/Y _08179_/X _06792_/Y _08180_/X VGND VGND VPWR VPWR _08181_/X sky130_fd_sc_hd__o22a_1
X_07132_ _10261_/Q VGND VGND VPWR VPWR _09507_/A sky130_fd_sc_hd__clkinv_4
X_05393_ _05406_/A VGND VGND VPWR VPWR _05394_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07063_ _09499_/A _05839_/B _07059_/Y _06351_/B _07062_/X VGND VGND VPWR VPWR _07063_/X
+ sky130_fd_sc_hd__o221a_4
Xoutput233 _09518_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput222 _09498_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_06014_ _06014_/A VGND VGND VPWR VPWR _06014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput211 _09478_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput244 _09470_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput266 _09728_/Z VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput255 _09718_/Z VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput277 _09703_/Z VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_2
Xoutput299 _10433_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_2
Xoutput288 _07495_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_2
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07965_ _07012_/Y _07779_/A _07963_/Y _07781_/A _07964_/X VGND VGND VPWR VPWR _07965_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06916_ _10049_/Q _05084_/Y _10111_/Q _05094_/Y _06915_/X VGND VGND VPWR VPWR _06935_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09704_ _10280_/Q _09461_/A VGND VGND VPWR VPWR _09704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07896_ _07402_/Y _07755_/X _07365_/Y _07802_/X VGND VGND VPWR VPWR _07896_/X sky130_fd_sc_hd__o22a_1
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09635_ _09634_/X _09891_/Q _09776_/Q VGND VGND VPWR VPWR _09635_/X sky130_fd_sc_hd__mux2_1
X_06847_ input40/X _06770_/A _10456_/Q _05089_/X VGND VGND VPWR VPWR _06847_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06778_ _10478_/Q _06933_/B input50/X _06697_/X _06777_/X VGND VGND VPWR VPWR _06789_/A
+ sky130_fd_sc_hd__a221o_2
X_09566_ _07049_/Y input2/X input1/X VGND VGND VPWR VPWR _09566_/X sky130_fd_sc_hd__mux2_4
X_09497_ _09497_/A VGND VGND VPWR VPWR _09498_/A sky130_fd_sc_hd__clkbuf_1
X_05729_ _05730_/A VGND VGND VPWR VPWR _05729_/X sky130_fd_sc_hd__clkbuf_2
X_08517_ _08968_/B VGND VGND VPWR VPWR _08520_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08448_ _08621_/C VGND VGND VPWR VPWR _09372_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ _08485_/A _08379_/B _08492_/C VGND VGND VPWR VPWR _08621_/C sky130_fd_sc_hd__or3_4
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ _10411_/CLK _10410_/D repeater407/X VGND VGND VPWR VPWR _10410_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10341_ _10341_/CLK _10341_/D repeater409/X VGND VGND VPWR VPWR _10341_/Q sky130_fd_sc_hd__dfstp_2
X_10272_ _10504_/CLK _10272_/D repeater403/X VGND VGND VPWR VPWR _10272_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10504_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10062_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07750_ _06875_/Y _07749_/X _06885_/Y _07629_/X VGND VGND VPWR VPWR _07750_/X sky130_fd_sc_hd__o22a_1
X_04962_ _09678_/X _04959_/Y _09536_/A3 _10467_/Q _04960_/X VGND VGND VPWR VPWR _10467_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06701_ _06701_/A _06701_/B _06701_/C _06701_/D VGND VGND VPWR VPWR _06758_/A sky130_fd_sc_hd__or4_4
X_04893_ _10492_/Q _04887_/X _09547_/A1 _04889_/X VGND VGND VPWR VPWR _10492_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07681_ _07189_/Y _07639_/X _07190_/Y _07641_/X _07680_/X VGND VGND VPWR VPWR _07684_/C
+ sky130_fd_sc_hd__o221a_1
X_09420_ _09420_/A _09420_/B _09420_/C _09420_/D VGND VGND VPWR VPWR _09421_/B sky130_fd_sc_hd__or4_1
XFILLER_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06632_ _06632_/A VGND VGND VPWR VPWR _09798_/D sky130_fd_sc_hd__clkbuf_1
X_09351_ _08808_/X _09096_/B _09307_/C _09062_/A _09284_/C VGND VGND VPWR VPWR _09389_/D
+ sky130_fd_sc_hd__a2111o_1
X_06563_ _09808_/Q _09807_/Q _09809_/Q VGND VGND VPWR VPWR _06563_/X sky130_fd_sc_hd__o21a_1
X_05514_ _05518_/A VGND VGND VPWR VPWR _05515_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08302_ _07059_/Y _08193_/A _07061_/Y _08194_/A _08301_/X VGND VGND VPWR VPWR _08309_/A
+ sky130_fd_sc_hd__o221a_1
X_09282_ _08897_/B _09048_/X _09046_/B _08957_/B _09058_/B VGND VGND VPWR VPWR _09284_/C
+ sky130_fd_sc_hd__o221ai_2
X_06494_ _06635_/A _06494_/B VGND VGND VPWR VPWR _06496_/A sky130_fd_sc_hd__or2_2
X_08233_ _06722_/Y _08207_/X _06719_/Y _08208_/X VGND VGND VPWR VPWR _08233_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05445_ _10398_/Q _05436_/A _09659_/A1 _05437_/A VGND VGND VPWR VPWR _10398_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08164_ _06887_/Y _08074_/X _06863_/Y _08075_/X _08163_/X VGND VGND VPWR VPWR _08171_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05376_ _06602_/B VGND VGND VPWR VPWR _05376_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08095_ _08214_/A VGND VGND VPWR VPWR _08095_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07115_ _10066_/Q VGND VGND VPWR VPWR _09489_/A sky130_fd_sc_hd__inv_6
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07046_ input46/X _06697_/X input6/X _06838_/X _07045_/X VGND VGND VPWR VPWR _07047_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08997_ _08997_/A VGND VGND VPWR VPWR _09425_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07948_ _10340_/Q VGND VGND VPWR VPWR _07948_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07879_ _05315_/Y _07818_/X _07878_/Y _07819_/X VGND VGND VPWR VPWR _07879_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09618_ _07717_/Y _10332_/Q _09682_/S VGND VGND VPWR VPWR _09618_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09549_ hold46/A _10301_/Q _09677_/S VGND VGND VPWR VPWR _09549_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10324_ _10510_/CLK _10324_/D _05034_/A VGND VGND VPWR VPWR _10324_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10255_ _10257_/CLK _10255_/D repeater407/X VGND VGND VPWR VPWR _10255_/Q sky130_fd_sc_hd__dfstp_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10186_ _10191_/CLK _10186_/D repeater410/X VGND VGND VPWR VPWR _10186_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05230_ _09969_/Q VGND VGND VPWR VPWR _07881_/A sky130_fd_sc_hd__clkinv_4
X_05161_ _06066_/B VGND VGND VPWR VPWR _05162_/A sky130_fd_sc_hd__inv_2
X_05092_ _05164_/B VGND VGND VPWR VPWR _06630_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08920_ _08921_/B _08933_/A VGND VGND VPWR VPWR _09283_/B sky130_fd_sc_hd__nor2_1
X_08851_ _08851_/A _08851_/B VGND VGND VPWR VPWR _09342_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07802_ _07802_/A VGND VGND VPWR VPWR _07802_/X sky130_fd_sc_hd__buf_2
X_05994_ _05995_/A VGND VGND VPWR VPWR _05994_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08782_ _08783_/B VGND VGND VPWR VPWR _08782_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07733_ _06942_/Y _07652_/X _07010_/Y _07653_/X VGND VGND VPWR VPWR _07733_/X sky130_fd_sc_hd__o22a_1
X_04945_ _10472_/Q _04936_/A _09536_/A3 _04937_/A VGND VGND VPWR VPWR _10472_/D sky130_fd_sc_hd__a22o_1
X_04876_ _10498_/Q _04872_/X _06683_/B1 _04873_/Y VGND VGND VPWR VPWR _10498_/D sky130_fd_sc_hd__a22o_1
X_07664_ _07377_/Y _06232_/X _07412_/Y _07533_/A _07663_/X VGND VGND VPWR VPWR _07671_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09403_ _09425_/A _09401_/X _09347_/Y _09402_/Y VGND VGND VPWR VPWR _09403_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06615_ _06615_/A VGND VGND VPWR VPWR _06615_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07595_ _07595_/A _07595_/B _07595_/C _07595_/D VGND VGND VPWR VPWR _07616_/B sky130_fd_sc_hd__and4_1
X_09334_ _08645_/A _08809_/B _09336_/B _09105_/A _09103_/B VGND VGND VPWR VPWR _09334_/X
+ sky130_fd_sc_hd__o311a_1
X_06546_ _09823_/Q _06539_/X _09658_/A1 _06541_/X VGND VGND VPWR VPWR _09823_/D sky130_fd_sc_hd__a22o_1
X_06477_ _09864_/Q _06473_/X _09576_/X _06474_/Y VGND VGND VPWR VPWR _09864_/D sky130_fd_sc_hd__a22o_1
X_09265_ _09265_/A _09265_/B VGND VGND VPWR VPWR _09421_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09196_ _09196_/A VGND VGND VPWR VPWR _09196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08216_ _06804_/Y _08211_/X _07823_/A _08212_/X _08215_/X VGND VGND VPWR VPWR _08217_/D
+ sky130_fd_sc_hd__o221a_1
X_05428_ _05428_/A VGND VGND VPWR VPWR _05428_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08147_ _06979_/Y _08080_/X _06927_/Y _08081_/X _08146_/X VGND VGND VPWR VPWR _08152_/B
+ sky130_fd_sc_hd__o221a_1
X_05359_ _05359_/A _05359_/B VGND VGND VPWR VPWR _06528_/A sky130_fd_sc_hd__or2_1
XFILLER_134_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08078_ _07344_/Y _08076_/X _07326_/Y _08077_/X VGND VGND VPWR VPWR _08078_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07029_ _07029_/A _07029_/B _07028_/X VGND VGND VPWR VPWR _07030_/A sky130_fd_sc_hd__or3b_2
XFILLER_121_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10040_ _10404_/CLK _10040_/D hold41/X VGND VGND VPWR VPWR _10040_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 hold9/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 _05297_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10307_ _10508_/CLK _10307_/D repeater402/X VGND VGND VPWR VPWR _10307_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10238_ _10238_/CLK _10238_/D repeater403/X VGND VGND VPWR VPWR _10238_/Q sky130_fd_sc_hd__dfstp_1
X_10169_ _10491_/CLK _10169_/D repeater403/X VGND VGND VPWR VPWR _10169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06400_ _09902_/Q _06394_/X _09574_/X _06395_/Y VGND VGND VPWR VPWR _09902_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ _07375_/Y _06206_/B _07376_/Y _05883_/B _07379_/X VGND VGND VPWR VPWR _07393_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06331_ _06331_/A VGND VGND VPWR VPWR _06331_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09050_ _08977_/A _09057_/B _09277_/A _08977_/C _09015_/B VGND VGND VPWR VPWR _09058_/A
+ sky130_fd_sc_hd__o32a_1
X_06262_ _09778_/Q _06262_/B _06288_/A VGND VGND VPWR VPWR _06262_/X sky130_fd_sc_hd__and3_1
X_05213_ _05213_/A _05213_/B _09672_/X VGND VGND VPWR VPWR _05277_/A sky130_fd_sc_hd__or3_4
X_08001_ _08043_/B VGND VGND VPWR VPWR _08032_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06193_ _07989_/B VGND VGND VPWR VPWR _06193_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05144_ _05144_/A VGND VGND VPWR VPWR _05144_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05075_ _05638_/C VGND VGND VPWR VPWR _06770_/A sky130_fd_sc_hd__inv_2
X_09952_ _10191_/CLK _09952_/D repeater405/X VGND VGND VPWR VPWR _09952_/Q sky130_fd_sc_hd__dfrtp_1
X_08903_ _08906_/B VGND VGND VPWR VPWR _08943_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09883_ _10023_/CLK _09883_/D repeater409/X VGND VGND VPWR VPWR _09883_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A _09286_/A _09067_/A _09442_/A VGND VGND VPWR VPWR _08838_/A sky130_fd_sc_hd__or4_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08765_ _09223_/B _09145_/B _08764_/Y VGND VGND VPWR VPWR _08767_/A sky130_fd_sc_hd__o21ai_1
X_05977_ _10117_/Q _05970_/A _09576_/X _05971_/A VGND VGND VPWR VPWR _10117_/D sky130_fd_sc_hd__a22o_1
Xrepeater396 _09576_/X VGND VGND VPWR VPWR _09660_/A1 sky130_fd_sc_hd__buf_12
XFILLER_122_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07716_ _07716_/A _07716_/B _07716_/C _07716_/D VGND VGND VPWR VPWR _07717_/C sky130_fd_sc_hd__and4_1
XFILLER_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08696_ _09231_/A _09225_/A VGND VGND VPWR VPWR _08697_/B sky130_fd_sc_hd__or2_1
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04928_ _09536_/A3 _10480_/Q _04928_/S VGND VGND VPWR VPWR _04929_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04859_ _10502_/Q _04851_/A _09549_/X _04852_/A VGND VGND VPWR VPWR _10502_/D sky130_fd_sc_hd__o22a_1
X_07647_ _07807_/A VGND VGND VPWR VPWR _07647_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07578_ _05302_/Y _07777_/A _05285_/Y _07778_/A _07577_/X VGND VGND VPWR VPWR _07616_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06529_ _06635_/A _06529_/B VGND VGND VPWR VPWR _06531_/A sky130_fd_sc_hd__or2_1
X_09317_ _09317_/A _09317_/B VGND VGND VPWR VPWR _09419_/B sky130_fd_sc_hd__or2_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ _09248_/A _09433_/C _09247_/X VGND VGND VPWR VPWR _09417_/D sky130_fd_sc_hd__or3b_2
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09179_ _09247_/C VGND VGND VPWR VPWR _09179_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput111 sram_ro_data[26] VGND VGND VPWR VPWR input111/X sky130_fd_sc_hd__clkbuf_2
Xinput100 sram_ro_data[16] VGND VGND VPWR VPWR input100/X sky130_fd_sc_hd__clkbuf_2
Xinput144 wb_adr_i[20] VGND VGND VPWR VPWR _08492_/B sky130_fd_sc_hd__buf_2
Xinput133 wb_adr_i[10] VGND VGND VPWR VPWR _08402_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput122 sram_ro_data[7] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_2
X_10023_ _10023_/CLK _10023_/D _05034_/A VGND VGND VPWR VPWR _10023_/Q sky130_fd_sc_hd__dfrtp_1
Xinput177 wb_dat_i[20] VGND VGND VPWR VPWR _08365_/B sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_dat_i[10] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_adr_i[30] VGND VGND VPWR VPWR _06461_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput199 wb_sel_i[1] VGND VGND VPWR VPWR _05489_/B sky130_fd_sc_hd__clkbuf_1
Xinput188 wb_dat_i[30] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05900_ _10166_/Q _05897_/X _09581_/X _05899_/X VGND VGND VPWR VPWR _10166_/D sky130_fd_sc_hd__a22o_1
X_06880_ _06880_/A _06880_/B _06880_/C _06880_/D VGND VGND VPWR VPWR _06880_/X sky130_fd_sc_hd__and4_2
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05831_ _05832_/A VGND VGND VPWR VPWR _05831_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05762_ _05794_/A _05762_/B VGND VGND VPWR VPWR _05764_/A sky130_fd_sc_hd__or2_2
X_08550_ _08813_/A VGND VGND VPWR VPWR _08553_/B sky130_fd_sc_hd__inv_2
X_05693_ _10288_/Q _05690_/X _09579_/X _05692_/X VGND VGND VPWR VPWR _10288_/D sky130_fd_sc_hd__a22o_1
X_08481_ _08787_/B _09372_/B _08621_/C VGND VGND VPWR VPWR _08482_/A sky130_fd_sc_hd__or3_1
X_07501_ _10297_/Q input74/X VGND VGND VPWR VPWR _07502_/A sky130_fd_sc_hd__and2b_1
X_07432_ _07030_/X _07426_/X _09754_/Q _07428_/X VGND VGND VPWR VPWR _09754_/D sky130_fd_sc_hd__o22a_2
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07363_ _09961_/Q VGND VGND VPWR VPWR _07363_/Y sky130_fd_sc_hd__clkinv_2
X_09102_ _09102_/A _09102_/B _09102_/C _09102_/D VGND VGND VPWR VPWR _09103_/B sky130_fd_sc_hd__or4_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07294_ _10470_/Q _04947_/Y input101/X _05153_/A VGND VGND VPWR VPWR _07294_/X sky130_fd_sc_hd__a22o_1
X_06314_ _06315_/A VGND VGND VPWR VPWR _06314_/X sky130_fd_sc_hd__clkbuf_2
X_09033_ _08504_/B _09000_/B _09032_/Y VGND VGND VPWR VPWR _09034_/C sky130_fd_sc_hd__o21ai_1
X_06245_ _09989_/Q _06245_/B VGND VGND VPWR VPWR _07546_/C sky130_fd_sc_hd__or2_1
X_06176_ _06176_/A _09777_/Q VGND VGND VPWR VPWR _06177_/A sky130_fd_sc_hd__or2_2
XFILLER_190_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05127_ _05297_/B VGND VGND VPWR VPWR _05349_/A sky130_fd_sc_hd__buf_4
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09935_ _10310_/CLK _09935_/D repeater404/X VGND VGND VPWR VPWR _09935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05058_ _05378_/A VGND VGND VPWR VPWR _05059_/A sky130_fd_sc_hd__clkbuf_1
X_09866_ _10283_/CLK _09866_/D repeater406/X VGND VGND VPWR VPWR _09866_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08817_ _09102_/C _08494_/A _09101_/A _08811_/X _08816_/X VGND VGND VPWR VPWR _08817_/X
+ sky130_fd_sc_hd__a41o_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09797_ _10483_/CLK _09797_/D _05034_/A VGND VGND VPWR VPWR _09797_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08775_/A VGND VGND VPWR VPWR _08753_/B sky130_fd_sc_hd__inv_2
XFILLER_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08809_/B _08679_/B VGND VGND VPWR VPWR _08807_/A sky130_fd_sc_hd__or2_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10006_ _10006_/CLK _10006_/D repeater407/X VGND VGND VPWR VPWR _10006_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06030_ _10086_/Q _06025_/X _09579_/X _06027_/X VGND VGND VPWR VPWR _10086_/D sky130_fd_sc_hd__a22o_1
XFILLER_126_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07981_ _06956_/Y _07818_/A _07980_/Y _07659_/A VGND VGND VPWR VPWR _07981_/X sky130_fd_sc_hd__o22a_1
X_09720_ _10506_/Q _09493_/A VGND VGND VPWR VPWR _09720_/Z sky130_fd_sc_hd__ebufn_1
X_06932_ _09964_/Q VGND VGND VPWR VPWR _06932_/Y sky130_fd_sc_hd__inv_4
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06863_ _10216_/Q VGND VGND VPWR VPWR _06863_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09651_ _08345_/X _09804_/Q _09773_/Q VGND VGND VPWR VPWR _09651_/X sky130_fd_sc_hd__mux2_1
X_05814_ _10216_/Q _05809_/X _09579_/X _05811_/X VGND VGND VPWR VPWR _10216_/D sky130_fd_sc_hd__a22o_1
X_09582_ _07505_/Y _10356_/Q _10299_/Q VGND VGND VPWR VPWR _09582_/X sky130_fd_sc_hd__mux2_1
X_08602_ _09082_/A _08602_/B VGND VGND VPWR VPWR _08603_/B sky130_fd_sc_hd__or2_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06794_ _06792_/Y _05794_/B _06793_/Y _06206_/B VGND VGND VPWR VPWR _06794_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05745_ _10255_/Q _05741_/X _06683_/B1 _05742_/Y VGND VGND VPWR VPWR _10255_/D sky130_fd_sc_hd__a22o_1
X_08533_ _08921_/C _08936_/A VGND VGND VPWR VPWR _08942_/B sky130_fd_sc_hd__or2_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _10382_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08464_ _08684_/A VGND VGND VPWR VPWR _08661_/A sky130_fd_sc_hd__clkbuf_2
X_05676_ _05806_/A VGND VGND VPWR VPWR _05794_/A sky130_fd_sc_hd__clkbuf_4
X_08395_ _08633_/A VGND VGND VPWR VPWR _08884_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07415_ _10399_/Q VGND VGND VPWR VPWR _07415_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07346_ _10246_/Q VGND VGND VPWR VPWR _07346_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07277_ _10078_/Q VGND VGND VPWR VPWR _07277_/Y sky130_fd_sc_hd__inv_2
X_09016_ _09014_/X _09388_/B _09304_/A _09016_/D VGND VGND VPWR VPWR _09016_/X sky130_fd_sc_hd__and4bb_1
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06228_ _09993_/Q _06228_/B VGND VGND VPWR VPWR _07602_/D sky130_fd_sc_hd__or2_2
XFILLER_163_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06159_ _10018_/Q _06155_/X _09580_/X _06157_/X VGND VGND VPWR VPWR _10018_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09918_ _09919_/CLK _09918_/D repeater409/X VGND VGND VPWR VPWR _09918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09849_ _10283_/CLK _09849_/D repeater406/X VGND VGND VPWR VPWR _09849_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10486_ _10486_/CLK _10486_/D _05034_/A VGND VGND VPWR VPWR _10486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05530_ _05530_/A VGND VGND VPWR VPWR _05531_/A sky130_fd_sc_hd__inv_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05461_ _09695_/X _05449_/X _10394_/Q _05451_/X VGND VGND VPWR VPWR _10394_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07200_ _10239_/Q VGND VGND VPWR VPWR _07200_/Y sky130_fd_sc_hd__inv_2
X_08180_ _08180_/A VGND VGND VPWR VPWR _08180_/X sky130_fd_sc_hd__buf_2
X_05392_ _09809_/Q _09770_/Q input58/X _05389_/Y _05391_/X VGND VGND VPWR VPWR _10419_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_158_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07131_ _09489_/A _06893_/B _07118_/X _07124_/X _07130_/X VGND VGND VPWR VPWR _07157_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07062_ _07060_/Y _06635_/B _07061_/Y _05785_/B VGND VGND VPWR VPWR _07062_/X sky130_fd_sc_hd__o22a_1
Xoutput234 _09520_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput223 _09500_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_06013_ _06013_/A VGND VGND VPWR VPWR _06014_/A sky130_fd_sc_hd__inv_2
Xoutput212 _09480_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_114_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput245 _09559_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput256 _09562_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_2
Xoutput267 _09701_/Z VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_141_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput278 _09704_/Z VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_2
Xoutput289 _07495_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_2
X_07964_ _06996_/Y _07782_/A _07006_/Y _07783_/A VGND VGND VPWR VPWR _07964_/X sky130_fd_sc_hd__o22a_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06915_ input24/X _06704_/X _10455_/Q _05089_/X VGND VGND VPWR VPWR _06915_/X sky130_fd_sc_hd__a22o_1
X_07895_ _10046_/Q VGND VGND VPWR VPWR _07895_/Y sky130_fd_sc_hd__clkinv_4
X_09703_ _10279_/Q _09459_/A VGND VGND VPWR VPWR _09703_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09634_ _07962_/Y _10327_/Q _09682_/S VGND VGND VPWR VPWR _09634_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06846_ input49/X _06697_/X input120/X _06696_/X _06845_/X VGND VGND VPWR VPWR _06855_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09565_ _10288_/Q input91/X input76/X VGND VGND VPWR VPWR _09565_/X sky130_fd_sc_hd__mux2_2
X_06777_ input107/X _05153_/A _09558_/X _06633_/A VGND VGND VPWR VPWR _06777_/X sky130_fd_sc_hd__a22o_1
X_09496_ _09496_/A VGND VGND VPWR VPWR _09496_/X sky130_fd_sc_hd__clkbuf_1
X_05728_ _05794_/A _05728_/B VGND VGND VPWR VPWR _05730_/A sky130_fd_sc_hd__or2_4
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_csclk clkbuf_leaf_4_csclk/A VGND VGND VPWR VPWR _10500_/CLK sky130_fd_sc_hd__clkbuf_16
X_08516_ _09029_/A _09103_/A VGND VGND VPWR VPWR _08968_/B sky130_fd_sc_hd__or2_1
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05659_ _10304_/Q _05653_/X _09578_/X _05655_/X VGND VGND VPWR VPWR _10304_/D sky130_fd_sc_hd__a22o_1
X_08447_ _08883_/B _09336_/B VGND VGND VPWR VPWR _09273_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08378_ _08378_/A VGND VGND VPWR VPWR _08379_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07329_ _07327_/Y _06537_/A _07328_/Y _05419_/B VGND VGND VPWR VPWR _07329_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10340_ _10341_/CLK _10340_/D repeater409/X VGND VGND VPWR VPWR _10340_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10271_ _10313_/CLK _10271_/D repeater403/X VGND VGND VPWR VPWR _10271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10469_ _10471_/CLK _10469_/D repeater409/X VGND VGND VPWR VPWR _10469_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04961_ _09678_/X _04959_/Y _06684_/B1 _10468_/Q _04960_/X VGND VGND VPWR VPWR _10468_/D
+ sky130_fd_sc_hd__a32o_1
X_06700_ input122/X _06696_/X input51/X _06697_/X _06699_/X VGND VGND VPWR VPWR _06701_/D
+ sky130_fd_sc_hd__a221o_1
X_07680_ _07276_/Y _07568_/B _07270_/Y _07642_/X VGND VGND VPWR VPWR _07680_/X sky130_fd_sc_hd__o22a_4
X_04892_ _10493_/Q _04887_/X _09579_/X _04889_/X VGND VGND VPWR VPWR _10493_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06631_ _09536_/A3 _09798_/Q _06631_/S VGND VGND VPWR VPWR _06632_/A sky130_fd_sc_hd__mux2_1
X_09350_ _09433_/B VGND VGND VPWR VPWR _09350_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06562_ _09814_/Q _09813_/Q VGND VGND VPWR VPWR _06601_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05513_ _05513_/A VGND VGND VPWR VPWR _10381_/D sky130_fd_sc_hd__clkbuf_1
X_09281_ _09352_/A _09280_/X _08918_/A _09058_/C VGND VGND VPWR VPWR _09431_/A sky130_fd_sc_hd__o211ai_4
X_08301_ _07065_/Y _08195_/A _07080_/Y _08196_/A VGND VGND VPWR VPWR _08301_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08232_ _06747_/Y _08199_/X _06718_/Y _08200_/X _08231_/X VGND VGND VPWR VPWR _08237_/B
+ sky130_fd_sc_hd__o221a_1
X_06493_ _06493_/A VGND VGND VPWR VPWR _06494_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05444_ _10399_/Q _05436_/A _09661_/A1 _05437_/A VGND VGND VPWR VPWR _10399_/D sky130_fd_sc_hd__a22o_1
X_08163_ _06869_/Y _08076_/X _06893_/A _08077_/X VGND VGND VPWR VPWR _08163_/X sky130_fd_sc_hd__o22a_1
X_05375_ _06561_/A VGND VGND VPWR VPWR _06602_/B sky130_fd_sc_hd__inv_2
X_08094_ _08213_/A VGND VGND VPWR VPWR _08094_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07114_ _07114_/A _07114_/B _07114_/C _07114_/D VGND VGND VPWR VPWR _07157_/B sky130_fd_sc_hd__and4_1
XFILLER_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07045_ input29/X _05129_/X input14/X _06698_/X VGND VGND VPWR VPWR _07045_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08996_ _08996_/A VGND VGND VPWR VPWR _09432_/A sky130_fd_sc_hd__buf_2
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07947_ _07945_/Y _07639_/A _07134_/Y _07801_/A _07946_/X VGND VGND VPWR VPWR _07951_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07878_ _10123_/Q VGND VGND VPWR VPWR _07878_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09617_ _09616_/X _09882_/Q _09776_/Q VGND VGND VPWR VPWR _09617_/X sky130_fd_sc_hd__mux2_1
X_06829_ _09926_/Q VGND VGND VPWR VPWR _06829_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09548_ _10313_/Q _09579_/X _09699_/S VGND VGND VPWR VPWR _09548_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09479_ _09479_/A VGND VGND VPWR VPWR _09480_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10323_ _10405_/CLK _10323_/D hold41/X VGND VGND VPWR VPWR _10323_/Q sky130_fd_sc_hd__dfrtp_1
X_10254_ _10254_/CLK _10254_/D repeater407/X VGND VGND VPWR VPWR _10254_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10185_ _10224_/CLK _10185_/D repeater405/X VGND VGND VPWR VPWR _10185_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05160_ _05160_/A _05325_/A VGND VGND VPWR VPWR _06066_/B sky130_fd_sc_hd__or2_1
XFILLER_170_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05091_ _05091_/A VGND VGND VPWR VPWR _05091_/X sky130_fd_sc_hd__buf_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08850_ _08850_/A _09290_/A VGND VGND VPWR VPWR _08852_/A sky130_fd_sc_hd__or2_1
X_07801_ _07801_/A VGND VGND VPWR VPWR _07801_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08781_ _09233_/A _08781_/B _09092_/A VGND VGND VPWR VPWR _08783_/B sky130_fd_sc_hd__or3_2
X_05993_ _05993_/A _05993_/B VGND VGND VPWR VPWR _05995_/A sky130_fd_sc_hd__or2_2
Xclkbuf_opt_6_0_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_4_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
X_07732_ _07732_/A _07732_/B _07732_/C _07732_/D VGND VGND VPWR VPWR _07744_/B sky130_fd_sc_hd__and4_1
X_04944_ _10473_/Q _04936_/A _06684_/B1 _04937_/A VGND VGND VPWR VPWR _10473_/D sky130_fd_sc_hd__a22o_1
X_04875_ _10499_/Q _04872_/X _09658_/A1 _04873_/Y VGND VGND VPWR VPWR _10499_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07663_ _07663_/A _07770_/B VGND VGND VPWR VPWR _07663_/X sky130_fd_sc_hd__or2_1
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09402_ _09426_/C VGND VGND VPWR VPWR _09402_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06614_ _06614_/A VGND VGND VPWR VPWR _06615_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09333_ _09425_/D VGND VGND VPWR VPWR _09333_/Y sky130_fd_sc_hd__inv_2
X_07594_ _05200_/Y _07645_/A _05239_/Y _07523_/A _07593_/X VGND VGND VPWR VPWR _07595_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06545_ _09824_/Q _06539_/X _09545_/A1 _06541_/X VGND VGND VPWR VPWR _09824_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06476_ _09865_/Q _06473_/X _09550_/A0 _06474_/Y VGND VGND VPWR VPWR _09865_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09264_ _09264_/A _09339_/D _09398_/C _09342_/D VGND VGND VPWR VPWR _09270_/A sky130_fd_sc_hd__or4_2
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09195_ _09195_/A _09194_/X VGND VGND VPWR VPWR _09196_/A sky130_fd_sc_hd__or2b_1
X_08215_ _06827_/Y _08213_/X _06802_/Y _08214_/X VGND VGND VPWR VPWR _08215_/X sky130_fd_sc_hd__o22a_1
X_05427_ _05588_/A VGND VGND VPWR VPWR _05428_/A sky130_fd_sc_hd__clkbuf_1
X_08146_ _07021_/Y _08082_/X _06991_/Y _08083_/X VGND VGND VPWR VPWR _08146_/X sky130_fd_sc_hd__o22a_1
XFILLER_181_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05358_ _09828_/Q VGND VGND VPWR VPWR _05358_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08077_ _08196_/A VGND VGND VPWR VPWR _08077_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05289_ _05285_/Y _05807_/A _05287_/Y _05873_/A VGND VGND VPWR VPWR _05289_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07028_ _07028_/A _07028_/B _07028_/C _07028_/D VGND VGND VPWR VPWR _07028_/X sky130_fd_sc_hd__and4_4
Xclkbuf_leaf_22_csclk clkbuf_opt_8_0_csclk/X VGND VGND VPWR VPWR _10508_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold22 hold22/A VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_08979_ _09390_/A _08979_/B VGND VGND VPWR VPWR _08981_/A sky130_fd_sc_hd__or2_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10404_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _05968_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10306_ _10508_/CLK _10306_/D repeater402/X VGND VGND VPWR VPWR _10306_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10237_ _10238_/CLK _10237_/D repeater403/X VGND VGND VPWR VPWR _10237_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_152_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10168_ _10491_/CLK _10168_/D repeater403/X VGND VGND VPWR VPWR _10168_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10099_ _10127_/CLK _10099_/D _07492_/B VGND VGND VPWR VPWR _10099_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06330_ _06331_/A VGND VGND VPWR VPWR _06330_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06261_ _10023_/Q _10022_/Q _10021_/Q VGND VGND VPWR VPWR _06288_/A sky130_fd_sc_hd__or3_1
X_05212_ _09833_/Q VGND VGND VPWR VPWR _05212_/Y sky130_fd_sc_hd__inv_2
X_08000_ _10005_/Q _08000_/B VGND VGND VPWR VPWR _08043_/B sky130_fd_sc_hd__or2_1
X_06192_ _10004_/Q VGND VGND VPWR VPWR _08000_/B sky130_fd_sc_hd__inv_2
X_05143_ _10480_/Q _10419_/Q _10298_/Q VGND VGND VPWR VPWR _05144_/A sky130_fd_sc_hd__or3_1
XFILLER_171_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09951_ _10062_/CLK _09951_/D repeater405/X VGND VGND VPWR VPWR _09951_/Q sky130_fd_sc_hd__dfrtp_1
X_05074_ _05178_/A _05167_/A VGND VGND VPWR VPWR _05638_/C sky130_fd_sc_hd__or2_2
X_08902_ _08902_/A _08905_/B VGND VGND VPWR VPWR _08906_/B sky130_fd_sc_hd__or2_1
XFILLER_143_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09882_ _10023_/CLK _09882_/D repeater409/X VGND VGND VPWR VPWR _09882_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08833_ _08835_/A _08853_/B VGND VGND VPWR VPWR _09442_/A sky130_fd_sc_hd__nor2_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05976_ _10118_/Q _05969_/X _09550_/A0 _05971_/X VGND VGND VPWR VPWR _10118_/D sky130_fd_sc_hd__a22o_1
X_08764_ _09297_/B _08764_/B VGND VGND VPWR VPWR _08764_/Y sky130_fd_sc_hd__nor2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07715_ _09489_/A _07665_/X _07504_/Y _07666_/X _07714_/X VGND VGND VPWR VPWR _07716_/D
+ sky130_fd_sc_hd__o221a_1
X_04927_ _05346_/A _05139_/B _06630_/C VGND VGND VPWR VPWR _04928_/S sky130_fd_sc_hd__or3_1
X_08695_ _08695_/A _08695_/B _08695_/C VGND VGND VPWR VPWR _09231_/A sky130_fd_sc_hd__or3_4
Xrepeater397 _09576_/X VGND VGND VPWR VPWR _06683_/B1 sky130_fd_sc_hd__buf_12
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04858_ _10503_/Q _04851_/A _09551_/X _04852_/A VGND VGND VPWR VPWR _10503_/D sky130_fd_sc_hd__o22a_1
X_07646_ _07646_/A VGND VGND VPWR VPWR _07646_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07577_ _05354_/Y _07779_/A _05172_/Y _07781_/A _07576_/X VGND VGND VPWR VPWR _07577_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09316_ _09316_/A VGND VGND VPWR VPWR _09316_/X sky130_fd_sc_hd__clkbuf_1
X_06528_ _06528_/A VGND VGND VPWR VPWR _06529_/B sky130_fd_sc_hd__buf_2
XFILLER_193_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09247_ _09295_/A _09247_/B _09247_/C _09247_/D VGND VGND VPWR VPWR _09247_/X sky130_fd_sc_hd__or4_1
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06459_ _08412_/A _08412_/B VGND VGND VPWR VPWR _08492_/C sky130_fd_sc_hd__or2_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09178_ _09178_/A _09178_/B _09410_/A VGND VGND VPWR VPWR _09182_/A sky130_fd_sc_hd__or3_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08129_ _09469_/A _08080_/X _09493_/A _08081_/X _08128_/X VGND VGND VPWR VPWR _08134_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput101 sram_ro_data[17] VGND VGND VPWR VPWR input101/X sky130_fd_sc_hd__buf_2
Xinput145 wb_adr_i[21] VGND VGND VPWR VPWR _08485_/A sky130_fd_sc_hd__buf_2
Xinput134 wb_adr_i[11] VGND VGND VPWR VPWR _08402_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput112 sram_ro_data[27] VGND VGND VPWR VPWR input112/X sky130_fd_sc_hd__buf_2
Xinput123 sram_ro_data[8] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10022_ _10023_/CLK _10022_/D _05034_/A VGND VGND VPWR VPWR _10022_/Q sky130_fd_sc_hd__dfrtp_1
Xinput178 wb_dat_i[21] VGND VGND VPWR VPWR _08367_/B sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_dat_i[11] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_adr_i[31] VGND VGND VPWR VPWR _06461_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput189 wb_dat_i[31] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05830_ _05874_/A _05830_/B VGND VGND VPWR VPWR _05832_/A sky130_fd_sc_hd__or2_2
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05761_ _05761_/A VGND VGND VPWR VPWR _05762_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07500_ _07500_/A VGND VGND VPWR VPWR _07500_/X sky130_fd_sc_hd__buf_6
XFILLER_35_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05692_ _05692_/A VGND VGND VPWR VPWR _05692_/X sky130_fd_sc_hd__clkbuf_2
X_08480_ _08974_/B VGND VGND VPWR VPWR _09372_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07431_ _06906_/X _07426_/X _09755_/Q _07428_/X VGND VGND VPWR VPWR _09755_/D sky130_fd_sc_hd__o22a_1
XFILLER_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07362_ _09984_/Q VGND VGND VPWR VPWR _07362_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09101_ _09101_/A VGND VGND VPWR VPWR _09101_/Y sky130_fd_sc_hd__inv_2
X_06313_ _06313_/A _06313_/B VGND VGND VPWR VPWR _06315_/A sky130_fd_sc_hd__or2_4
XFILLER_175_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07293_ _10460_/Q _06853_/B _10098_/Q _05070_/Y _07292_/X VGND VGND VPWR VPWR _07303_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ _09032_/A _09311_/C _09214_/C _09405_/C VGND VGND VPWR VPWR _09032_/Y sky130_fd_sc_hd__nor4_2
X_06244_ _07524_/A VGND VGND VPWR VPWR _07611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06175_ _09775_/Q VGND VGND VPWR VPWR _06176_/A sky130_fd_sc_hd__inv_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05126_ _05595_/B VGND VGND VPWR VPWR _05126_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09934_ _10310_/CLK _09934_/D repeater403/X VGND VGND VPWR VPWR _09934_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_77_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05057_ _06572_/A VGND VGND VPWR VPWR _05378_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09865_ _10283_/CLK _09865_/D repeater406/X VGND VGND VPWR VPWR _09865_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08553_/B _09278_/A _09256_/A _08815_/Y VGND VGND VPWR VPWR _08816_/X sky130_fd_sc_hd__o31a_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _10283_/CLK _09796_/D repeater406/X VGND VGND VPWR VPWR _09796_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05959_ _10128_/Q _05953_/X _09659_/A1 _05954_/Y VGND VGND VPWR VPWR _10128_/D sky130_fd_sc_hd__a22o_1
X_08747_ _09229_/B VGND VGND VPWR VPWR _08750_/A sky130_fd_sc_hd__inv_2
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08824_/B VGND VGND VPWR VPWR _08678_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07629_ _07629_/A VGND VGND VPWR VPWR _07629_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10005_ _10006_/CLK _10005_/D repeater409/X VGND VGND VPWR VPWR _10005_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07980_ _10127_/Q VGND VGND VPWR VPWR _07980_/Y sky130_fd_sc_hd__clkinv_2
X_06931_ _06926_/Y _05874_/B _06927_/Y _05968_/B _06930_/X VGND VGND VPWR VPWR _06931_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_101_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09650_ _09777_/Q _09554_/X _09776_/Q VGND VGND VPWR VPWR _09650_/X sky130_fd_sc_hd__mux2_8
X_08601_ _08980_/C _08491_/C _08484_/Y _08600_/X VGND VGND VPWR VPWR _08602_/B sky130_fd_sc_hd__a31o_1
X_06862_ _09979_/Q VGND VGND VPWR VPWR _07770_/A sky130_fd_sc_hd__inv_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09581_ _10418_/Q _10385_/Q _10299_/Q VGND VGND VPWR VPWR _09581_/X sky130_fd_sc_hd__mux2_8
X_05813_ _10217_/Q _05809_/X _09580_/X _05811_/X VGND VGND VPWR VPWR _10217_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06793_ _10000_/Q VGND VGND VPWR VPWR _06793_/Y sky130_fd_sc_hd__clkinv_2
X_08532_ _08537_/C _09236_/A _08640_/A _08561_/B VGND VGND VPWR VPWR _08936_/A sky130_fd_sc_hd__or4_4
X_05744_ _10256_/Q _05741_/X _09577_/X _05742_/Y VGND VGND VPWR VPWR _10256_/D sky130_fd_sc_hd__a22o_1
X_08463_ _08697_/A VGND VGND VPWR VPWR _08684_/A sky130_fd_sc_hd__buf_2
X_07414_ _10497_/Q VGND VGND VPWR VPWR _07414_/Y sky130_fd_sc_hd__clkinv_2
X_05675_ _05390_/X _05592_/B _09774_/Q _10297_/Q VGND VGND VPWR VPWR _10297_/D sky130_fd_sc_hd__a31o_1
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08394_ _08561_/B VGND VGND VPWR VPWR _08633_/A sky130_fd_sc_hd__inv_2
X_07345_ _10387_/Q VGND VGND VPWR VPWR _07345_/Y sky130_fd_sc_hd__clkinv_2
X_07276_ _10161_/Q VGND VGND VPWR VPWR _07276_/Y sky130_fd_sc_hd__clkinv_2
X_09015_ _09277_/A _09015_/B VGND VGND VPWR VPWR _09304_/A sky130_fd_sc_hd__or2_2
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06227_ _06228_/B _06227_/B _07534_/A VGND VGND VPWR VPWR _06227_/Y sky130_fd_sc_hd__nor3_1
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06158_ _10019_/Q _06155_/X _09581_/X _06157_/X VGND VGND VPWR VPWR _10019_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06089_ _06089_/A VGND VGND VPWR VPWR _06089_/Y sky130_fd_sc_hd__inv_2
X_05109_ _09674_/X _05109_/B _09670_/X _05109_/D VGND VGND VPWR VPWR _05325_/A sky130_fd_sc_hd__or4_4
X_09917_ _09919_/CLK _09917_/D repeater409/X VGND VGND VPWR VPWR _09917_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09848_ _10350_/CLK _09848_/D repeater405/X VGND VGND VPWR VPWR _09848_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09779_ _10006_/CLK _09779_/D _05034_/A VGND VGND VPWR VPWR _09779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10485_ _10486_/CLK _10485_/D _05034_/A VGND VGND VPWR VPWR _10485_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05460_ _05460_/A VGND VGND VPWR VPWR _05460_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05391_ _05429_/A _05390_/X _06593_/A _10419_/Q VGND VGND VPWR VPWR _05391_/X sky130_fd_sc_hd__o31a_1
X_07130_ _09481_/A _06266_/A _07126_/Y _06551_/B _07129_/X VGND VGND VPWR VPWR _07130_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07061_ _10230_/Q VGND VGND VPWR VPWR _07061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_145_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput224 _09502_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_2
Xoutput235 _09568_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_2
X_06012_ _06013_/A VGND VGND VPWR VPWR _06012_/X sky130_fd_sc_hd__clkbuf_2
Xoutput213 _09482_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_2
Xoutput268 _09729_/Z VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_2
Xoutput257 _09719_/Z VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput246 _09709_/Z VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_99_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput279 _09705_/Z VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_2
X_07963_ _10101_/Q VGND VGND VPWR VPWR _07963_/Y sky130_fd_sc_hd__inv_2
X_07894_ _07339_/Y _07792_/X _07390_/Y _07793_/X _07893_/X VGND VGND VPWR VPWR _07901_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09702_ _10278_/Q _09455_/A VGND VGND VPWR VPWR _09702_/Z sky130_fd_sc_hd__ebufn_1
X_06914_ input105/X _05153_/X _06908_/X _06911_/X _06913_/X VGND VGND VPWR VPWR _07029_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09633_ _09632_/X _09890_/Q _09776_/Q VGND VGND VPWR VPWR _09633_/X sky130_fd_sc_hd__mux2_1
X_06845_ input66/X _06844_/X _10034_/Q _05080_/A VGND VGND VPWR VPWR _06845_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09564_ _10287_/Q input89/X input76/X VGND VGND VPWR VPWR _09564_/X sky130_fd_sc_hd__mux2_4
X_08515_ _08586_/A VGND VGND VPWR VPWR _08746_/A sky130_fd_sc_hd__buf_2
X_06776_ _06776_/A VGND VGND VPWR VPWR _06933_/B sky130_fd_sc_hd__buf_2
X_09495_ _09495_/A VGND VGND VPWR VPWR _09496_/A sky130_fd_sc_hd__clkbuf_1
X_05727_ _05727_/A VGND VGND VPWR VPWR _05728_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05658_ _10305_/Q _05653_/X _09579_/X _05655_/X VGND VGND VPWR VPWR _10305_/D sky130_fd_sc_hd__a22o_1
X_08446_ _08732_/A VGND VGND VPWR VPWR _09336_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08377_ _08965_/A VGND VGND VPWR VPWR _08999_/A sky130_fd_sc_hd__inv_2
XFILLER_139_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07328_ _10408_/Q VGND VGND VPWR VPWR _07328_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05589_ _05589_/A VGND VGND VPWR VPWR _05589_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07259_ _09822_/Q VGND VGND VPWR VPWR _07259_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10270_ _10313_/CLK _10270_/D repeater404/X VGND VGND VPWR VPWR _10270_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10468_ _10471_/CLK _10468_/D repeater409/X VGND VGND VPWR VPWR _10468_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10399_ _10404_/CLK _10399_/D repeater410/X VGND VGND VPWR VPWR _10399_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04960_ _05031_/A _04960_/B VGND VGND VPWR VPWR _04960_/X sky130_fd_sc_hd__or2_1
X_04891_ _10494_/Q _04887_/X _09580_/X _04889_/X VGND VGND VPWR VPWR _10494_/D sky130_fd_sc_hd__a22o_1
X_06630_ _06630_/A _06630_/B _06630_/C VGND VGND VPWR VPWR _06631_/S sky130_fd_sc_hd__or3_1
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06561_ _06561_/A VGND VGND VPWR VPWR _07489_/A sky130_fd_sc_hd__clkbuf_2
X_05512_ _09687_/X _10381_/Q _05512_/S VGND VGND VPWR VPWR _05513_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09280_ _08897_/B _09352_/C _08910_/X VGND VGND VPWR VPWR _09280_/X sky130_fd_sc_hd__o21a_1
X_06492_ _09854_/Q _06483_/A _09659_/A1 _06484_/A VGND VGND VPWR VPWR _09854_/D sky130_fd_sc_hd__a22o_1
X_08300_ _07067_/Y _08183_/A _08297_/X _08299_/X VGND VGND VPWR VPWR _08310_/C sky130_fd_sc_hd__o211a_1
XFILLER_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08231_ _06716_/Y _08201_/X _06725_/Y _08202_/X VGND VGND VPWR VPWR _08231_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05443_ _10400_/Q _05436_/A _09660_/A1 _05437_/A VGND VGND VPWR VPWR _10400_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05374_ _05429_/A _05429_/D _06579_/B VGND VGND VPWR VPWR _06561_/A sky130_fd_sc_hd__or3_1
Xclkbuf_opt_2_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_08162_ _06852_/Y _08064_/X _08159_/X _08161_/X VGND VGND VPWR VPWR _08172_/C sky130_fd_sc_hd__o211a_1
X_08093_ _08212_/A VGND VGND VPWR VPWR _08093_/X sky130_fd_sc_hd__clkbuf_2
X_07113_ _09485_/A _06153_/A _09483_/A _06205_/A _07112_/X VGND VGND VPWR VPWR _07114_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07044_ input128/X _05118_/Y _10484_/Q _06633_/X _07043_/X VGND VGND VPWR VPWR _07047_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08995_ _09363_/A _09318_/B VGND VGND VPWR VPWR _09385_/A sky130_fd_sc_hd__or2_2
XFILLER_114_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07946_ _07085_/Y _07512_/A _07119_/Y _07642_/A VGND VGND VPWR VPWR _07946_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07877_ _05350_/Y _07762_/X _05337_/Y _07811_/X _07876_/X VGND VGND VPWR VPWR _07885_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06828_ _10199_/Q VGND VGND VPWR VPWR _06828_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09616_ _07695_/Y _10331_/Q _09682_/S VGND VGND VPWR VPWR _09616_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09547_ _10312_/Q _09547_/A1 _09699_/S VGND VGND VPWR VPWR _09547_/X sky130_fd_sc_hd__mux2_1
X_06759_ _06759_/A VGND VGND VPWR VPWR _06759_/X sky130_fd_sc_hd__buf_6
XFILLER_169_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09478_ _09478_/A VGND VGND VPWR VPWR _09478_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08429_ _09236_/B _08568_/A VGND VGND VPWR VPWR _09247_/C sky130_fd_sc_hd__nand2_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10322_ _10405_/CLK _10322_/D hold41/X VGND VGND VPWR VPWR _10322_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10253_ _10254_/CLK _10253_/D repeater407/X VGND VGND VPWR VPWR _10253_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10184_ _10184_/CLK _10184_/D repeater407/X VGND VGND VPWR VPWR _10184_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06665__1 _09572_/A1 VGND VGND VPWR VPWR _09780_/CLK sky130_fd_sc_hd__inv_2
X_05090_ _05090_/A VGND VGND VPWR VPWR _05091_/A sky130_fd_sc_hd__inv_2
XFILLER_69_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10366_/CLK sky130_fd_sc_hd__clkbuf_16
X_08780_ _08895_/A _08786_/B _08643_/A _08814_/A VGND VGND VPWR VPWR _09092_/A sky130_fd_sc_hd__or4bb_4
XFILLER_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07800_ _10139_/Q VGND VGND VPWR VPWR _07800_/Y sky130_fd_sc_hd__inv_2
X_05992_ _05992_/A VGND VGND VPWR VPWR _05993_/B sky130_fd_sc_hd__clkbuf_4
X_07731_ _06976_/Y _07645_/X _06991_/Y _07533_/B _07730_/X VGND VGND VPWR VPWR _07732_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04943_ _10474_/Q _04936_/A _06683_/B1 _04937_/A VGND VGND VPWR VPWR _10474_/D sky130_fd_sc_hd__a22o_1
X_04874_ _10500_/Q _04872_/X _09545_/A1 _04873_/Y VGND VGND VPWR VPWR _10500_/D sky130_fd_sc_hd__a22o_1
X_07662_ _07983_/B VGND VGND VPWR VPWR _07770_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09401_ _09401_/A _09421_/D _09425_/C _09426_/D VGND VGND VPWR VPWR _09401_/X sky130_fd_sc_hd__or4_1
X_07593_ _05322_/Y _07646_/A _05273_/Y _07807_/A VGND VGND VPWR VPWR _07593_/X sky130_fd_sc_hd__o22a_1
X_06613_ _09804_/Q _06604_/X _09649_/X _06606_/X VGND VGND VPWR VPWR _09804_/D sky130_fd_sc_hd__a22o_1
X_09332_ _09418_/A _09417_/B _09415_/B _09332_/D VGND VGND VPWR VPWR _09332_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06544_ _09825_/Q _06539_/X _09579_/X _06541_/X VGND VGND VPWR VPWR _09825_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06475_ _09866_/Q _06473_/X _09578_/X _06474_/Y VGND VGND VPWR VPWR _09866_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09263_ _09263_/A _09265_/B VGND VGND VPWR VPWR _09342_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09194_ _09222_/B _09193_/X VGND VGND VPWR VPWR _09194_/X sky130_fd_sc_hd__or2b_1
X_08214_ _08214_/A VGND VGND VPWR VPWR _08214_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05426_ _10407_/Q _05420_/X _09574_/X _05421_/Y VGND VGND VPWR VPWR _10407_/D sky130_fd_sc_hd__a22o_1
X_08145_ _07022_/Y _08074_/X _06987_/Y _08075_/X _08144_/X VGND VGND VPWR VPWR _08152_/A
+ sky130_fd_sc_hd__o221a_1
X_05357_ _05357_/A _05357_/B VGND VGND VPWR VPWR _05527_/A sky130_fd_sc_hd__or2_2
XFILLER_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08076_ _08195_/A VGND VGND VPWR VPWR _08076_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05288_ _05313_/A _05351_/A VGND VGND VPWR VPWR _05873_/A sky130_fd_sc_hd__or2_1
X_07027_ _07027_/A _07027_/B _07027_/C _07027_/D VGND VGND VPWR VPWR _07028_/D sky130_fd_sc_hd__and4_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold12 hold12/A VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _08973_/X _08978_/B _08978_/C VGND VGND VPWR VPWR _08979_/B sky130_fd_sc_hd__nand3b_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold34 hold34/A VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__clkdlybuf4s50_1
X_07929_ _10125_/Q VGND VGND VPWR VPWR _07929_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_56_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _05184_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10305_ _10508_/CLK _10305_/D repeater402/X VGND VGND VPWR VPWR _10305_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10236_ _10355_/CLK _10236_/D repeater406/X VGND VGND VPWR VPWR _10236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10167_ _10313_/CLK _10167_/D repeater403/X VGND VGND VPWR VPWR _10167_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10098_ _10127_/CLK _10098_/D _07492_/B VGND VGND VPWR VPWR _10098_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06260_ _10023_/Q _10022_/Q _06260_/C _10020_/Q VGND VGND VPWR VPWR _06262_/B sky130_fd_sc_hd__or4_2
X_05211_ _05197_/Y _05748_/A _05200_/Y _06401_/A _05210_/X VGND VGND VPWR VPWR _05236_/B
+ sky130_fd_sc_hd__o221a_1
X_06191_ _06184_/Y _06190_/X _06177_/A VGND VGND VPWR VPWR _10005_/D sky130_fd_sc_hd__o21a_1
X_05142_ _05346_/A VGND VGND VPWR VPWR _05142_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05073_ _05960_/B VGND VGND VPWR VPWR _05073_/Y sky130_fd_sc_hd__clkinv_2
X_09950_ _10062_/CLK _09950_/D repeater410/X VGND VGND VPWR VPWR _09950_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08901_ _08938_/A _08921_/B _08905_/B VGND VGND VPWR VPWR _09307_/B sky130_fd_sc_hd__nor3_1
XFILLER_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09881_ _10023_/CLK _09881_/D repeater409/X VGND VGND VPWR VPWR _09881_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08832_ _08837_/A _08835_/A VGND VGND VPWR VPWR _09067_/A sky130_fd_sc_hd__nor2_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05975_ _10119_/Q _05969_/X _09578_/X _05971_/X VGND VGND VPWR VPWR _10119_/D sky130_fd_sc_hd__a22o_1
X_08763_ _08763_/A _09416_/A VGND VGND VPWR VPWR _08764_/B sky130_fd_sc_hd__or2_1
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07714_ _09503_/A _07667_/X _09501_/A _07668_/X VGND VGND VPWR VPWR _07714_/X sky130_fd_sc_hd__o22a_1
X_04926_ _06780_/A VGND VGND VPWR VPWR _05139_/B sky130_fd_sc_hd__buf_2
X_08694_ _08529_/A _08775_/A _08693_/X VGND VGND VPWR VPWR _08700_/B sky130_fd_sc_hd__o21ai_1
Xrepeater398 _09661_/A1 VGND VGND VPWR VPWR _06684_/B1 sky130_fd_sc_hd__buf_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04857_ _10504_/Q _04851_/X _09550_/X _04852_/X VGND VGND VPWR VPWR _10504_/D sky130_fd_sc_hd__o22a_1
X_07645_ _07645_/A VGND VGND VPWR VPWR _07645_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07576_ _05134_/Y _07782_/A _05283_/Y _07783_/A VGND VGND VPWR VPWR _07576_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09315_ _09315_/A _09315_/B _09315_/C _09315_/D VGND VGND VPWR VPWR _09316_/A sky130_fd_sc_hd__or4_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06527_ _09833_/Q _06518_/A _09659_/A1 _06519_/A VGND VGND VPWR VPWR _09833_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06458_ _08405_/C _08405_/D _06458_/C VGND VGND VPWR VPWR _06466_/C sky130_fd_sc_hd__or3_1
XFILLER_166_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09246_ _08491_/A _08999_/B _08750_/C _09245_/Y _09182_/B VGND VGND VPWR VPWR _09329_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05409_ _06572_/A VGND VGND VPWR VPWR _05588_/A sky130_fd_sc_hd__buf_6
XFILLER_193_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09177_ _08504_/B _08883_/A _08466_/A _09265_/A VGND VGND VPWR VPWR _09410_/A sky130_fd_sc_hd__o22ai_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06389_ _09700_/X VGND VGND VPWR VPWR _06389_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08128_ _09485_/A _08082_/X _07135_/Y _08083_/X VGND VGND VPWR VPWR _08128_/X sky130_fd_sc_hd__o22a_1
X_08059_ _08178_/A VGND VGND VPWR VPWR _08059_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 sram_ro_data[18] VGND VGND VPWR VPWR input102/X sky130_fd_sc_hd__clkbuf_2
X_10021_ _10023_/CLK _10021_/D repeater409/X VGND VGND VPWR VPWR _10021_/Q sky130_fd_sc_hd__dfrtp_1
Xinput135 wb_adr_i[12] VGND VGND VPWR VPWR _08402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput113 sram_ro_data[28] VGND VGND VPWR VPWR input113/X sky130_fd_sc_hd__buf_2
Xinput124 sram_ro_data[9] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__clkbuf_2
Xinput168 wb_dat_i[12] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_adr_i[22] VGND VGND VPWR VPWR _08412_/B sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_adr_i[3] VGND VGND VPWR VPWR _09085_/D sky130_fd_sc_hd__buf_4
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput179 wb_dat_i[22] VGND VGND VPWR VPWR _08369_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10219_ _10349_/CLK _10219_/D repeater405/X VGND VGND VPWR VPWR _10219_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05760_ _10245_/Q _05751_/A _09659_/A1 _05752_/A VGND VGND VPWR VPWR _10245_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05691_ _05691_/A VGND VGND VPWR VPWR _05692_/A sky130_fd_sc_hd__inv_2
X_07430_ _06835_/X _07426_/X _09756_/Q _07428_/X VGND VGND VPWR VPWR _09756_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07361_ _07356_/Y _05793_/A _07357_/Y _06503_/B _07360_/X VGND VGND VPWR VPWR _07374_/B
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_21_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10296_/CLK sky130_fd_sc_hd__clkbuf_16
X_09100_ _09100_/A VGND VGND VPWR VPWR _09420_/A sky130_fd_sc_hd__inv_2
X_06312_ _06312_/A VGND VGND VPWR VPWR _06313_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09031_ _09176_/A _09427_/B VGND VGND VPWR VPWR _09405_/C sky130_fd_sc_hd__or2_1
X_07292_ input21/X _06704_/A input35/X _06838_/X VGND VGND VPWR VPWR _07292_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06243_ _06243_/A _09988_/Q VGND VGND VPWR VPWR _07524_/A sky130_fd_sc_hd__or2_1
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06174_ _10007_/Q _06168_/X _09536_/A3 _06169_/Y VGND VGND VPWR VPWR _10007_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_36_csclk clkbuf_opt_5_0_csclk/X VGND VGND VPWR VPWR _10405_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05125_ _05149_/A _05338_/A VGND VGND VPWR VPWR _05595_/B sky130_fd_sc_hd__or2_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09933_ _10310_/CLK _09933_/D repeater404/X VGND VGND VPWR VPWR _09933_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_89_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05056_ _06668_/A VGND VGND VPWR VPWR _06572_/A sky130_fd_sc_hd__buf_2
X_09864_ _10157_/CLK _09864_/D repeater406/X VGND VGND VPWR VPWR _09864_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _09105_/A _09105_/B _08788_/A VGND VGND VPWR VPWR _08815_/Y sky130_fd_sc_hd__o21ai_2
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _10157_/CLK _09795_/D repeater406/X VGND VGND VPWR VPWR _09795_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05958_ _10129_/Q _05953_/X _09661_/A1 _05954_/Y VGND VGND VPWR VPWR _10129_/D sky130_fd_sc_hd__a22o_1
X_08746_ _08746_/A VGND VGND VPWR VPWR _09229_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05889_ _10172_/Q _05884_/X _09579_/X _05886_/X VGND VGND VPWR VPWR _10172_/D sky130_fd_sc_hd__a22o_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08823_/A VGND VGND VPWR VPWR _08824_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04909_ _10483_/Q _04902_/X _09545_/A1 _04904_/X VGND VGND VPWR VPWR _10483_/D sky130_fd_sc_hd__a22o_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07788_/A VGND VGND VPWR VPWR _07628_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07559_ _09989_/Q _09988_/Q _07585_/C _07562_/B VGND VGND VPWR VPWR _07583_/A sky130_fd_sc_hd__or4_1
XFILLER_166_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09229_ _09229_/A _09229_/B VGND VGND VPWR VPWR _09229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10004_ _10006_/CLK _10004_/D repeater409/X VGND VGND VPWR VPWR _10004_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06930_ _06928_/Y _05740_/B _06929_/Y _05918_/B VGND VGND VPWR VPWR _06930_/X sky130_fd_sc_hd__o22a_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08600_ _09374_/A _08600_/B VGND VGND VPWR VPWR _08600_/X sky130_fd_sc_hd__or2_1
X_06861_ _06856_/Y _04886_/B _06857_/Y _05928_/B _06860_/X VGND VGND VPWR VPWR _06880_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09580_ _10417_/Q _10384_/Q _10299_/Q VGND VGND VPWR VPWR _09580_/X sky130_fd_sc_hd__mux2_8
X_05812_ _10218_/Q _05809_/X _09581_/X _05811_/X VGND VGND VPWR VPWR _10218_/D sky130_fd_sc_hd__a22o_1
X_06792_ _10225_/Q VGND VGND VPWR VPWR _06792_/Y sky130_fd_sc_hd__inv_2
X_05743_ _10257_/Q _05741_/X _09578_/X _05742_/Y VGND VGND VPWR VPWR _10257_/D sky130_fd_sc_hd__a22o_1
X_08531_ _08582_/B VGND VGND VPWR VPWR _09024_/A sky130_fd_sc_hd__clkbuf_2
X_08462_ _09085_/C _08494_/A _08505_/A _08472_/B VGND VGND VPWR VPWR _08697_/A sky130_fd_sc_hd__or4_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05674_ _05674_/A VGND VGND VPWR VPWR _05674_/X sky130_fd_sc_hd__clkbuf_1
X_07413_ _09855_/Q VGND VGND VPWR VPWR _07413_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08393_ _08972_/A VGND VGND VPWR VPWR _09218_/A sky130_fd_sc_hd__buf_2
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07344_ _10090_/Q VGND VGND VPWR VPWR _07344_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07275_ _10151_/Q VGND VGND VPWR VPWR _07275_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09014_ _09283_/B _09014_/B _09205_/A _09013_/X VGND VGND VPWR VPWR _09014_/X sky130_fd_sc_hd__or4b_1
X_06226_ _06238_/A _07558_/A VGND VGND VPWR VPWR _07534_/A sky130_fd_sc_hd__or2_2
XFILLER_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06157_ _06157_/A VGND VGND VPWR VPWR _06157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06088_ _06089_/A VGND VGND VPWR VPWR _06088_/X sky130_fd_sc_hd__clkbuf_2
X_05108_ _05108_/A _05108_/B _05108_/C _05108_/D VGND VGND VPWR VPWR _05366_/A sky130_fd_sc_hd__or4_2
XFILLER_104_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09916_ _10397_/CLK _09916_/D repeater409/X VGND VGND VPWR VPWR _09916_/Q sky130_fd_sc_hd__dfrtp_1
X_05039_ _05713_/A _05395_/A VGND VGND VPWR VPWR _05041_/A sky130_fd_sc_hd__or2_2
XFILLER_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09847_ _10350_/CLK _09847_/D repeater405/X VGND VGND VPWR VPWR _09847_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09778_ _10023_/CLK _09778_/D _05034_/A VGND VGND VPWR VPWR _09778_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08729_ _08466_/A _09263_/A _08728_/X VGND VGND VPWR VPWR _08731_/A sky130_fd_sc_hd__o21ai_1
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10484_ _10510_/CLK _10484_/D _05034_/A VGND VGND VPWR VPWR _10484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05390_ _06585_/A VGND VGND VPWR VPWR _05390_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07060_ _09795_/Q VGND VGND VPWR VPWR _07060_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06011_ _06011_/A _06011_/B VGND VGND VPWR VPWR _06013_/A sky130_fd_sc_hd__or2_4
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput225 _09504_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_173_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput214 _09484_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput203 _09526_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_2
Xoutput258 _09720_/Z VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput236 _09569_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_160_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput247 _09710_/Z VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_99_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput269 _09730_/Z VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07962_ _07962_/A _07962_/B _07962_/C VGND VGND VPWR VPWR _07962_/Y sky130_fd_sc_hd__nand3_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09701_ _10277_/Q _09457_/A VGND VGND VPWR VPWR _09701_/Z sky130_fd_sc_hd__ebufn_1
X_07893_ _07378_/Y _07794_/X _07343_/Y _07795_/X VGND VGND VPWR VPWR _07893_/X sky130_fd_sc_hd__o22a_1
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06913_ input113/X _05112_/X _10483_/Q _06633_/X _06912_/X VGND VGND VPWR VPWR _06913_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09632_ _07937_/Y _10326_/Q _09682_/S VGND VGND VPWR VPWR _09632_/X sky130_fd_sc_hd__mux2_1
X_06844_ _06844_/A VGND VGND VPWR VPWR _06844_/X sky130_fd_sc_hd__clkbuf_4
X_09563_ _10286_/Q input81/X input79/X VGND VGND VPWR VPWR _09563_/X sky130_fd_sc_hd__mux2_4
X_08514_ _08575_/A VGND VGND VPWR VPWR _08586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06775_ _06775_/A _06775_/B _06775_/C _06775_/D VGND VGND VPWR VPWR _06834_/A sky130_fd_sc_hd__or4_2
X_09494_ _09494_/A VGND VGND VPWR VPWR _09494_/X sky130_fd_sc_hd__clkbuf_1
X_05726_ _10266_/Q _05717_/A _09544_/X _05718_/A VGND VGND VPWR VPWR _10266_/D sky130_fd_sc_hd__o22a_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05657_ _10306_/Q _05653_/X _09580_/X _05655_/X VGND VGND VPWR VPWR _10306_/D sky130_fd_sc_hd__a22o_1
X_08445_ _08710_/A VGND VGND VPWR VPWR _08732_/A sky130_fd_sc_hd__buf_2
X_08376_ _09085_/D _08472_/B _08389_/A VGND VGND VPWR VPWR _08965_/A sky130_fd_sc_hd__or3_2
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05588_ _05588_/A VGND VGND VPWR VPWR _05589_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07327_ _09821_/Q VGND VGND VPWR VPWR _07327_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07258_ _09930_/Q VGND VGND VPWR VPWR _07258_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07189_ _10031_/Q VGND VGND VPWR VPWR _07189_/Y sky130_fd_sc_hd__clkinv_2
X_06209_ _06209_/A VGND VGND VPWR VPWR _06209_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10467_ _10471_/CLK _10467_/D repeater409/X VGND VGND VPWR VPWR _10467_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_170_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10398_ _10404_/CLK _10398_/D hold41/A VGND VGND VPWR VPWR _10398_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04890_ _10495_/Q _04887_/X _09581_/X _04889_/X VGND VGND VPWR VPWR _10495_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06560_ _06560_/A VGND VGND VPWR VPWR _06560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05511_ _05511_/A VGND VGND VPWR VPWR _05511_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06491_ _09855_/Q _06483_/A _09661_/A1 _06484_/A VGND VGND VPWR VPWR _09855_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08230_ _06711_/Y _08193_/X _06745_/Y _08194_/X _08229_/X VGND VGND VPWR VPWR _08237_/A
+ sky130_fd_sc_hd__o221a_1
X_05442_ _10401_/Q _05435_/X _09658_/A1 _05437_/X VGND VGND VPWR VPWR _10401_/D sky130_fd_sc_hd__a22o_1
XFILLER_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05373_ _09807_/Q VGND VGND VPWR VPWR _06579_/B sky130_fd_sc_hd__inv_2
X_08161_ _06885_/Y _08067_/X _06856_/Y _08068_/X _08160_/X VGND VGND VPWR VPWR _08161_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08092_ _08211_/A VGND VGND VPWR VPWR _08092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07112_ _07110_/Y _05821_/B _07111_/Y _06529_/B VGND VGND VPWR VPWR _07112_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07043_ _10435_/Q _05121_/Y input118/X _06696_/X VGND VGND VPWR VPWR _07043_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08994_ _08994_/A _08994_/B VGND VGND VPWR VPWR _08994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07945_ _10048_/Q VGND VGND VPWR VPWR _07945_/Y sky130_fd_sc_hd__inv_2
X_07876_ _05218_/Y _07812_/X _05345_/Y _07813_/X VGND VGND VPWR VPWR _07876_/X sky130_fd_sc_hd__o22a_1
X_09615_ _09614_/X _09881_/Q _09776_/Q VGND VGND VPWR VPWR _09615_/X sky130_fd_sc_hd__mux2_1
X_06827_ _10251_/Q VGND VGND VPWR VPWR _06827_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_141_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ _10311_/Q _09550_/A0 _09699_/S VGND VGND VPWR VPWR _09546_/X sky130_fd_sc_hd__mux2_1
X_06758_ _06758_/A _06758_/B _06740_/X _06757_/X VGND VGND VPWR VPWR _06759_/A sky130_fd_sc_hd__or4bb_4
X_09477_ _09477_/A VGND VGND VPWR VPWR _09478_/A sky130_fd_sc_hd__clkbuf_1
X_05709_ _10276_/Q _05701_/A _09661_/X _05702_/A VGND VGND VPWR VPWR _10276_/D sky130_fd_sc_hd__o22a_1
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08428_ _08571_/C _08476_/A _09236_/A _08556_/D _08424_/X VGND VGND VPWR VPWR _08568_/A
+ sky130_fd_sc_hd__a32o_1
X_06689_ _06689_/A VGND VGND VPWR VPWR _06853_/B sky130_fd_sc_hd__buf_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08359_ _09788_/Q _08359_/B VGND VGND VPWR VPWR _08359_/X sky130_fd_sc_hd__and2_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10321_ _10405_/CLK _10321_/D hold41/X VGND VGND VPWR VPWR _10321_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10252_ _10504_/CLK _10252_/D repeater403/X VGND VGND VPWR VPWR _10252_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10183_ _10184_/CLK _10183_/D repeater407/X VGND VGND VPWR VPWR _10183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _07017_/Y _07646_/X _06961_/Y _07647_/X VGND VGND VPWR VPWR _07730_/X sky130_fd_sc_hd__o22a_1
X_05991_ _10107_/Q _05982_/A _09536_/A3 _05983_/A VGND VGND VPWR VPWR _10107_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04942_ _10475_/Q _04935_/X _09658_/A1 _04937_/X VGND VGND VPWR VPWR _10475_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04873_ _04873_/A VGND VGND VPWR VPWR _04873_/Y sky130_fd_sc_hd__inv_2
X_07661_ _07415_/Y _07656_/X _07408_/Y _07657_/X _07660_/X VGND VGND VPWR VPWR _07671_/B
+ sky130_fd_sc_hd__o221a_1
X_09400_ _09400_/A _09400_/B _09400_/C VGND VGND VPWR VPWR _09426_/D sky130_fd_sc_hd__or3_1
X_07592_ _07592_/A _07612_/B _07612_/C VGND VGND VPWR VPWR _07807_/A sky130_fd_sc_hd__or3_4
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06612_ _06612_/A VGND VGND VPWR VPWR _06612_/X sky130_fd_sc_hd__clkbuf_1
X_09331_ _09331_/A _09419_/A _09418_/B _09331_/D VGND VGND VPWR VPWR _09332_/D sky130_fd_sc_hd__or4_1
XFILLER_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06543_ _09826_/Q _06539_/X _09580_/X _06541_/X VGND VGND VPWR VPWR _09826_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06474_ _06474_/A VGND VGND VPWR VPWR _06474_/Y sky130_fd_sc_hd__inv_2
X_09262_ _09262_/A _09265_/B VGND VGND VPWR VPWR _09398_/C sky130_fd_sc_hd__nor2_1
XFILLER_159_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09193_ _09193_/A _09222_/C VGND VGND VPWR VPWR _09193_/X sky130_fd_sc_hd__or2_1
X_08213_ _08213_/A VGND VGND VPWR VPWR _08213_/X sky130_fd_sc_hd__clkbuf_2
X_05425_ _10408_/Q _05420_/X _09661_/A1 _05421_/Y VGND VGND VPWR VPWR _10408_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08144_ _06937_/Y _08076_/X _06963_/Y _08077_/X VGND VGND VPWR VPWR _08144_/X sky130_fd_sc_hd__o22a_1
X_05356_ _10370_/Q VGND VGND VPWR VPWR _05356_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05287_ _10175_/Q VGND VGND VPWR VPWR _05287_/Y sky130_fd_sc_hd__clkinv_2
X_08075_ _08194_/A VGND VGND VPWR VPWR _08075_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07026_ _07021_/Y _06153_/A _07022_/Y _06338_/A _07025_/X VGND VGND VPWR VPWR _07027_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__buf_12
X_08977_ _08977_/A _09084_/B _08977_/C VGND VGND VPWR VPWR _08978_/C sky130_fd_sc_hd__or3_1
XFILLER_152_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold24 hold24/A VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07278_/Y _07532_/A _07272_/Y _07811_/X _07927_/X VGND VGND VPWR VPWR _07936_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07859_ _07859_/A _07859_/B _07859_/C _07859_/D VGND VGND VPWR VPWR _07860_/C sky130_fd_sc_hd__and4_1
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _10510_/Q input39/X VGND VGND VPWR VPWR _09530_/A sky130_fd_sc_hd__and2_1
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10304_ _10508_/CLK _10304_/D repeater402/X VGND VGND VPWR VPWR _10304_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10235_ _10254_/CLK _10235_/D repeater406/X VGND VGND VPWR VPWR _10235_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10166_ _10244_/CLK _10166_/D repeater403/X VGND VGND VPWR VPWR _10166_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10097_ _10127_/CLK _10097_/D _07492_/B VGND VGND VPWR VPWR _10097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05210_ _05204_/Y _06429_/A _05208_/Y _05774_/A VGND VGND VPWR VPWR _05210_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06190_ _10004_/Q _07989_/B _06184_/A _10005_/Q VGND VGND VPWR VPWR _06190_/X sky130_fd_sc_hd__o31a_1
XFILLER_190_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05141_ _05141_/A _05141_/B _05141_/C _05140_/X VGND VGND VPWR VPWR _05366_/B sky130_fd_sc_hd__or4b_1
XFILLER_143_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05072_ _05167_/A _05205_/A VGND VGND VPWR VPWR _05960_/B sky130_fd_sc_hd__or2_1
X_08900_ _08900_/A _09277_/A VGND VGND VPWR VPWR _09390_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09880_ _10409_/CLK _09880_/D repeater407/X VGND VGND VPWR VPWR _09880_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08831_ _08836_/A _08831_/B VGND VGND VPWR VPWR _09286_/A sky130_fd_sc_hd__nor2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05974_ _10120_/Q _05969_/X _09579_/X _05971_/X VGND VGND VPWR VPWR _10120_/D sky130_fd_sc_hd__a22o_1
X_08762_ _08997_/A _09249_/A VGND VGND VPWR VPWR _09416_/A sky130_fd_sc_hd__or2_1
XFILLER_111_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _08693_/A _08749_/A VGND VGND VPWR VPWR _08693_/X sky130_fd_sc_hd__or2_1
X_07713_ _09513_/A _06232_/X _09455_/A _07533_/A _07712_/X VGND VGND VPWR VPWR _07716_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04925_ _05318_/A VGND VGND VPWR VPWR _05346_/A sky130_fd_sc_hd__buf_4
Xrepeater399 hold46/A VGND VGND VPWR VPWR _09661_/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07644_ _07638_/Y _07639_/X _07640_/Y _07641_/X _07643_/X VGND VGND VPWR VPWR _07650_/C
+ sky130_fd_sc_hd__o221a_1
X_04856_ _10505_/Q _04851_/X _09552_/X _04852_/X VGND VGND VPWR VPWR _10505_/D sky130_fd_sc_hd__o22a_1
XFILLER_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07575_ _07608_/A _07575_/B VGND VGND VPWR VPWR _07783_/A sky130_fd_sc_hd__or2_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09314_ _08457_/X _08461_/X _09372_/C _08548_/A _09039_/X VGND VGND VPWR VPWR _09315_/D
+ sky130_fd_sc_hd__o221ai_1
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06526_ _09834_/Q _06518_/A _09661_/A1 _06519_/A VGND VGND VPWR VPWR _09834_/D sky130_fd_sc_hd__a22o_1
X_06457_ _08402_/A _08402_/B _08402_/C _08402_/D VGND VGND VPWR VPWR _06458_/C sky130_fd_sc_hd__or4_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09245_ _09245_/A VGND VGND VPWR VPWR _09245_/Y sky130_fd_sc_hd__inv_2
X_05408_ hold45/A _05396_/X hold50/A _05398_/X VGND VGND VPWR VPWR _10415_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09176_ _09176_/A _09342_/A VGND VGND VPWR VPWR _09178_/B sky130_fd_sc_hd__or2_1
X_06388_ _06386_/X _09591_/X _09650_/X _09908_/Q VGND VGND VPWR VPWR _09908_/D sky130_fd_sc_hd__o22a_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ _09475_/A _08074_/X _09511_/A _08075_/X _08126_/X VGND VGND VPWR VPWR _08134_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05339_ _10386_/Q VGND VGND VPWR VPWR _05339_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08058_ _08177_/A VGND VGND VPWR VPWR _08058_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07009_ _10223_/Q VGND VGND VPWR VPWR _07009_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_163_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10020_ _10023_/CLK _10020_/D _05034_/A VGND VGND VPWR VPWR _10020_/Q sky130_fd_sc_hd__dfrtp_2
Xinput136 wb_adr_i[13] VGND VGND VPWR VPWR _08402_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput125 trap VGND VGND VPWR VPWR _05179_/A sky130_fd_sc_hd__buf_6
Xinput114 sram_ro_data[29] VGND VGND VPWR VPWR input114/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput103 sram_ro_data[19] VGND VGND VPWR VPWR input103/X sky130_fd_sc_hd__buf_2
Xinput169 wb_dat_i[13] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_adr_i[23] VGND VGND VPWR VPWR _08412_/A sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_adr_i[4] VGND VGND VPWR VPWR _08561_/B sky130_fd_sc_hd__buf_2
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_csclk clkbuf_leaf_2_csclk/A VGND VGND VPWR VPWR _10369_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10218_ _10491_/CLK _10218_/D repeater402/X VGND VGND VPWR VPWR _10218_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10149_ _10257_/CLK _10149_/D repeater407/X VGND VGND VPWR VPWR _10149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05690_ _05691_/A VGND VGND VPWR VPWR _05690_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07360_ _07358_/Y _05865_/B _07359_/Y _05927_/A VGND VGND VPWR VPWR _07360_/X sky130_fd_sc_hd__o22a_1
X_06311_ _09955_/Q _06305_/X _09574_/X _06306_/Y VGND VGND VPWR VPWR _09955_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09030_ _09030_/A VGND VGND VPWR VPWR _09176_/A sky130_fd_sc_hd__inv_2
X_07291_ _06763_/A _07290_/X _09760_/Q _06764_/A VGND VGND VPWR VPWR _09760_/D sky130_fd_sc_hd__o22a_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06242_ _06184_/A _07592_/A _07551_/B _06177_/A _06241_/X VGND VGND VPWR VPWR _09990_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_156_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06173_ _10008_/Q _06168_/X _06684_/B1 _06169_/Y VGND VGND VPWR VPWR _10008_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05124_ _05124_/A VGND VGND VPWR VPWR _06633_/A sky130_fd_sc_hd__inv_2
X_09932_ _10119_/CLK _09932_/D repeater402/X VGND VGND VPWR VPWR _09932_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05055_ _10425_/Q _05040_/X _09643_/X _05042_/X VGND VGND VPWR VPWR _10425_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09863_ _10157_/CLK _09863_/D repeater406/X VGND VGND VPWR VPWR _09863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08814_/A _08814_/B VGND VGND VPWR VPWR _09105_/B sky130_fd_sc_hd__or2_4
X_09794_ _10119_/CLK _09794_/D repeater403/X VGND VGND VPWR VPWR _09794_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08745_/A _09245_/A VGND VGND VPWR VPWR _08751_/A sky130_fd_sc_hd__nand2_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05957_ _10130_/Q _05953_/X _09660_/A1 _05954_/Y VGND VGND VPWR VPWR _10130_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05888_ _10173_/Q _05884_/X _09580_/X _05886_/X VGND VGND VPWR VPWR _10173_/D sky130_fd_sc_hd__a22o_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08809_/B _08676_/B VGND VGND VPWR VPWR _08823_/A sky130_fd_sc_hd__or2_1
XFILLER_81_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04908_ _10484_/Q _04902_/X _09658_/A1 _04904_/X VGND VGND VPWR VPWR _10484_/D sky130_fd_sc_hd__a22o_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07627_/A VGND VGND VPWR VPWR _07627_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04839_ _09678_/X _04822_/Y _06684_/B1 _10509_/Q _04827_/X VGND VGND VPWR VPWR _10509_/D
+ sky130_fd_sc_hd__a32o_1
X_07558_ _07558_/A VGND VGND VPWR VPWR _07585_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_06509_ _09846_/Q _06504_/X _09579_/X _06506_/X VGND VGND VPWR VPWR _09846_/D sky130_fd_sc_hd__a22o_1
XFILLER_158_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07489_ _07489_/A _07489_/B VGND VGND VPWR VPWR _07489_/X sky130_fd_sc_hd__or2_1
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09228_ _09180_/Y _09225_/Y _09237_/A _09152_/B VGND VGND VPWR VPWR _09324_/B sky130_fd_sc_hd__a31o_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09159_ _09159_/A _09395_/A VGND VGND VPWR VPWR _09161_/C sky130_fd_sc_hd__or2_1
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10003_ _10006_/CLK _10003_/D repeater409/X VGND VGND VPWR VPWR _10003_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06860_ _06858_/Y _06708_/B _06859_/Y _05749_/B VGND VGND VPWR VPWR _06860_/X sky130_fd_sc_hd__o22a_1
X_05811_ _05811_/A VGND VGND VPWR VPWR _05811_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06791_ _09860_/Q VGND VGND VPWR VPWR _06791_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08530_ _08537_/C _09236_/A _09233_/A _08530_/D VGND VGND VPWR VPWR _08582_/B sky130_fd_sc_hd__or4_4
X_05742_ _05742_/A VGND VGND VPWR VPWR _05742_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08461_ _09046_/A VGND VGND VPWR VPWR _08461_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05673_ _06568_/A VGND VGND VPWR VPWR _05674_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07412_ _10371_/Q VGND VGND VPWR VPWR _07412_/Y sky130_fd_sc_hd__inv_2
X_08392_ _08938_/A VGND VGND VPWR VPWR _08972_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07343_ _09793_/Q VGND VGND VPWR VPWR _07343_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07274_ _07269_/Y _06304_/B _07270_/Y _06290_/A _07273_/X VGND VGND VPWR VPWR _07287_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_191_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09013_ _09010_/X _09206_/A _09046_/B _09001_/A VGND VGND VPWR VPWR _09013_/X sky130_fd_sc_hd__o22a_1
X_06225_ _07528_/A _06237_/A VGND VGND VPWR VPWR _07558_/A sky130_fd_sc_hd__or2_1
XFILLER_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06156_ _06156_/A VGND VGND VPWR VPWR _06157_/A sky130_fd_sc_hd__inv_2
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06087_ _06087_/A _06087_/B VGND VGND VPWR VPWR _06089_/A sky130_fd_sc_hd__or2_1
X_05107_ input36/X _06693_/A input123/X _05101_/X _05106_/Y VGND VGND VPWR VPWR _05108_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09915_ _10397_/CLK _09915_/D repeater407/X VGND VGND VPWR VPWR _09915_/Q sky130_fd_sc_hd__dfrtp_1
X_05038_ _09772_/Q VGND VGND VPWR VPWR _05395_/A sky130_fd_sc_hd__inv_2
X_09846_ _10350_/CLK _09846_/D repeater404/X VGND VGND VPWR VPWR _09846_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _06987_/Y _05808_/B _07738_/A _06267_/B VGND VGND VPWR VPWR _06989_/X sky130_fd_sc_hd__o22a_1
X_09777_ _10023_/CLK _09777_/D _05034_/A VGND VGND VPWR VPWR _09777_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _08743_/A _09263_/A _08727_/Y VGND VGND VPWR VPWR _08728_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08845_/A VGND VGND VPWR VPWR _08849_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10483_ _10483_/CLK _10483_/D _05034_/A VGND VGND VPWR VPWR _10483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06010_ _06010_/A VGND VGND VPWR VPWR _06011_/B sky130_fd_sc_hd__clkbuf_4
Xoutput226 _09506_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput215 _09486_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_173_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput204 _10482_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_2
Xoutput259 _09721_/Z VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput237 _09570_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput248 _09711_/Z VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07961_ _07961_/A _07961_/B _07961_/C _07961_/D VGND VGND VPWR VPWR _07962_/C sky130_fd_sc_hd__and4_1
XFILLER_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06912_ input39/X _09699_/S _10436_/Q _05121_/Y VGND VGND VPWR VPWR _06912_/X sky130_fd_sc_hd__a22o_1
X_09700_ _08051_/X _07506_/Y _09700_/S VGND VGND VPWR VPWR _09700_/X sky130_fd_sc_hd__mux2_1
X_07892_ _07368_/Y _07787_/X _07401_/Y _07788_/X _07891_/X VGND VGND VPWR VPWR _07901_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09631_ _09630_/X _09889_/Q _09776_/Q VGND VGND VPWR VPWR _09631_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06843_ input31/X _05129_/X _06837_/X _06840_/X _06842_/X VGND VGND VPWR VPWR _06905_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09562_ _09561_/X input74/X _10297_/Q VGND VGND VPWR VPWR _09562_/X sky130_fd_sc_hd__mux2_1
X_06774_ input59/X _05114_/X _10061_/Q _05162_/X _06773_/X VGND VGND VPWR VPWR _06775_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08513_ _09085_/D _09085_/B _09102_/C _08624_/A VGND VGND VPWR VPWR _08575_/A sky130_fd_sc_hd__or4_4
X_05725_ _10267_/Q _05717_/A _09585_/X _05718_/A VGND VGND VPWR VPWR _10267_/D sky130_fd_sc_hd__o22a_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09493_ _09493_/A VGND VGND VPWR VPWR _09494_/A sky130_fd_sc_hd__clkbuf_1
X_05656_ _10307_/Q _05653_/X _09581_/X _05655_/X VGND VGND VPWR VPWR _10307_/D sky130_fd_sc_hd__a22o_1
X_08444_ _08703_/A VGND VGND VPWR VPWR _08710_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08375_ _09102_/C _08494_/A VGND VGND VPWR VPWR _08389_/A sky130_fd_sc_hd__or2_1
X_05587_ _10343_/Q _05578_/A _09659_/A1 _05579_/A VGND VGND VPWR VPWR _10343_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07326_ _10064_/Q VGND VGND VPWR VPWR _07326_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07257_ _09935_/Q VGND VGND VPWR VPWR _07257_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07188_ _10057_/Q VGND VGND VPWR VPWR _07188_/Y sky130_fd_sc_hd__inv_2
X_06208_ _06208_/A VGND VGND VPWR VPWR _06209_/A sky130_fd_sc_hd__inv_2
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06139_ _06139_/A VGND VGND VPWR VPWR _06150_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09829_ _10354_/CLK _09829_/D repeater406/X VGND VGND VPWR VPWR _09829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10466_ _10471_/CLK _10466_/D repeater409/X VGND VGND VPWR VPWR _10466_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _04811_/A1 sky130_fd_sc_hd__clkbuf_2
X_10397_ _10397_/CLK _10397_/D _05447_/X VGND VGND VPWR VPWR _10397_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05510_ _05518_/A VGND VGND VPWR VPWR _05511_/A sky130_fd_sc_hd__clkbuf_1
X_06490_ _09856_/Q _06483_/A _09660_/A1 _06484_/A VGND VGND VPWR VPWR _09856_/D sky130_fd_sc_hd__a22o_1
X_05441_ _10402_/Q _05435_/X _09545_/A1 _05437_/X VGND VGND VPWR VPWR _10402_/D sky130_fd_sc_hd__a22o_1
X_08160_ _06898_/Y _08069_/X _06894_/Y _08070_/X VGND VGND VPWR VPWR _08160_/X sky130_fd_sc_hd__o22a_1
X_07111_ _09831_/Q VGND VGND VPWR VPWR _07111_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05372_ _09808_/Q VGND VGND VPWR VPWR _05429_/D sky130_fd_sc_hd__inv_2
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08091_ _07413_/Y _08086_/X _07389_/Y _08087_/X _08090_/X VGND VGND VPWR VPWR _08098_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07042_ input23/X _06704_/X _10136_/Q _06705_/Y _07041_/X VGND VGND VPWR VPWR _07047_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08993_ _08993_/A _08993_/B VGND VGND VPWR VPWR _08994_/B sky130_fd_sc_hd__and2_1
X_07944_ _07071_/Y _07792_/A _07059_/Y _07793_/A _07943_/X VGND VGND VPWR VPWR _07951_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07875_ _07875_/A _07875_/B _07875_/C _07875_/D VGND VGND VPWR VPWR _07886_/B sky130_fd_sc_hd__and4_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06826_ _06821_/Y _05928_/B _06822_/Y _06893_/B _06825_/X VGND VGND VPWR VPWR _06833_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09614_ _07672_/Y _10330_/Q _09682_/S VGND VGND VPWR VPWR _09614_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06757_ _06741_/Y _05434_/B _06744_/X _06750_/X _06756_/X VGND VGND VPWR VPWR _06757_/X
+ sky130_fd_sc_hd__o2111a_1
X_09545_ _10320_/Q _09545_/A1 _09679_/S VGND VGND VPWR VPWR _09545_/X sky130_fd_sc_hd__mux2_1
X_09476_ _09476_/A VGND VGND VPWR VPWR _09476_/X sky130_fd_sc_hd__clkbuf_1
X_05708_ _10277_/Q _05701_/A _09660_/X _05702_/A VGND VGND VPWR VPWR _10277_/D sky130_fd_sc_hd__o22a_1
X_06688_ _06688_/A VGND VGND VPWR VPWR _06688_/X sky130_fd_sc_hd__clkbuf_2
X_08427_ _08888_/A VGND VGND VPWR VPWR _08556_/D sky130_fd_sc_hd__clkbuf_2
X_05639_ _05639_/A VGND VGND VPWR VPWR _05641_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08358_ _09790_/Q input181/X _09789_/Q input195/X _08357_/X VGND VGND VPWR VPWR _08358_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08289_ _07266_/Y _08213_/X _07269_/Y _08214_/X VGND VGND VPWR VPWR _08289_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07309_ input104/X _06696_/A _10325_/Q _05156_/Y VGND VGND VPWR VPWR _07309_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10320_ _10405_/CLK _10320_/D hold41/X VGND VGND VPWR VPWR _10320_/Q sky130_fd_sc_hd__dfrtp_1
X_10251_ _10504_/CLK _10251_/D repeater403/X VGND VGND VPWR VPWR _10251_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10182_ _10257_/CLK _10182_/D repeater407/X VGND VGND VPWR VPWR _10182_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10449_ _10487_/CLK _10449_/D repeater409/X VGND VGND VPWR VPWR _10449_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05990_ _10108_/Q _05982_/A _06684_/B1 _05983_/A VGND VGND VPWR VPWR _10108_/D sky130_fd_sc_hd__a22o_1
X_04941_ _10476_/Q _04935_/X _09545_/A1 _04937_/X VGND VGND VPWR VPWR _10476_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04872_ _04873_/A VGND VGND VPWR VPWR _04872_/X sky130_fd_sc_hd__clkbuf_2
X_07660_ _07321_/Y _07658_/X _07298_/Y _07659_/X VGND VGND VPWR VPWR _07660_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06611_ _06614_/A VGND VGND VPWR VPWR _06612_/A sky130_fd_sc_hd__clkbuf_1
X_07591_ _07588_/Y _07639_/A _05102_/Y _07801_/A _07590_/X VGND VGND VPWR VPWR _07595_/C
+ sky130_fd_sc_hd__o221a_1
X_09330_ _09223_/A _08761_/A _09229_/A _09223_/A VGND VGND VPWR VPWR _09418_/B sky130_fd_sc_hd__o22ai_1
X_06542_ _09827_/Q _06539_/X _09581_/X _06541_/X VGND VGND VPWR VPWR _09827_/D sky130_fd_sc_hd__a22o_1
X_09261_ _09261_/A VGND VGND VPWR VPWR _09265_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06473_ _06474_/A VGND VGND VPWR VPWR _06473_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08212_ _08212_/A VGND VGND VPWR VPWR _08212_/X sky130_fd_sc_hd__buf_2
X_09192_ _08883_/B _09093_/A _08776_/B VGND VGND VPWR VPWR _09222_/C sky130_fd_sc_hd__o21ai_1
X_05424_ _10409_/Q _05420_/X _06683_/B1 _05421_/Y VGND VGND VPWR VPWR _10409_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05355_ _05355_/A _05355_/B VGND VGND VPWR VPWR _06312_/A sky130_fd_sc_hd__or2_2
X_08143_ _07016_/Y _08064_/X _08140_/X _08142_/X VGND VGND VPWR VPWR _08153_/C sky130_fd_sc_hd__o211a_1
XFILLER_174_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08074_ _08193_/A VGND VGND VPWR VPWR _08074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05286_ _05286_/A _05286_/B VGND VGND VPWR VPWR _05807_/A sky130_fd_sc_hd__or2_2
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07025_ _07023_/Y _06537_/A _07024_/Y _05821_/B VGND VGND VPWR VPWR _07025_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08976_ _09051_/A _09295_/C _09051_/B VGND VGND VPWR VPWR _08977_/A sky130_fd_sc_hd__or3b_2
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold25 hold25/A VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07927_ _07246_/Y _07812_/X _07182_/Y _07813_/X VGND VGND VPWR VPWR _07927_/X sky130_fd_sc_hd__o22a_1
X_07858_ _06746_/Y _07825_/X _07856_/Y _07827_/X _07857_/X VGND VGND VPWR VPWR _07859_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07789_ _07789_/A VGND VGND VPWR VPWR _07789_/X sky130_fd_sc_hd__buf_4
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06809_ _10363_/Q VGND VGND VPWR VPWR _06809_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09528_ _09528_/A VGND VGND VPWR VPWR _09528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09459_ _09459_/A VGND VGND VPWR VPWR _09460_/A sky130_fd_sc_hd__clkbuf_1
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10303_ _10508_/CLK _10303_/D repeater402/X VGND VGND VPWR VPWR _10303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10234_ _10254_/CLK _10234_/D repeater406/X VGND VGND VPWR VPWR _10234_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10165_ _10244_/CLK _10165_/D repeater403/X VGND VGND VPWR VPWR _10165_/Q sky130_fd_sc_hd__dfrtp_1
X_10096_ _10289_/CLK _10096_/D repeater402/X VGND VGND VPWR VPWR _10096_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05140_ _05133_/Y _04827_/B _05134_/Y _05968_/B _05139_/X VGND VGND VPWR VPWR _05140_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05071_ _05164_/B VGND VGND VPWR VPWR _05167_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08830_ _08830_/A _09064_/A _09354_/A _09065_/A VGND VGND VPWR VPWR _08834_/A sky130_fd_sc_hd__or4_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05973_ _10121_/Q _05969_/X _09580_/X _05971_/X VGND VGND VPWR VPWR _10121_/D sky130_fd_sc_hd__a22o_1
X_08761_ _08761_/A _08766_/B VGND VGND VPWR VPWR _09249_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08692_ _08895_/A _08913_/B _08692_/C VGND VGND VPWR VPWR _08749_/A sky130_fd_sc_hd__or3_4
X_04924_ _09683_/X _04923_/A _10481_/Q _04923_/Y VGND VGND VPWR VPWR _10481_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07712_ _09481_/A _07770_/B VGND VGND VPWR VPWR _07712_/X sky130_fd_sc_hd__or2_1
X_04855_ _10506_/Q _04851_/X _09553_/X _04852_/X VGND VGND VPWR VPWR _10506_/D sky130_fd_sc_hd__o22a_1
X_07643_ _07400_/Y _07568_/B _07363_/Y _07642_/X VGND VGND VPWR VPWR _07643_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09313_ _09313_/A _09408_/A _09374_/C _09313_/D VGND VGND VPWR VPWR _09315_/B sky130_fd_sc_hd__or4_1
X_07574_ _07608_/A _07574_/B VGND VGND VPWR VPWR _07782_/A sky130_fd_sc_hd__or2_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06525_ _09835_/Q _06518_/A _09660_/A1 _06519_/A VGND VGND VPWR VPWR _09835_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06456_ _08401_/A _08401_/B _08399_/A _08399_/B VGND VGND VPWR VPWR _06466_/B sky130_fd_sc_hd__or4_1
XFILLER_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09244_ _09244_/A _09380_/C _09327_/D _09411_/A VGND VGND VPWR VPWR _09250_/A sky130_fd_sc_hd__or4_2
XFILLER_178_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05407_ _05407_/A VGND VGND VPWR VPWR _05407_/X sky130_fd_sc_hd__clkbuf_1
X_09175_ _09175_/A VGND VGND VPWR VPWR _09342_/A sky130_fd_sc_hd__inv_2
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08126_ _09491_/A _08076_/X _09489_/A _08077_/X VGND VGND VPWR VPWR _08126_/X sky130_fd_sc_hd__o22a_1
X_06387_ _06386_/X _09593_/X _09650_/X _09909_/Q VGND VGND VPWR VPWR _09909_/D sky130_fd_sc_hd__o22a_1
XFILLER_147_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05338_ _05338_/A _05338_/B VGND VGND VPWR VPWR _06166_/A sky130_fd_sc_hd__or2_2
X_05269_ _05265_/Y _06095_/A _05267_/Y _05909_/A VGND VGND VPWR VPWR _05269_/X sky130_fd_sc_hd__o22a_1
X_08057_ _07408_/Y _08052_/X _07384_/Y _08053_/X _08056_/X VGND VGND VPWR VPWR _08099_/A
+ sky130_fd_sc_hd__o221a_1
X_07008_ _07003_/Y _05838_/A _07004_/Y _06351_/B _07007_/X VGND VGND VPWR VPWR _07027_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput126 uart_enabled VGND VGND VPWR VPWR _09521_/B sky130_fd_sc_hd__buf_4
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput104 sram_ro_data[1] VGND VGND VPWR VPWR input104/X sky130_fd_sc_hd__clkbuf_2
Xinput115 sram_ro_data[2] VGND VGND VPWR VPWR input115/X sky130_fd_sc_hd__clkbuf_2
Xinput148 wb_adr_i[24] VGND VGND VPWR VPWR _06455_/C sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_adr_i[14] VGND VGND VPWR VPWR _08401_/B sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_adr_i[5] VGND VGND VPWR VPWR _09233_/A sky130_fd_sc_hd__buf_6
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08959_ _09046_/A _08959_/B VGND VGND VPWR VPWR _09075_/B sky130_fd_sc_hd__nor2_2
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10217_ _10290_/CLK _10217_/D repeater402/X VGND VGND VPWR VPWR _10217_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10148_ _10491_/CLK _10148_/D repeater403/X VGND VGND VPWR VPWR _10148_/Q sky130_fd_sc_hd__dfrtp_1
X_10079_ _10411_/CLK _10079_/D repeater407/X VGND VGND VPWR VPWR _10079_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06310_ _09956_/Q _06305_/X hold46/X _06306_/Y VGND VGND VPWR VPWR _09956_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07290_ _07290_/A VGND VGND VPWR VPWR _07290_/X sky130_fd_sc_hd__clkbuf_8
X_06241_ _09989_/Q _09988_/Q _09777_/Q _09990_/Q VGND VGND VPWR VPWR _06241_/X sky130_fd_sc_hd__a31o_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06172_ _10009_/Q _06168_/X _06683_/B1 _06169_/Y VGND VGND VPWR VPWR _10009_/D sky130_fd_sc_hd__a22o_1
X_05123_ _10430_/Q _05030_/Y input131/X _05118_/Y _05122_/X VGND VGND VPWR VPWR _05141_/B
+ sky130_fd_sc_hd__a221o_1
X_09931_ _10119_/CLK _09931_/D repeater402/X VGND VGND VPWR VPWR _09931_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05054_ _05054_/A VGND VGND VPWR VPWR _05054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09862_ _10157_/CLK _09862_/D repeater406/X VGND VGND VPWR VPWR _09862_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _10157_/CLK _09793_/D repeater406/X VGND VGND VPWR VPWR _09793_/Q sky130_fd_sc_hd__dfrtp_1
X_08813_ _08813_/A VGND VGND VPWR VPWR _09105_/A sky130_fd_sc_hd__buf_2
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05956_ _10131_/Q _05953_/X _09577_/X _05954_/Y VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__a22o_1
X_08744_ _09093_/A _08860_/A VGND VGND VPWR VPWR _09245_/A sky130_fd_sc_hd__or2_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04907_ _10485_/Q _04902_/X _06683_/B1 _04904_/X VGND VGND VPWR VPWR _10485_/D sky130_fd_sc_hd__a22o_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08675_/A _08675_/B VGND VGND VPWR VPWR _08809_/B sky130_fd_sc_hd__nand2_4
X_05887_ _10174_/Q _05884_/X _09581_/X _05886_/X VGND VGND VPWR VPWR _10174_/D sky130_fd_sc_hd__a22o_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _07396_/Y _07618_/X _07395_/Y _07619_/X _07625_/X VGND VGND VPWR VPWR _07672_/A
+ sky130_fd_sc_hd__o221a_1
X_04838_ _09678_/X _04835_/Y _06684_/B1 _10510_/Q _04836_/X VGND VGND VPWR VPWR _10510_/D
+ sky130_fd_sc_hd__a32o_1
X_07557_ _07565_/A _07596_/B VGND VGND VPWR VPWR _07589_/A sky130_fd_sc_hd__or2_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06508_ _09847_/Q _06504_/X _09580_/X _06506_/X VGND VGND VPWR VPWR _09847_/D sky130_fd_sc_hd__a22o_1
XFILLER_158_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07488_ _07487_/Y _07468_/Y _05430_/Y _09773_/Q _07489_/A VGND VGND VPWR VPWR _09773_/D
+ sky130_fd_sc_hd__a32o_1
X_06439_ _06481_/A _06439_/B VGND VGND VPWR VPWR _06441_/A sky130_fd_sc_hd__or2_2
X_09227_ _09224_/Y _09225_/Y _09237_/A _09161_/C VGND VGND VPWR VPWR _09319_/A sky130_fd_sc_hd__a31o_1
XFILLER_154_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09158_ _09158_/A VGND VGND VPWR VPWR _09395_/A sky130_fd_sc_hd__inv_2
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09089_ _09275_/A _09222_/A VGND VGND VPWR VPWR _09363_/B sky130_fd_sc_hd__or2_1
XFILLER_135_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08109_ _07257_/Y _08074_/X _07245_/Y _08075_/X _08108_/X VGND VGND VPWR VPWR _08116_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10002_ _10006_/CLK _10002_/D repeater409/X VGND VGND VPWR VPWR _10002_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05810_ _05810_/A VGND VGND VPWR VPWR _05811_/A sky130_fd_sc_hd__inv_2
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06790_ _09874_/Q VGND VGND VPWR VPWR _06790_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05741_ _05742_/A VGND VGND VPWR VPWR _05741_/X sky130_fd_sc_hd__clkbuf_2
X_08460_ _08951_/A VGND VGND VPWR VPWR _09046_/A sky130_fd_sc_hd__clkbuf_4
X_05672_ _09770_/Q _05671_/B _10419_/Q _10298_/Q _05671_/Y VGND VGND VPWR VPWR _10298_/D
+ sky130_fd_sc_hd__a32o_1
X_08391_ _08916_/A VGND VGND VPWR VPWR _08938_/A sky130_fd_sc_hd__clkbuf_4
X_07411_ _07406_/Y _05575_/A _07407_/Y _06359_/A _07410_/X VGND VGND VPWR VPWR _07418_/C
+ sky130_fd_sc_hd__o221a_1
X_07342_ _07337_/Y _06122_/B _07338_/Y _04886_/B _07341_/X VGND VGND VPWR VPWR _07349_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07273_ _07271_/Y _05830_/B _07272_/Y _06167_/B VGND VGND VPWR VPWR _07273_/X sky130_fd_sc_hd__o22a_2
XFILLER_136_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ _09012_/A VGND VGND VPWR VPWR _09046_/B sky130_fd_sc_hd__buf_2
X_06224_ _09990_/Q VGND VGND VPWR VPWR _06237_/A sky130_fd_sc_hd__inv_2
X_06155_ _06156_/A VGND VGND VPWR VPWR _06155_/X sky130_fd_sc_hd__clkbuf_2
X_05106_ _05102_/Y _06705_/A _05105_/X VGND VGND VPWR VPWR _05106_/Y sky130_fd_sc_hd__o21ai_1
X_06086_ _10050_/Q _06080_/X _09536_/A3 _06081_/Y VGND VGND VPWR VPWR _10050_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09914_ _10397_/CLK _09914_/D repeater407/X VGND VGND VPWR VPWR _09914_/Q sky130_fd_sc_hd__dfrtp_1
X_05037_ _09811_/Q VGND VGND VPWR VPWR _05713_/A sky130_fd_sc_hd__clkinv_4
X_09845_ _10350_/CLK _09845_/D repeater404/X VGND VGND VPWR VPWR _09845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10336_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06988_ _09978_/Q VGND VGND VPWR VPWR _07738_/A sky130_fd_sc_hd__inv_2
X_09776_ _10023_/CLK _09776_/D _05034_/A VGND VGND VPWR VPWR _09776_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05939_ _10141_/Q _05930_/A _09659_/A1 _05931_/A VGND VGND VPWR VPWR _10141_/D sky130_fd_sc_hd__a22o_1
X_08727_ _08727_/A _09397_/A VGND VGND VPWR VPWR _08727_/Y sky130_fd_sc_hd__nor2_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08676_/B _08672_/B VGND VGND VPWR VPWR _08845_/A sky130_fd_sc_hd__or2_1
XFILLER_54_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07609_ _10055_/Q VGND VGND VPWR VPWR _07609_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08589_ _08490_/A _08999_/B _08527_/Y _08588_/Y VGND VGND VPWR VPWR _08590_/B sky130_fd_sc_hd__a31o_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10482_ _10482_/CLK _10482_/D repeater405/X VGND VGND VPWR VPWR _10482_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _09572_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput216 _09488_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xoutput205 _09528_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_2
Xoutput227 _09508_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_2
Xoutput249 _09712_/Z VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput238 _09456_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07960_ _07080_/Y _07825_/A _07054_/Y _07827_/A _07959_/X VGND VGND VPWR VPWR _07961_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06911_ _10447_/Q _06688_/X _10033_/Q _05080_/X _06910_/X VGND VGND VPWR VPWR _06911_/X
+ sky130_fd_sc_hd__a221o_1
X_07891_ _07370_/Y _07749_/X _07353_/Y _07789_/X VGND VGND VPWR VPWR _07891_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09630_ _07912_/Y _10325_/Q _09682_/S VGND VGND VPWR VPWR _09630_/X sky130_fd_sc_hd__mux2_1
X_06842_ input57/X _05114_/X input97/X _05101_/X _06841_/X VGND VGND VPWR VPWR _06842_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_82_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06773_ _10139_/Q _06705_/Y input32/X _05129_/X VGND VGND VPWR VPWR _06773_/X sky130_fd_sc_hd__a22o_1
X_09561_ _09560_/X input38/X _10342_/Q VGND VGND VPWR VPWR _09561_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05724_ _10268_/Q _05717_/A _09586_/X _05718_/A VGND VGND VPWR VPWR _10268_/D sky130_fd_sc_hd__o22a_1
X_08512_ _08512_/A _08752_/A VGND VGND VPWR VPWR _08596_/A sky130_fd_sc_hd__or2_1
X_09492_ _09492_/A VGND VGND VPWR VPWR _09492_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05655_ _05655_/A VGND VGND VPWR VPWR _05655_/X sky130_fd_sc_hd__clkbuf_2
X_08443_ _09102_/B _08783_/A VGND VGND VPWR VPWR _08703_/A sky130_fd_sc_hd__or2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08374_ _08631_/C VGND VGND VPWR VPWR _08472_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05586_ _10344_/Q _05578_/A _09661_/A1 _05579_/A VGND VGND VPWR VPWR _10344_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07325_ _09934_/Q VGND VGND VPWR VPWR _07325_/Y sky130_fd_sc_hd__clkinv_2
X_07256_ _10091_/Q VGND VGND VPWR VPWR _07256_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06207_ _06208_/A VGND VGND VPWR VPWR _06207_/X sky130_fd_sc_hd__clkbuf_2
X_07187_ _07182_/Y _05419_/B _07183_/Y _05794_/B _07186_/X VGND VGND VPWR VPWR _07187_/X
+ sky130_fd_sc_hd__o221a_1
X_06138_ _10023_/Q VGND VGND VPWR VPWR _06140_/A sky130_fd_sc_hd__inv_2
X_06069_ _06069_/A VGND VGND VPWR VPWR _06069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09828_ _10354_/CLK _09828_/D repeater406/X VGND VGND VPWR VPWR _09828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09759_ _09919_/CLK _09759_/D VGND VGND VPWR VPWR _09759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10465_ _10471_/CLK _10465_/D repeater409/X VGND VGND VPWR VPWR _10465_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10396_ _10397_/CLK _10396_/D _05454_/X VGND VGND VPWR VPWR _10396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05440_ _10403_/Q _05435_/X _09579_/X _05437_/X VGND VGND VPWR VPWR _10403_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05371_ _09809_/Q VGND VGND VPWR VPWR _05429_/A sky130_fd_sc_hd__inv_2
X_07110_ _10209_/Q VGND VGND VPWR VPWR _07110_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08090_ _07381_/Y _08088_/X _07396_/Y _08089_/X VGND VGND VPWR VPWR _08090_/X sky130_fd_sc_hd__o22a_1
X_07041_ input112/X _05112_/A _10454_/Q _05089_/X VGND VGND VPWR VPWR _07041_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08992_ _08992_/A _09362_/C VGND VGND VPWR VPWR _08993_/B sky130_fd_sc_hd__or2_1
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07943_ _07074_/Y _07794_/A _07060_/Y _07795_/A VGND VGND VPWR VPWR _07943_/X sky130_fd_sc_hd__o22a_1
X_07874_ _05204_/Y _07805_/X _07872_/Y _07758_/X _07873_/X VGND VGND VPWR VPWR _07875_/D
+ sky130_fd_sc_hd__o221a_1
X_06825_ _06823_/Y _05968_/B _06824_/Y _05896_/B VGND VGND VPWR VPWR _06825_/X sky130_fd_sc_hd__o22a_1
X_09613_ _09612_/X _09918_/Q _09776_/Q VGND VGND VPWR VPWR _09613_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09544_ _10308_/Q _09659_/A1 _09699_/S VGND VGND VPWR VPWR _09544_/X sky130_fd_sc_hd__mux2_1
X_06756_ _06751_/Y _05928_/B _06752_/Y _05883_/B _06755_/X VGND VGND VPWR VPWR _06756_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_70_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09475_ _09475_/A VGND VGND VPWR VPWR _09476_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05707_ _10278_/Q _05701_/X _09658_/X _05702_/X VGND VGND VPWR VPWR _10278_/D sky130_fd_sc_hd__o22a_1
X_06687_ _10036_/Q _05080_/X input108/X _05153_/X _06686_/X VGND VGND VPWR VPWR _06701_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08426_ _08426_/A VGND VGND VPWR VPWR _08888_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05638_ _05651_/A _05651_/B _05638_/C VGND VGND VPWR VPWR _05639_/A sky130_fd_sc_hd__or3_4
X_08357_ _09788_/Q _08357_/B VGND VGND VPWR VPWR _08357_/X sky130_fd_sc_hd__and2_1
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05569_ _05569_/A VGND VGND VPWR VPWR _05569_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08288_ _07278_/Y _08205_/X _07215_/Y _08206_/X _08287_/X VGND VGND VPWR VPWR _08291_/C
+ sky130_fd_sc_hd__o221a_1
X_07308_ _10473_/Q _06933_/B _09791_/Q _06633_/X _07307_/Y VGND VGND VPWR VPWR _07324_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07239_ _10353_/Q VGND VGND VPWR VPWR _07239_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_137_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10250_ _10504_/CLK _10250_/D repeater403/X VGND VGND VPWR VPWR _10250_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_34_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _10369_/CLK _10181_/D repeater407/X VGND VGND VPWR VPWR _10181_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_49_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10448_ _10487_/CLK _10448_/D _05034_/A VGND VGND VPWR VPWR _10448_/Q sky130_fd_sc_hd__dfstp_2
X_10379_ _10382_/CLK _10379_/D _05519_/X VGND VGND VPWR VPWR _10379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04940_ _10477_/Q _04935_/X _09579_/X _04937_/X VGND VGND VPWR VPWR _10477_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04871_ _05541_/A _04871_/B VGND VGND VPWR VPWR _04873_/A sky130_fd_sc_hd__or2_1
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07590_ _05271_/Y _07512_/A _05274_/Y _07642_/A VGND VGND VPWR VPWR _07590_/X sky130_fd_sc_hd__o22a_2
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06610_ _09805_/Q _06604_/X _09651_/X _06606_/X VGND VGND VPWR VPWR _09805_/D sky130_fd_sc_hd__a22o_1
X_06541_ _06541_/A VGND VGND VPWR VPWR _06541_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06472_ _06472_/A _06472_/B VGND VGND VPWR VPWR _06474_/A sky130_fd_sc_hd__or2_2
X_09260_ _09260_/A _09261_/A VGND VGND VPWR VPWR _09339_/D sky130_fd_sc_hd__nor2_1
X_05423_ _10410_/Q _05420_/X _09577_/X _05421_/Y VGND VGND VPWR VPWR _10410_/D sky130_fd_sc_hd__a22o_1
X_08211_ _08211_/A VGND VGND VPWR VPWR _08211_/X sky130_fd_sc_hd__buf_2
X_09191_ _09191_/A _09317_/A VGND VGND VPWR VPWR _09193_/A sky130_fd_sc_hd__or2_1
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05354_ _09947_/Q VGND VGND VPWR VPWR _05354_/Y sky130_fd_sc_hd__clkinv_2
X_08142_ _06970_/Y _08067_/X _06961_/Y _08068_/X _08141_/X VGND VGND VPWR VPWR _08142_/X
+ sky130_fd_sc_hd__o221a_1
X_05285_ _10211_/Q VGND VGND VPWR VPWR _05285_/Y sky130_fd_sc_hd__clkinv_4
X_08073_ _07415_/Y _08064_/X _08066_/X _08072_/X VGND VGND VPWR VPWR _08099_/C sky130_fd_sc_hd__o211a_1
XFILLER_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07024_ _10210_/Q VGND VGND VPWR VPWR _07024_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08975_ _09233_/A _08483_/D _08849_/A _08695_/A _08884_/Y VGND VGND VPWR VPWR _09051_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07926_ _07926_/A _07926_/B _07926_/C _07926_/D VGND VGND VPWR VPWR _07937_/B sky130_fd_sc_hd__and4_1
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold15 hold15/A VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07857_ _06729_/Y _07828_/X _06737_/Y _07829_/X VGND VGND VPWR VPWR _07857_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07788_ _07788_/A VGND VGND VPWR VPWR _07788_/X sky130_fd_sc_hd__buf_2
XFILLER_71_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06808_ _10376_/Q VGND VGND VPWR VPWR _06808_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06739_ _06734_/Y _06538_/B _06735_/Y _06360_/B _06738_/X VGND VGND VPWR VPWR _06740_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09527_ _10511_/Q input70/X VGND VGND VPWR VPWR _09528_/A sky130_fd_sc_hd__and2_2
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09458_ _09458_/A VGND VGND VPWR VPWR _09458_/X sky130_fd_sc_hd__clkbuf_1
X_08409_ _08379_/B _08408_/Y _08492_/B _08408_/A VGND VGND VPWR VPWR _08564_/A sky130_fd_sc_hd__o22a_1
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09389_ _09389_/A _09389_/B _09389_/C _09389_/D VGND VGND VPWR VPWR _09443_/D sky130_fd_sc_hd__or4_2
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10302_ _10508_/CLK hold43/X repeater404/X VGND VGND VPWR VPWR _10302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10233_ _10254_/CLK _10233_/D repeater406/X VGND VGND VPWR VPWR _10233_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10164_ _10238_/CLK _10164_/D repeater403/X VGND VGND VPWR VPWR _10164_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10095_ _10289_/CLK _10095_/D repeater402/X VGND VGND VPWR VPWR _10095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05070_ _06002_/B VGND VGND VPWR VPWR _05070_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05972_ _10122_/Q _05969_/X _09581_/X _05971_/X VGND VGND VPWR VPWR _10122_/D sky130_fd_sc_hd__a22o_1
X_08760_ _08897_/A _08766_/A VGND VGND VPWR VPWR _08997_/A sky130_fd_sc_hd__nor2_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04923_ _04923_/A VGND VGND VPWR VPWR _04923_/Y sky130_fd_sc_hd__inv_2
X_08691_ _08686_/Y _09278_/B _08753_/C VGND VGND VPWR VPWR _08700_/A sky130_fd_sc_hd__o21a_1
XFILLER_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07711_ _09459_/A _07656_/X _09487_/A _07657_/X _07710_/X VGND VGND VPWR VPWR _07716_/B
+ sky130_fd_sc_hd__o221a_1
X_04854_ _10507_/Q _04851_/X _09583_/X _04852_/X VGND VGND VPWR VPWR _10507_/D sky130_fd_sc_hd__o22a_1
X_07642_ _07642_/A VGND VGND VPWR VPWR _07642_/X sky130_fd_sc_hd__buf_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09312_ _09312_/A _09312_/B VGND VGND VPWR VPWR _09374_/C sky130_fd_sc_hd__or2_1
X_07573_ _07573_/A VGND VGND VPWR VPWR _07781_/A sky130_fd_sc_hd__buf_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06524_ _09836_/Q _06517_/X _09658_/A1 _06519_/X VGND VGND VPWR VPWR _09836_/D sky130_fd_sc_hd__a22o_1
X_06455_ _08399_/C _08399_/D _06455_/C input149/X VGND VGND VPWR VPWR _06466_/A sky130_fd_sc_hd__or4b_1
XFILLER_166_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ _09179_/Y _09231_/Y _09237_/X _09178_/B VGND VGND VPWR VPWR _09411_/A sky130_fd_sc_hd__a31o_1
XFILLER_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05406_ _05406_/A VGND VGND VPWR VPWR _05407_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09174_ _09174_/A _09327_/C VGND VGND VPWR VPWR _09178_/A sky130_fd_sc_hd__or2_1
X_06386_ _06417_/A VGND VGND VPWR VPWR _06386_/X sky130_fd_sc_hd__clkbuf_2
X_05337_ _10007_/Q VGND VGND VPWR VPWR _05337_/Y sky130_fd_sc_hd__clkinv_2
X_08125_ _09459_/A _08064_/X _08122_/X _08124_/X VGND VGND VPWR VPWR _08135_/C sky130_fd_sc_hd__o211a_1
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05268_ _05346_/A _05307_/B VGND VGND VPWR VPWR _05909_/A sky130_fd_sc_hd__or2_1
X_08056_ _07359_/Y _08054_/X _07412_/Y _08055_/X VGND VGND VPWR VPWR _08056_/X sky130_fd_sc_hd__o22a_1
X_07007_ _07983_/A _06280_/B _07006_/Y _06037_/B VGND VGND VPWR VPWR _07007_/X sky130_fd_sc_hd__o22a_1
X_05199_ _05305_/A _06780_/B VGND VGND VPWR VPWR _05748_/A sky130_fd_sc_hd__or2_2
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput127 user_clock VGND VGND VPWR VPWR input127/X sky130_fd_sc_hd__buf_2
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput116 sram_ro_data[30] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__buf_2
Xinput105 sram_ro_data[20] VGND VGND VPWR VPWR input105/X sky130_fd_sc_hd__clkbuf_2
Xinput149 wb_adr_i[25] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__clkbuf_1
Xinput138 wb_adr_i[15] VGND VGND VPWR VPWR _08401_/A sky130_fd_sc_hd__clkbuf_1
X_08958_ _08958_/A _09290_/B VGND VGND VPWR VPWR _08960_/A sky130_fd_sc_hd__or2_1
X_08889_ _08900_/A VGND VGND VPWR VPWR _09052_/B sky130_fd_sc_hd__inv_2
X_07909_ _07409_/Y _07828_/X _07364_/Y _07829_/X VGND VGND VPWR VPWR _07909_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10216_ _10290_/CLK _10216_/D repeater402/X VGND VGND VPWR VPWR _10216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10147_ _10491_/CLK _10147_/D repeater403/X VGND VGND VPWR VPWR _10147_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10078_ _10411_/CLK _10078_/D repeater407/X VGND VGND VPWR VPWR _10078_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06240_ _07528_/A _06235_/Y _06147_/X _07584_/B VGND VGND VPWR VPWR _09991_/D sky130_fd_sc_hd__o22ai_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06171_ _10010_/Q _06168_/X _09658_/A1 _06169_/Y VGND VGND VPWR VPWR _10010_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05122_ _05119_/Y _05120_/Y _10469_/Q _10432_/Q _05121_/Y VGND VGND VPWR VPWR _05122_/X
+ sky130_fd_sc_hd__a32o_1
X_09930_ _10119_/CLK _09930_/D repeater402/X VGND VGND VPWR VPWR _09930_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05053_ _05053_/A VGND VGND VPWR VPWR _05054_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09861_ _10268_/CLK _09861_/D repeater404/X VGND VGND VPWR VPWR _09861_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10119_/CLK _09792_/D repeater403/X VGND VGND VPWR VPWR _09792_/Q sky130_fd_sc_hd__dfrtp_1
X_08812_ _08812_/A VGND VGND VPWR VPWR _09256_/A sky130_fd_sc_hd__inv_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05955_ _10132_/Q _05953_/X _09547_/A1 _05954_/Y VGND VGND VPWR VPWR _10132_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08743_ _08743_/A VGND VGND VPWR VPWR _09093_/A sky130_fd_sc_hd__clkbuf_4
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04906_ _10486_/Q _04902_/X _09579_/X _04904_/X VGND VGND VPWR VPWR _10486_/D sky130_fd_sc_hd__a22o_1
X_05886_ _05886_/A VGND VGND VPWR VPWR _05886_/X sky130_fd_sc_hd__clkbuf_2
X_08674_ _08831_/B VGND VGND VPWR VPWR _08674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _07384_/Y _07620_/X _07306_/Y _07621_/X _07624_/X VGND VGND VPWR VPWR _07625_/X
+ sky130_fd_sc_hd__o221a_1
X_04837_ _09678_/X _04835_/Y _09536_/A3 _10511_/Q _04836_/X VGND VGND VPWR VPWR _10511_/D
+ sky130_fd_sc_hd__a32o_1
X_07556_ _07565_/A _07575_/B VGND VGND VPWR VPWR _07610_/A sky130_fd_sc_hd__or2_1
XFILLER_22_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06507_ _09848_/Q _06504_/X _09581_/X _06506_/X VGND VGND VPWR VPWR _09848_/D sky130_fd_sc_hd__a22o_1
X_09226_ _09226_/A _09226_/B VGND VGND VPWR VPWR _09237_/A sky130_fd_sc_hd__or2_2
X_07487_ _10420_/Q VGND VGND VPWR VPWR _07487_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06438_ _06438_/A VGND VGND VPWR VPWR _06439_/B sky130_fd_sc_hd__buf_2
XFILLER_135_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09157_ _09157_/A _09157_/B VGND VGND VPWR VPWR _09161_/B sky130_fd_sc_hd__or2_1
X_06369_ _09922_/Q _06362_/A _09660_/A1 _06363_/A VGND VGND VPWR VPWR _09922_/D sky130_fd_sc_hd__a22o_1
XFILLER_181_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09088_ _09417_/A _09088_/B VGND VGND VPWR VPWR _09090_/A sky130_fd_sc_hd__or2_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08108_ _07256_/Y _08076_/X _07237_/Y _08077_/X VGND VGND VPWR VPWR _08108_/X sky130_fd_sc_hd__o22a_1
XFILLER_150_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08039_ _08046_/A _10002_/Q _08045_/C _10006_/Q VGND VGND VPWR VPWR _08207_/A sky130_fd_sc_hd__or4_4
XFILLER_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ _10364_/CLK _10001_/D repeater410/X VGND VGND VPWR VPWR _10001_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05740_ _05775_/A _05740_/B VGND VGND VPWR VPWR _05742_/A sky130_fd_sc_hd__or2_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05671_ _09770_/Q _05671_/B VGND VGND VPWR VPWR _05671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08390_ _08505_/A _09085_/B _08493_/B VGND VGND VPWR VPWR _08916_/A sky130_fd_sc_hd__or3_1
X_07410_ _07408_/Y _06095_/A _07409_/Y _05775_/B VGND VGND VPWR VPWR _07410_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07341_ _07339_/Y _05952_/B _07340_/Y _06037_/B VGND VGND VPWR VPWR _07341_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_148_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07272_ _10009_/Q VGND VGND VPWR VPWR _07272_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09011_ _09011_/A VGND VGND VPWR VPWR _09206_/A sky130_fd_sc_hd__clkbuf_2
X_06223_ _09991_/Q VGND VGND VPWR VPWR _07528_/A sky130_fd_sc_hd__inv_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06154_ _06313_/A _06154_/B VGND VGND VPWR VPWR _06156_/A sky130_fd_sc_hd__or2_2
XFILLER_191_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05105_ _06630_/A _06630_/B _09798_/Q VGND VGND VPWR VPWR _05105_/X sky130_fd_sc_hd__or3b_1
X_06085_ _10051_/Q _06080_/X _06684_/B1 _06081_/Y VGND VGND VPWR VPWR _10051_/D sky130_fd_sc_hd__a22o_1
X_09913_ _10397_/CLK _09913_/D repeater407/X VGND VGND VPWR VPWR _09913_/Q sky130_fd_sc_hd__dfrtp_1
X_05036_ _06668_/A VGND VGND VPWR VPWR _05053_/A sky130_fd_sc_hd__clkbuf_2
X_09844_ _10350_/CLK _09844_/D repeater405/X VGND VGND VPWR VPWR _09844_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06987_ _10215_/Q VGND VGND VPWR VPWR _06987_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09775_ _10023_/CLK _09775_/D _05034_/A VGND VGND VPWR VPWR _09775_/Q sky130_fd_sc_hd__dfstp_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05938_ _10142_/Q _05930_/A _09661_/A1 _05931_/A VGND VGND VPWR VPWR _10142_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08726_ _08732_/A _08849_/B VGND VGND VPWR VPWR _09397_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08657_ _09236_/A _08675_/A VGND VGND VPWR VPWR _08672_/B sky130_fd_sc_hd__or2_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05869_ _10183_/Q _05866_/X _09658_/A1 _05867_/Y VGND VGND VPWR VPWR _10183_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07608_/A _07608_/B VGND VGND VPWR VPWR _07825_/A sky130_fd_sc_hd__or2_2
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08588_ _08752_/A _08959_/B _08587_/X VGND VGND VPWR VPWR _08588_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07539_ _07539_/A _07601_/B VGND VGND VPWR VPWR _07819_/A sky130_fd_sc_hd__or2_1
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ _04811_/A1 _10481_/D _05459_/A VGND VGND VPWR VPWR _10481_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09209_ _09306_/A _09407_/C _09209_/C _09209_/D VGND VGND VPWR VPWR _09209_/X sky130_fd_sc_hd__or4_1
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput217 _09490_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_173_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _09530_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_2
Xoutput228 _09510_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_126_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput239 _09460_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_175_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06910_ _06909_/Y _06045_/B _10333_/Q _05151_/X VGND VGND VPWR VPWR _06910_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07890_ _07403_/Y _07777_/X _07371_/Y _07778_/X _07889_/X VGND VGND VPWR VPWR _07912_/A
+ sky130_fd_sc_hd__o221a_1
X_06841_ input106/X _05153_/A input17/X _06698_/X VGND VGND VPWR VPWR _06841_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06772_ input18/X _06698_/X input41/X _09699_/S _06771_/X VGND VGND VPWR VPWR _06775_/C
+ sky130_fd_sc_hd__a221o_1
X_09560_ _10429_/Q _10276_/Q hold1/A VGND VGND VPWR VPWR _09560_/X sky130_fd_sc_hd__mux2_1
X_09491_ _09491_/A VGND VGND VPWR VPWR _09492_/A sky130_fd_sc_hd__clkbuf_1
X_05723_ _10269_/Q _05717_/X _09546_/X _05718_/X VGND VGND VPWR VPWR _10269_/D sky130_fd_sc_hd__o22a_1
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08511_ _08583_/A VGND VGND VPWR VPWR _08752_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08442_ _09085_/C _08494_/A _09085_/D VGND VGND VPWR VPWR _08783_/A sky130_fd_sc_hd__or3_4
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05654_ _05654_/A VGND VGND VPWR VPWR _05655_/A sky130_fd_sc_hd__inv_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08373_ _09085_/B VGND VGND VPWR VPWR _08631_/C sky130_fd_sc_hd__inv_2
X_05585_ _10345_/Q _05578_/A _09660_/A1 _05579_/A VGND VGND VPWR VPWR _10345_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07324_ _07324_/A _07324_/B _07324_/C _07323_/X VGND VGND VPWR VPWR _07420_/B sky130_fd_sc_hd__or4b_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07255_ _07932_/A _06280_/B _07251_/Y _05138_/A _07254_/X VGND VGND VPWR VPWR _07262_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_149_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06206_ _06313_/A _06206_/B VGND VGND VPWR VPWR _06208_/A sky130_fd_sc_hd__or2_4
XFILLER_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07186_ _07184_/Y _05728_/B _07185_/Y _06472_/B VGND VGND VPWR VPWR _07186_/X sky130_fd_sc_hd__o22a_2
XFILLER_129_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06137_ _06137_/A _06139_/A _06260_/C VGND VGND VPWR VPWR _06137_/X sky130_fd_sc_hd__or3_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06068_ _06068_/A VGND VGND VPWR VPWR _06069_/A sky130_fd_sc_hd__inv_2
X_05019_ _05541_/A _05121_/A VGND VGND VPWR VPWR _05021_/A sky130_fd_sc_hd__or2_2
XFILLER_132_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09827_ _10405_/CLK _09827_/D hold41/X VGND VGND VPWR VPWR _09827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09758_ _09919_/CLK _09758_/D VGND VGND VPWR VPWR _09758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _08717_/A _08831_/B VGND VGND VPWR VPWR _09115_/A sky130_fd_sc_hd__or2_1
X_09689_ _08368_/X input192/X _09698_/S VGND VGND VPWR VPWR _09689_/X sky130_fd_sc_hd__mux2_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10464_ _10471_/CLK _10464_/D repeater409/X VGND VGND VPWR VPWR _10464_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_163_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10395_ _04811_/A1 _10395_/D _05457_/X VGND VGND VPWR VPWR _10395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05370_ _05370_/A VGND VGND VPWR VPWR _05370_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07040_ _07040_/A _07040_/B _07040_/C _07040_/D VGND VGND VPWR VPWR _07158_/A sky130_fd_sc_hd__or4_2
XFILLER_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08991_ _09083_/C _08900_/A _09789_/Q VGND VGND VPWR VPWR _09362_/C sky130_fd_sc_hd__o21ai_4
XFILLER_141_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07942_ _07122_/Y _07627_/A _07126_/Y _07788_/A _07941_/X VGND VGND VPWR VPWR _07951_/A
+ sky130_fd_sc_hd__o221a_1
X_07873_ _05326_/Y _07806_/X _05282_/Y _07807_/X VGND VGND VPWR VPWR _07873_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06824_ _10165_/Q VGND VGND VPWR VPWR _06824_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09612_ _08328_/Y _10328_/Q _09700_/S VGND VGND VPWR VPWR _09612_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09543_ _10323_/Q _09581_/X _09679_/S VGND VGND VPWR VPWR _09543_/X sky130_fd_sc_hd__mux2_1
X_06755_ _06753_/Y _05728_/B _06754_/Y _05839_/B VGND VGND VPWR VPWR _06755_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09474_ _09474_/A VGND VGND VPWR VPWR _09474_/X sky130_fd_sc_hd__clkbuf_1
X_06686_ input10/X _06838_/A _10458_/Q _05089_/A VGND VGND VPWR VPWR _06686_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05706_ _10279_/Q _05701_/X _09545_/X _05702_/X VGND VGND VPWR VPWR _10279_/D sky130_fd_sc_hd__o22a_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08425_ _08571_/C _08476_/A _08424_/X VGND VGND VPWR VPWR _09236_/B sky130_fd_sc_hd__o21ai_2
X_05637_ _10316_/Q _05628_/A _09659_/A1 _05629_/A VGND VGND VPWR VPWR _10316_/D sky130_fd_sc_hd__a22o_1
X_08356_ _08356_/A VGND VGND VPWR VPWR _09698_/S sky130_fd_sc_hd__clkinv_8
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05568_ _05569_/A VGND VGND VPWR VPWR _05568_/X sky130_fd_sc_hd__clkbuf_2
X_07307_ _07306_/Y _06024_/B _06780_/X VGND VGND VPWR VPWR _07307_/Y sky130_fd_sc_hd__o21ai_2
X_05499_ _09690_/X _10384_/Q _05512_/S VGND VGND VPWR VPWR _05500_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08287_ _07194_/Y _08207_/X _07209_/Y _08208_/X VGND VGND VPWR VPWR _08287_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07238_ _10026_/Q VGND VGND VPWR VPWR _07238_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07169_ _10099_/Q _05070_/Y _10445_/Q _06688_/X _07168_/X VGND VGND VPWR VPWR _07193_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10180_ _10184_/CLK _10180_/D repeater407/X VGND VGND VPWR VPWR _10180_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10447_ _10487_/CLK _10447_/D repeater409/X VGND VGND VPWR VPWR _10447_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_108_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10378_ _04811_/A1 _10378_/D _05524_/X VGND VGND VPWR VPWR _10378_/Q sky130_fd_sc_hd__dfrtp_1
X_04870_ _04870_/A VGND VGND VPWR VPWR _04871_/B sky130_fd_sc_hd__buf_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06540_ _06540_/A VGND VGND VPWR VPWR _06541_/A sky130_fd_sc_hd__inv_2
X_06471_ _06471_/A VGND VGND VPWR VPWR _06472_/B sky130_fd_sc_hd__buf_2
X_08210_ _06791_/Y _08205_/X _06803_/Y _08206_/X _08209_/X VGND VGND VPWR VPWR _08217_/C
+ sky130_fd_sc_hd__o221a_1
X_05422_ _10411_/Q _05420_/X _09578_/X _05421_/Y VGND VGND VPWR VPWR _10411_/D sky130_fd_sc_hd__a22o_1
XANTENNA_190 _07779_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09190_ _09273_/A _09362_/B VGND VGND VPWR VPWR _09317_/A sky130_fd_sc_hd__or2_1
X_05353_ _05343_/Y _05549_/A _05345_/Y _05419_/B _05352_/X VGND VGND VPWR VPWR _05364_/C
+ sky130_fd_sc_hd__o221a_1
X_08141_ _07003_/Y _08069_/X _06967_/Y _08070_/X VGND VGND VPWR VPWR _08141_/X sky130_fd_sc_hd__o22a_1
X_05284_ _05311_/B _05284_/B VGND VGND VPWR VPWR _06010_/A sky130_fd_sc_hd__or2_2
X_08072_ _07387_/Y _08067_/X _07338_/Y _08068_/X _08071_/X VGND VGND VPWR VPWR _08072_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07023_ _09824_/Q VGND VGND VPWR VPWR _07023_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08974_ _09372_/A _08974_/B _09005_/A VGND VGND VPWR VPWR _08978_/B sky130_fd_sc_hd__or3_2
XFILLER_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07925_ _07194_/Y _07805_/X _07923_/Y _07523_/A _07924_/X VGND VGND VPWR VPWR _07926_/D
+ sky130_fd_sc_hd__o221a_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07856_ _10062_/Q VGND VGND VPWR VPWR _07856_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06807_ _06802_/Y _06291_/B _06803_/Y _05728_/B _06806_/X VGND VGND VPWR VPWR _06814_/C
+ sky130_fd_sc_hd__o221a_1
X_07787_ _07787_/A VGND VGND VPWR VPWR _07787_/X sky130_fd_sc_hd__buf_4
X_04999_ _10448_/Q _04994_/X _09579_/X _04996_/X VGND VGND VPWR VPWR _10448_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06738_ _06736_/Y _05852_/B _06737_/Y _05794_/B VGND VGND VPWR VPWR _06738_/X sky130_fd_sc_hd__o22a_1
X_09526_ _09526_/A VGND VGND VPWR VPWR _09526_/X sky130_fd_sc_hd__clkbuf_2
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09457_ _09457_/A VGND VGND VPWR VPWR _09458_/A sky130_fd_sc_hd__clkbuf_1
X_08408_ _08408_/A VGND VGND VPWR VPWR _08408_/Y sky130_fd_sc_hd__inv_2
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06669_ _06677_/A VGND VGND VPWR VPWR _06670_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09388_ _09388_/A _09388_/B VGND VGND VPWR VPWR _09389_/B sky130_fd_sc_hd__or2_1
X_08339_ _09803_/Q _08338_/B _08340_/A VGND VGND VPWR VPWR _08339_/X sky130_fd_sc_hd__o21a_1
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10301_ _10504_/CLK hold47/X repeater404/X VGND VGND VPWR VPWR _10301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10232_ _10288_/CLK _10232_/D repeater406/X VGND VGND VPWR VPWR _10232_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10163_ _10238_/CLK _10163_/D repeater403/X VGND VGND VPWR VPWR _10163_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10094_ _10289_/CLK _10094_/D repeater402/X VGND VGND VPWR VPWR _10094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05971_ _05971_/A VGND VGND VPWR VPWR _05971_/X sky130_fd_sc_hd__clkbuf_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _09499_/A _07658_/X _09519_/A _07659_/X VGND VGND VPWR VPWR _07710_/X sky130_fd_sc_hd__o22a_1
X_04922_ _09533_/A _09683_/S VGND VGND VPWR VPWR _04923_/A sky130_fd_sc_hd__nand2_1
X_08690_ _09233_/C VGND VGND VPWR VPWR _08753_/C sky130_fd_sc_hd__inv_2
X_04853_ _10508_/Q _04851_/X _09584_/X _04852_/X VGND VGND VPWR VPWR _10508_/D sky130_fd_sc_hd__o22a_1
X_07641_ _07801_/A VGND VGND VPWR VPWR _07641_/X sky130_fd_sc_hd__clkbuf_2
X_07572_ _07572_/A VGND VGND VPWR VPWR _07779_/A sky130_fd_sc_hd__buf_4
XFILLER_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09311_ _09311_/A _09311_/B _09311_/C _09311_/D VGND VGND VPWR VPWR _09408_/A sky130_fd_sc_hd__or4_4
X_06523_ _09837_/Q _06517_/X _09547_/A1 _06519_/X VGND VGND VPWR VPWR _09837_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_33_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10224_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06454_ _09787_/D VGND VGND VPWR VPWR _07450_/B sky130_fd_sc_hd__inv_2
X_09242_ _09224_/Y _09236_/Y _09237_/X _09172_/D VGND VGND VPWR VPWR _09327_/D sky130_fd_sc_hd__a31o_1
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05405_ _10416_/Q _05396_/X hold45/A _05398_/X VGND VGND VPWR VPWR _10416_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09173_ _08883_/A _08520_/B _08466_/A _09263_/A VGND VGND VPWR VPWR _09327_/C sky130_fd_sc_hd__o22ai_1
X_06385_ _06380_/X _09595_/X _09650_/X _09910_/Q VGND VGND VPWR VPWR _09910_/D sky130_fd_sc_hd__o22a_1
X_05336_ _05336_/A _05357_/B VGND VGND VPWR VPWR _06502_/A sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_48_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10471_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08124_ _09463_/A _08067_/X _09505_/A _08068_/X _08123_/X VGND VGND VPWR VPWR _08124_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05267_ _10154_/Q VGND VGND VPWR VPWR _05267_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08055_ _08174_/A VGND VGND VPWR VPWR _08055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07006_ _10080_/Q VGND VGND VPWR VPWR _07006_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05198_ _05198_/A VGND VGND VPWR VPWR _06780_/B sky130_fd_sc_hd__buf_2
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput117 sram_ro_data[31] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__buf_2
Xinput106 sram_ro_data[21] VGND VGND VPWR VPWR input106/X sky130_fd_sc_hd__buf_2
Xinput128 usr1_vcc_pwrgood VGND VGND VPWR VPWR input128/X sky130_fd_sc_hd__buf_6
Xinput139 wb_adr_i[16] VGND VGND VPWR VPWR _08399_/B sky130_fd_sc_hd__clkbuf_1
X_08957_ _08957_/A _08957_/B VGND VGND VPWR VPWR _09290_/B sky130_fd_sc_hd__nor2_1
X_08888_ _08888_/A _08888_/B _08890_/A VGND VGND VPWR VPWR _08900_/A sky130_fd_sc_hd__or3_4
X_07908_ _07332_/Y _07768_/X _07382_/Y _07769_/X _07907_/X VGND VGND VPWR VPWR _07911_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07839_ _06747_/Y _07787_/X _06734_/Y _07788_/X _07838_/X VGND VGND VPWR VPWR _07848_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09509_ _09509_/A VGND VGND VPWR VPWR _09510_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10215_ _10508_/CLK _10215_/D repeater402/X VGND VGND VPWR VPWR _10215_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10146_ _10491_/CLK _10146_/D repeater403/X VGND VGND VPWR VPWR _10146_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10077_ _10411_/CLK _10077_/D repeater407/X VGND VGND VPWR VPWR _10077_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06170_ _10011_/Q _06168_/X _09545_/A1 _06169_/Y VGND VGND VPWR VPWR _10011_/D sky130_fd_sc_hd__a22o_1
XFILLER_171_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05121_ _05121_/A VGND VGND VPWR VPWR _05121_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05052_ _10426_/Q _05040_/X _09639_/X _05042_/X VGND VGND VPWR VPWR _10426_/D sky130_fd_sc_hd__a22o_2
X_09860_ _10268_/CLK _09860_/D repeater404/X VGND VGND VPWR VPWR _09860_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _09102_/A _09085_/B _08683_/A VGND VGND VPWR VPWR _08811_/X sky130_fd_sc_hd__or3b_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _10510_/CLK _09791_/D _05034_/A VGND VGND VPWR VPWR _09791_/Q sky130_fd_sc_hd__dfrtp_4
X_05954_ _05954_/A VGND VGND VPWR VPWR _05954_/Y sky130_fd_sc_hd__inv_2
X_08742_ _08742_/A _09420_/C VGND VGND VPWR VPWR _08745_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _08829_/A VGND VGND VPWR VPWR _08831_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04905_ _10487_/Q _04902_/X _09580_/X _04904_/X VGND VGND VPWR VPWR _10487_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05885_ _05885_/A VGND VGND VPWR VPWR _05886_/A sky130_fd_sc_hd__inv_2
X_07624_ _07319_/Y _07622_/X _07344_/Y _07623_/X VGND VGND VPWR VPWR _07624_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04836_ _05031_/A _04836_/B VGND VGND VPWR VPWR _04836_/X sky130_fd_sc_hd__or2_1
X_07555_ _07806_/A VGND VGND VPWR VPWR _07646_/A sky130_fd_sc_hd__buf_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06506_ _06506_/A VGND VGND VPWR VPWR _06506_/X sky130_fd_sc_hd__clkbuf_2
X_07486_ _10419_/Q _05376_/X _09770_/Q _09774_/Q VGND VGND VPWR VPWR _09774_/D sky130_fd_sc_hd__a31o_1
XFILLER_34_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06437_ _09876_/Q _06431_/X _09574_/X _06432_/Y VGND VGND VPWR VPWR _09876_/D sky130_fd_sc_hd__a22o_1
X_09225_ _09225_/A VGND VGND VPWR VPWR _09225_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09156_ _09324_/A _09156_/B _09156_/C _09155_/X VGND VGND VPWR VPWR _09157_/B sky130_fd_sc_hd__or4b_1
X_06368_ _09923_/Q _06361_/X _09550_/A0 _06363_/X VGND VGND VPWR VPWR _09923_/D sky130_fd_sc_hd__a22o_1
X_09087_ _09434_/A _09087_/B VGND VGND VPWR VPWR _09088_/B sky130_fd_sc_hd__or2_1
X_06299_ _09963_/Q _06292_/X _09550_/A0 _06294_/X VGND VGND VPWR VPWR _09963_/D sky130_fd_sc_hd__a22o_1
X_05319_ _05315_/Y _05864_/A _05317_/Y _05829_/A VGND VGND VPWR VPWR _05319_/X sky130_fd_sc_hd__o22a_1
X_08107_ _07221_/Y _08064_/X _08104_/X _08106_/X VGND VGND VPWR VPWR _08117_/C sky130_fd_sc_hd__o211a_1
XFILLER_107_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08038_ _08038_/A _08044_/B _08038_/C VGND VGND VPWR VPWR _08206_/A sky130_fd_sc_hd__or3_4
XFILLER_150_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10000_ _10000_/CLK _10000_/D repeater410/X VGND VGND VPWR VPWR _10000_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09989_ _10397_/CLK _09989_/D repeater407/X VGND VGND VPWR VPWR _09989_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10129_ _10238_/CLK _10129_/D repeater403/X VGND VGND VPWR VPWR _10129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05670_ _05670_/A VGND VGND VPWR VPWR _05670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07340_ _10077_/Q VGND VGND VPWR VPWR _07340_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09010_ _09010_/A VGND VGND VPWR VPWR _09010_/X sky130_fd_sc_hd__buf_2
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07271_ _10203_/Q VGND VGND VPWR VPWR _07271_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06222_ _06243_/A _06245_/B VGND VGND VPWR VPWR _06238_/A sky130_fd_sc_hd__or2_1
X_06153_ _06153_/A VGND VGND VPWR VPWR _06154_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_144_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05104_ _05338_/A VGND VGND VPWR VPWR _06630_/B sky130_fd_sc_hd__buf_4
XFILLER_171_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06084_ _10052_/Q _06080_/X _06683_/B1 _06081_/Y VGND VGND VPWR VPWR _10052_/D sky130_fd_sc_hd__a22o_1
X_09912_ _10397_/CLK _09912_/D repeater409/X VGND VGND VPWR VPWR _09912_/Q sky130_fd_sc_hd__dfrtp_1
X_05035_ _06679_/B split1/X VGND VGND VPWR VPWR _06668_/A sky130_fd_sc_hd__nor2_2
XFILLER_140_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09843_ _10350_/CLK _09843_/D repeater404/X VGND VGND VPWR VPWR _09843_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _10406_/CLK _09774_/D _06670_/X VGND VGND VPWR VPWR _09774_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _10054_/Q VGND VGND VPWR VPWR _06986_/Y sky130_fd_sc_hd__inv_4
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05937_ _10143_/Q _05930_/A _09660_/A1 _05931_/A VGND VGND VPWR VPWR _10143_/D sky130_fd_sc_hd__a22o_1
X_08725_ _08725_/A _09124_/A VGND VGND VPWR VPWR _08727_/A sky130_fd_sc_hd__nand2_1
X_08656_ _08656_/A VGND VGND VPWR VPWR _08675_/A sky130_fd_sc_hd__inv_2
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05868_ _10184_/Q _05866_/X _09545_/A1 _05867_/Y VGND VGND VPWR VPWR _10184_/D sky130_fd_sc_hd__a22o_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _05189_/Y _06232_/A _05356_/Y _07519_/A _07606_/X VGND VGND VPWR VPWR _07615_/C
+ sky130_fd_sc_hd__o221a_1
X_08587_ _09010_/A _09024_/A _08584_/Y _09200_/A _09025_/A VGND VGND VPWR VPWR _08587_/X
+ sky130_fd_sc_hd__o2111a_1
X_04819_ _04818_/Y _09666_/X _09665_/X VGND VGND VPWR VPWR _05213_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07538_ _07787_/A VGND VGND VPWR VPWR _07627_/A sky130_fd_sc_hd__clkbuf_4
X_05799_ _10225_/Q _05795_/X _09580_/X _05797_/X VGND VGND VPWR VPWR _10225_/D sky130_fd_sc_hd__a22o_1
X_07469_ _10420_/Q _05430_/Y _07468_/Y _09771_/Q VGND VGND VPWR VPWR _09771_/D sky130_fd_sc_hd__a31o_1
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ _09407_/A _09371_/A _09306_/B _08559_/X VGND VGND VPWR VPWR _09209_/D sky130_fd_sc_hd__or4b_1
X_10480_ _10483_/CLK _10480_/D _05034_/A VGND VGND VPWR VPWR _10480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09139_ _09139_/A _09139_/B VGND VGND VPWR VPWR _09140_/C sky130_fd_sc_hd__or2_1
XFILLER_185_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput207 _09566_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_2
Xoutput218 _09567_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_2
Xoutput229 _09458_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06840_ _10442_/Q _05091_/X _09557_/X _06633_/X _06839_/X VGND VGND VPWR VPWR _06840_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06771_ input9/X _06838_/A _10449_/Q _06688_/A VGND VGND VPWR VPWR _06771_/X sky130_fd_sc_hd__a22o_2
X_09490_ _09490_/A VGND VGND VPWR VPWR _09490_/X sky130_fd_sc_hd__clkbuf_1
X_05722_ _10270_/Q _05717_/X _09547_/X _05718_/X VGND VGND VPWR VPWR _10270_/D sky130_fd_sc_hd__o22a_1
X_08510_ _08685_/B VGND VGND VPWR VPWR _08583_/A sky130_fd_sc_hd__clkbuf_4
X_05653_ _05654_/A VGND VGND VPWR VPWR _05653_/X sky130_fd_sc_hd__clkbuf_2
X_08441_ _08631_/A VGND VGND VPWR VPWR _09085_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08372_ _09790_/Q input189/X _09789_/Q input171/X _08371_/X VGND VGND VPWR VPWR _08372_/X
+ sky130_fd_sc_hd__a221o_1
X_05584_ _10346_/Q _05577_/X _09550_/A0 _05579_/X VGND VGND VPWR VPWR _10346_/D sky130_fd_sc_hd__a22o_1
X_07323_ _07318_/Y _06167_/B _07319_/Y _05968_/B _07322_/X VGND VGND VPWR VPWR _07323_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07254_ _07252_/Y _06401_/A _07253_/Y _06393_/B VGND VGND VPWR VPWR _07254_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06205_ _06205_/A VGND VGND VPWR VPWR _06206_/B sky130_fd_sc_hd__buf_2
XFILLER_191_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07185_ _09864_/Q VGND VGND VPWR VPWR _07185_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06136_ _10021_/Q VGND VGND VPWR VPWR _06260_/C sky130_fd_sc_hd__inv_2
XFILLER_117_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06067_ _06068_/A VGND VGND VPWR VPWR _06067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05018_ _05118_/A _05198_/A VGND VGND VPWR VPWR _05121_/A sky130_fd_sc_hd__or2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09826_ _10405_/CLK _09826_/D hold41/X VGND VGND VPWR VPWR _09826_/Q sky130_fd_sc_hd__dfrtp_1
X_09757_ _09781_/CLK _09757_/D VGND VGND VPWR VPWR _09757_/Q sky130_fd_sc_hd__dfxtp_1
X_06969_ _10132_/Q VGND VGND VPWR VPWR _06969_/Y sky130_fd_sc_hd__inv_4
XFILLER_100_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _09095_/A _08824_/B _08705_/X _09111_/A _09158_/A VGND VGND VPWR VPWR _08708_/X
+ sky130_fd_sc_hd__o2111a_1
X_09688_ _08366_/X input191/X _09698_/S VGND VGND VPWR VPWR _09688_/X sky130_fd_sc_hd__mux2_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08556_/B _08789_/B _08641_/B VGND VGND VPWR VPWR _08781_/B sky130_fd_sc_hd__a21bo_2
XFILLER_120_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10463_ _10471_/CLK _10463_/D repeater409/X VGND VGND VPWR VPWR _10463_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10394_ _04811_/A1 _10394_/D _05460_/X VGND VGND VPWR VPWR _10394_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08990_ _09222_/A _08990_/B VGND VGND VPWR VPWR _08992_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07941_ _07128_/Y _07527_/A _07111_/Y _07629_/A VGND VGND VPWR VPWR _07941_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07872_ _10337_/Q VGND VGND VPWR VPWR _07872_/Y sky130_fd_sc_hd__inv_2
X_06823_ _10121_/Q VGND VGND VPWR VPWR _06823_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09611_ _09610_/X _09917_/Q _09776_/Q VGND VGND VPWR VPWR _09611_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06754_ _10200_/Q VGND VGND VPWR VPWR _06754_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09542_ _10322_/Q _09580_/X _09679_/S VGND VGND VPWR VPWR _09542_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05705_ _10280_/Q _05701_/X _09541_/X _05702_/X VGND VGND VPWR VPWR _10280_/D sky130_fd_sc_hd__o22a_1
X_09473_ _09473_/A VGND VGND VPWR VPWR _09474_/A sky130_fd_sc_hd__clkbuf_1
X_06685_ _09766_/Q _06681_/A _09536_/A3 _06681_/Y VGND VGND VPWR VPWR _09766_/D sky130_fd_sc_hd__a22o_1
X_08424_ _08537_/C _08424_/B VGND VGND VPWR VPWR _08424_/X sky130_fd_sc_hd__or2_1
X_05636_ _10317_/Q _05628_/A _09661_/A1 _05629_/A VGND VGND VPWR VPWR _10317_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08355_ _09789_/Q _05489_/X _08353_/X _08354_/X VGND VGND VPWR VPWR _08355_/X sky130_fd_sc_hd__a211o_1
X_05567_ _05775_/A _05567_/B VGND VGND VPWR VPWR _05569_/A sky130_fd_sc_hd__or2_1
X_07306_ _10082_/Q VGND VGND VPWR VPWR _07306_/Y sky130_fd_sc_hd__inv_4
XFILLER_192_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05498_ _05498_/A VGND VGND VPWR VPWR _05498_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08286_ _07185_/Y _08199_/X _07214_/Y _08200_/X _08285_/X VGND VGND VPWR VPWR _08291_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07237_ _10065_/Q VGND VGND VPWR VPWR _07237_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_164_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07168_ input5/X _06838_/X input63/X _06844_/X VGND VGND VPWR VPWR _07168_/X sky130_fd_sc_hd__a22o_1
X_06119_ _10029_/Q _06110_/A _09536_/A3 _06111_/A VGND VGND VPWR VPWR _10029_/D sky130_fd_sc_hd__a22o_1
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07099_ _09844_/Q VGND VGND VPWR VPWR _09465_/A sky130_fd_sc_hd__clkinv_4
XFILLER_160_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09809_ _09572_/A1 _09809_/D _06588_/X VGND VGND VPWR VPWR _09809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10446_ _10487_/CLK _10446_/D _05034_/A VGND VGND VPWR VPWR _10446_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10377_ _10404_/CLK _10377_/D hold41/X VGND VGND VPWR VPWR _10377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06470_ _09781_/Q _06453_/Y _09867_/Q _06468_/Y _06469_/X VGND VGND VPWR VPWR _09867_/D
+ sky130_fd_sc_hd__o221a_1
X_05421_ _05421_/A VGND VGND VPWR VPWR _05421_/Y sky130_fd_sc_hd__inv_2
XANTENNA_191 _07779_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_180 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08140_ _06950_/Y _08065_/X _06942_/Y _06188_/X VGND VGND VPWR VPWR _08140_/X sky130_fd_sc_hd__o22a_1
X_05352_ _05348_/Y _06328_/A _05350_/Y _06493_/A VGND VGND VPWR VPWR _05352_/X sky130_fd_sc_hd__o22a_1
X_05283_ _10089_/Q VGND VGND VPWR VPWR _05283_/Y sky130_fd_sc_hd__clkinv_4
X_08071_ _07321_/Y _08069_/X _07376_/Y _08070_/X VGND VGND VPWR VPWR _08071_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07022_ _09937_/Q VGND VGND VPWR VPWR _07022_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08973_ _08973_/A _09405_/B VGND VGND VPWR VPWR _08973_/X sky130_fd_sc_hd__or2_2
XFILLER_102_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07924_ _07253_/Y _07806_/X _07244_/Y _07807_/X VGND VGND VPWR VPWR _07924_/X sky130_fd_sc_hd__o22a_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold39 hold39/A VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _06736_/Y _07768_/X _06708_/A _07769_/X _07854_/X VGND VGND VPWR VPWR _07859_/C
+ sky130_fd_sc_hd__o221a_1
X_06806_ _06804_/Y _06503_/B _06805_/Y _05883_/B VGND VGND VPWR VPWR _06806_/X sky130_fd_sc_hd__o22a_1
X_07786_ _06830_/Y _07777_/X _06818_/Y _07778_/X _07785_/X VGND VGND VPWR VPWR _07833_/A
+ sky130_fd_sc_hd__o221a_2
X_04998_ _10449_/Q _04994_/X _09580_/X _04996_/X VGND VGND VPWR VPWR _10449_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06737_ _10226_/Q VGND VGND VPWR VPWR _06737_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09525_ input36/X input1/X VGND VGND VPWR VPWR _09526_/A sky130_fd_sc_hd__and2_1
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _09781_/CLK sky130_fd_sc_hd__clkbuf_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06668_ _06668_/A VGND VGND VPWR VPWR _06677_/A sky130_fd_sc_hd__clkbuf_2
X_09456_ _09456_/A VGND VGND VPWR VPWR _09456_/X sky130_fd_sc_hd__clkbuf_1
X_08407_ _08556_/B _08430_/B _08641_/A _08641_/C VGND VGND VPWR VPWR _08408_/A sky130_fd_sc_hd__or4_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05619_ _10327_/Q _05616_/X _09658_/A1 _05617_/Y VGND VGND VPWR VPWR _10327_/D sky130_fd_sc_hd__a22o_1
X_09387_ _09387_/A _09387_/B _09387_/C _09387_/D VGND VGND VPWR VPWR _09428_/D sky130_fd_sc_hd__or4_4
X_06599_ _06614_/A VGND VGND VPWR VPWR _06600_/A sky130_fd_sc_hd__clkbuf_1
X_08338_ _09803_/Q _08338_/B VGND VGND VPWR VPWR _08340_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08269_ _07351_/Y _08207_/X _07403_/Y _08208_/X VGND VGND VPWR VPWR _08269_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10300_ _10504_/CLK _10300_/D repeater404/X VGND VGND VPWR VPWR _10300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10231_ _10355_/CLK _10231_/D repeater406/X VGND VGND VPWR VPWR _10231_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10162_ _10238_/CLK _10162_/D repeater403/X VGND VGND VPWR VPWR _10162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10093_ _10289_/CLK _10093_/D repeater402/X VGND VGND VPWR VPWR _10093_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput390 _09742_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10429_ net399_2/A _10429_/D _05053_/A VGND VGND VPWR VPWR _10429_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _05970_/A VGND VGND VPWR VPWR _05971_/A sky130_fd_sc_hd__inv_2
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04921_ _09787_/Q _08356_/A VGND VGND VPWR VPWR _09683_/S sky130_fd_sc_hd__nor2_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04852_ _04852_/A VGND VGND VPWR VPWR _04852_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07640_ _10134_/Q VGND VGND VPWR VPWR _07640_/Y sky130_fd_sc_hd__inv_2
X_07571_ _07585_/C _07611_/A _07601_/A VGND VGND VPWR VPWR _07778_/A sky130_fd_sc_hd__or3_4
XFILLER_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09310_ _09407_/D _09371_/C _09439_/A _09369_/D VGND VGND VPWR VPWR _09313_/A sky130_fd_sc_hd__or4_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06522_ _09838_/Q _06517_/X _09579_/X _06519_/X VGND VGND VPWR VPWR _09838_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06453_ _09787_/Q VGND VGND VPWR VPWR _06453_/Y sky130_fd_sc_hd__inv_2
X_09241_ _09236_/Y _09233_/Y _09237_/X _09172_/B VGND VGND VPWR VPWR _09380_/C sky130_fd_sc_hd__a31o_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05404_ _05404_/A VGND VGND VPWR VPWR _05404_/X sky130_fd_sc_hd__clkbuf_1
X_09172_ _09172_/A _09172_/B _09380_/A _09172_/D VGND VGND VPWR VPWR _09174_/A sky130_fd_sc_hd__or4_1
X_06384_ _06380_/X _09597_/X _09650_/X _09911_/Q VGND VGND VPWR VPWR _09911_/D sky130_fd_sc_hd__o22a_1
X_05335_ _09841_/Q VGND VGND VPWR VPWR _05335_/Y sky130_fd_sc_hd__inv_2
X_08123_ _09499_/A _08069_/X _09497_/A _08070_/X VGND VGND VPWR VPWR _08123_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08054_ _08173_/A VGND VGND VPWR VPWR _08054_/X sky130_fd_sc_hd__clkbuf_2
X_07005_ _09973_/Q VGND VGND VPWR VPWR _07983_/A sky130_fd_sc_hd__clkinv_4
X_05266_ _06780_/B _05307_/B VGND VGND VPWR VPWR _06095_/A sky130_fd_sc_hd__or2_2
X_05197_ _10245_/Q VGND VGND VPWR VPWR _05197_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput118 sram_ro_data[3] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput107 sram_ro_data[22] VGND VGND VPWR VPWR input107/X sky130_fd_sc_hd__buf_2
Xinput129 usr1_vdd_pwrgood VGND VGND VPWR VPWR input129/X sky130_fd_sc_hd__buf_6
X_08956_ _08956_/A _09073_/B VGND VGND VPWR VPWR _08958_/A sky130_fd_sc_hd__or2_1
X_08887_ _08890_/A _08888_/B _08888_/A VGND VGND VPWR VPWR _09052_/A sky130_fd_sc_hd__o21a_1
X_07907_ _07907_/A _07932_/B VGND VGND VPWR VPWR _07907_/X sky130_fd_sc_hd__or2_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07838_ _06723_/Y _07749_/X _06712_/Y _07789_/X VGND VGND VPWR VPWR _07838_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09508_ _09508_/A VGND VGND VPWR VPWR _09508_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07769_ _07769_/A VGND VGND VPWR VPWR _07769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09439_ _09439_/A _09439_/B _09439_/C _09439_/D VGND VGND VPWR VPWR _09440_/A sky130_fd_sc_hd__or4_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_80 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10214_ _10508_/CLK _10214_/D repeater402/X VGND VGND VPWR VPWR _10214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10145_ _10491_/CLK _10145_/D repeater403/X VGND VGND VPWR VPWR _10145_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10076_ _10411_/CLK _10076_/D repeater407/X VGND VGND VPWR VPWR _10076_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05120_ _05292_/A VGND VGND VPWR VPWR _05120_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05051_ _05051_/A VGND VGND VPWR VPWR _05051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08810_ _09048_/A _08810_/B VGND VGND VPWR VPWR _09101_/A sky130_fd_sc_hd__nand2_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _10382_/CLK _09790_/D _06645_/X VGND VGND VPWR VPWR _09790_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05953_ _05954_/A VGND VGND VPWR VPWR _05953_/X sky130_fd_sc_hd__clkbuf_2
X_08741_ _09336_/B _08860_/A VGND VGND VPWR VPWR _09420_/C sky130_fd_sc_hd__nor2_2
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05884_ _05885_/A VGND VGND VPWR VPWR _05884_/X sky130_fd_sc_hd__clkbuf_2
X_08672_ _08809_/A _08672_/B VGND VGND VPWR VPWR _08829_/A sky130_fd_sc_hd__or2_1
X_04904_ _04904_/A VGND VGND VPWR VPWR _04904_/X sky130_fd_sc_hd__clkbuf_2
X_07623_ _07783_/A VGND VGND VPWR VPWR _07623_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04835_ _04836_/B VGND VGND VPWR VPWR _04835_/Y sky130_fd_sc_hd__inv_2
X_07554_ _07592_/A _07602_/C _07554_/C VGND VGND VPWR VPWR _07806_/A sky130_fd_sc_hd__or3_1
XFILLER_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06505_ _06505_/A VGND VGND VPWR VPWR _06506_/A sky130_fd_sc_hd__inv_2
X_07485_ _07485_/A VGND VGND VPWR VPWR _09770_/D sky130_fd_sc_hd__inv_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09224_ _09233_/C _09224_/B VGND VGND VPWR VPWR _09224_/Y sky130_fd_sc_hd__nor2_4
X_06436_ _09877_/Q _06431_/X _06684_/B1 _06432_/Y VGND VGND VPWR VPWR _09877_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09155_ _09155_/A _09155_/B VGND VGND VPWR VPWR _09155_/X sky130_fd_sc_hd__or2_1
X_06367_ _09924_/Q _06361_/X _09547_/A1 _06363_/X VGND VGND VPWR VPWR _09924_/D sky130_fd_sc_hd__a22o_1
XFILLER_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09086_ _09086_/A _09086_/B _09432_/C _09297_/A VGND VGND VPWR VPWR _09087_/B sky130_fd_sc_hd__or4_1
X_06298_ _09964_/Q _06292_/X _09547_/A1 _06294_/X VGND VGND VPWR VPWR _09964_/D sky130_fd_sc_hd__a22o_1
X_05318_ _05318_/A _05318_/B VGND VGND VPWR VPWR _05829_/A sky130_fd_sc_hd__or2_2
X_08106_ _07283_/Y _08067_/X _07208_/Y _08068_/X _08105_/X VGND VGND VPWR VPWR _08106_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08037_ _08038_/A _08037_/B _10006_/Q VGND VGND VPWR VPWR _08205_/A sky130_fd_sc_hd__or3_4
X_05249_ _05277_/A VGND VGND VPWR VPWR _05361_/B sky130_fd_sc_hd__buf_2
XFILLER_122_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09988_ _10006_/CLK _09988_/D repeater407/X VGND VGND VPWR VPWR _09988_/Q sky130_fd_sc_hd__dfstp_2
X_08939_ _08939_/A VGND VGND VPWR VPWR _09068_/B sky130_fd_sc_hd__inv_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10000_/CLK sky130_fd_sc_hd__clkbuf_16
X_10128_ _10238_/CLK _10128_/D repeater403/X VGND VGND VPWR VPWR _10128_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10127_/CLK sky130_fd_sc_hd__clkbuf_16
X_10059_ _10110_/CLK _10059_/D repeater405/X VGND VGND VPWR VPWR _10059_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07270_ _09962_/Q VGND VGND VPWR VPWR _07270_/Y sky130_fd_sc_hd__clkinv_2
X_06221_ _09988_/Q VGND VGND VPWR VPWR _06245_/B sky130_fd_sc_hd__inv_2
XFILLER_176_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06152_ _06337_/A VGND VGND VPWR VPWR _06313_/A sky130_fd_sc_hd__clkbuf_4
X_05103_ _05160_/A _05103_/B VGND VGND VPWR VPWR _06705_/A sky130_fd_sc_hd__or2_2
X_06083_ _10053_/Q _06080_/X _09658_/A1 _06081_/Y VGND VGND VPWR VPWR _10053_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09911_ _10006_/CLK _09911_/D repeater409/X VGND VGND VPWR VPWR _09911_/Q sky130_fd_sc_hd__dfrtp_1
X_05034_ _05034_/A VGND VGND VPWR VPWR _06679_/B sky130_fd_sc_hd__inv_2
XFILLER_171_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09842_ _10350_/CLK _09842_/D repeater404/X VGND VGND VPWR VPWR _09842_/Q sky130_fd_sc_hd__dfstp_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _10406_/CLK _09773_/D _06672_/X VGND VGND VPWR VPWR _09773_/Q sky130_fd_sc_hd__dfrtp_4
X_06985_ _06985_/A _06985_/B _06985_/C _06985_/D VGND VGND VPWR VPWR _07028_/B sky130_fd_sc_hd__and4_1
X_08724_ _08736_/A _08849_/B VGND VGND VPWR VPWR _09124_/A sky130_fd_sc_hd__or2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05936_ _10144_/Q _05929_/X _09550_/A0 _05931_/X VGND VGND VPWR VPWR _10144_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08786_/A _08788_/A VGND VGND VPWR VPWR _08676_/B sky130_fd_sc_hd__or2_1
X_05867_ _05867_/A VGND VGND VPWR VPWR _05867_/Y sky130_fd_sc_hd__inv_2
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07606_/A _07606_/B VGND VGND VPWR VPWR _07606_/X sky130_fd_sc_hd__or2_1
X_08586_ _08586_/A _08951_/B VGND VGND VPWR VPWR _09025_/A sky130_fd_sc_hd__or2_1
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04818_ _10299_/Q VGND VGND VPWR VPWR _04818_/Y sky130_fd_sc_hd__inv_2
X_07537_ _07612_/A _07612_/B _07562_/B VGND VGND VPWR VPWR _07787_/A sky130_fd_sc_hd__or3_1
X_05798_ _10226_/Q _05795_/X _09581_/X _05797_/X VGND VGND VPWR VPWR _10226_/D sky130_fd_sc_hd__a22o_1
XFILLER_169_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07468_ _10419_/Q VGND VGND VPWR VPWR _07468_/Y sky130_fd_sc_hd__inv_2
X_09207_ _09283_/B _09207_/B VGND VGND VPWR VPWR _09371_/A sky130_fd_sc_hd__or2_1
X_07399_ _07394_/Y _05549_/A _07395_/Y _05807_/A _07398_/X VGND VGND VPWR VPWR _07418_/A
+ sky130_fd_sc_hd__o221a_1
X_06419_ _06417_/X _09629_/X _09650_/X _09889_/Q VGND VGND VPWR VPWR _09889_/D sky130_fd_sc_hd__o22a_1
XFILLER_182_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09138_ _09138_/A _09271_/B VGND VGND VPWR VPWR _09139_/B sky130_fd_sc_hd__or2_1
XFILLER_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09069_ _09339_/B _09198_/B VGND VGND VPWR VPWR _09070_/D sky130_fd_sc_hd__or2_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput208 _09472_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput219 _09492_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_153_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06770_ _06770_/A VGND VGND VPWR VPWR _09699_/S sky130_fd_sc_hd__buf_12
XFILLER_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05721_ _10271_/Q _05717_/X _09548_/X _05718_/X VGND VGND VPWR VPWR _10271_/D sky130_fd_sc_hd__o22a_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05652_ _05652_/A VGND VGND VPWR VPWR _05654_/A sky130_fd_sc_hd__clkbuf_2
X_08440_ _09102_/C VGND VGND VPWR VPWR _08631_/A sky130_fd_sc_hd__inv_2
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08371_ _09788_/Q _08371_/B VGND VGND VPWR VPWR _08371_/X sky130_fd_sc_hd__and2_1
XFILLER_189_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05583_ _10347_/Q _05577_/X _09547_/A1 _05579_/X VGND VGND VPWR VPWR _10347_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07322_ _07320_/Y _05918_/B _07321_/Y _05838_/A VGND VGND VPWR VPWR _07322_/X sky130_fd_sc_hd__o22a_1
X_07253_ _09904_/Q VGND VGND VPWR VPWR _07253_/Y sky130_fd_sc_hd__inv_2
X_07184_ _10260_/Q VGND VGND VPWR VPWR _07184_/Y sky130_fd_sc_hd__inv_2
X_06204_ _07994_/B _09777_/Q _10002_/Q _06203_/Y VGND VGND VPWR VPWR _10002_/D sky130_fd_sc_hd__a22o_1
X_06135_ _07477_/A _06133_/Y _06227_/B _09776_/Q _09554_/X VGND VGND VPWR VPWR _06139_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06066_ _06108_/A _06066_/B VGND VGND VPWR VPWR _06068_/A sky130_fd_sc_hd__or2_2
X_05017_ _09674_/X _05109_/B _09670_/X _09668_/X VGND VGND VPWR VPWR _05198_/A sky130_fd_sc_hd__or4_2
X_09825_ _10405_/CLK _09825_/D hold41/X VGND VGND VPWR VPWR _09825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09756_ _09781_/CLK _09756_/D VGND VGND VPWR VPWR _09756_/Q sky130_fd_sc_hd__dfxtp_1
X_06968_ _10163_/Q VGND VGND VPWR VPWR _06968_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09687_ _08364_/X input190/X _09698_/S VGND VGND VPWR VPWR _09687_/X sky130_fd_sc_hd__mux2_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05919_ _05920_/A VGND VGND VPWR VPWR _05919_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08707_ _08710_/A _08824_/B VGND VGND VPWR VPWR _09158_/A sky130_fd_sc_hd__or2_1
XFILLER_100_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08638_ _08656_/A _08675_/B VGND VGND VPWR VPWR _08786_/B sky130_fd_sc_hd__or2_4
X_06899_ _10263_/Q VGND VGND VPWR VPWR _06899_/Y sky130_fd_sc_hd__inv_2
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08569_ _09180_/A _09225_/A VGND VGND VPWR VPWR _08570_/B sky130_fd_sc_hd__or2_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10462_ _10471_/CLK _10462_/D repeater409/X VGND VGND VPWR VPWR _10462_/Q sky130_fd_sc_hd__dfstp_1
X_10393_ _04811_/A1 _10393_/D _05465_/X VGND VGND VPWR VPWR _10393_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07940_ _07150_/Y _07777_/A _07061_/Y _07778_/A _07939_/X VGND VGND VPWR VPWR _07962_/A
+ sky130_fd_sc_hd__o221a_1
X_07871_ _07869_/Y _07799_/X _05251_/Y _07801_/X _07870_/X VGND VGND VPWR VPWR _07875_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09610_ _08310_/Y _10327_/Q _09700_/S VGND VGND VPWR VPWR _09610_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06822_ _10069_/Q VGND VGND VPWR VPWR _06822_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06753_ _10265_/Q VGND VGND VPWR VPWR _06753_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09541_ _10321_/Q _09579_/X _09679_/S VGND VGND VPWR VPWR _09541_/X sky130_fd_sc_hd__mux2_1
X_05704_ _10281_/Q _05701_/X _09542_/X _05702_/X VGND VGND VPWR VPWR _10281_/D sky130_fd_sc_hd__o22a_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09472_ _09472_/A VGND VGND VPWR VPWR _09472_/X sky130_fd_sc_hd__clkbuf_1
X_06684_ _09767_/Q _06681_/A _06684_/B1 _06681_/Y VGND VGND VPWR VPWR _09767_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08423_ _08634_/A VGND VGND VPWR VPWR _08537_/C sky130_fd_sc_hd__clkbuf_2
X_05635_ _10318_/Q _05628_/A _09660_/A1 _05629_/A VGND VGND VPWR VPWR _10318_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08354_ _08354_/A _08354_/B _09790_/Q VGND VGND VPWR VPWR _08354_/X sky130_fd_sc_hd__and3_1
X_05566_ _06630_/C VGND VGND VPWR VPWR _05775_/A sky130_fd_sc_hd__buf_4
XFILLER_177_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07305_ _10431_/Q _05030_/Y _10330_/Q _05151_/X _07304_/X VGND VGND VPWR VPWR _07324_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05497_ _05497_/A VGND VGND VPWR VPWR _05498_/A sky130_fd_sc_hd__clkbuf_1
X_08285_ _07272_/Y _08201_/X _07923_/Y _08202_/X VGND VGND VPWR VPWR _08285_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07236_ _07231_/Y _05910_/B _07232_/Y _06153_/A _07235_/X VGND VGND VPWR VPWR _07243_/C
+ sky130_fd_sc_hd__o221a_1
X_07167_ _07167_/A _07167_/B _07167_/C VGND VGND VPWR VPWR _07289_/A sky130_fd_sc_hd__or3_2
X_06118_ _10030_/Q _06110_/A _06684_/B1 _06111_/A VGND VGND VPWR VPWR _10030_/D sky130_fd_sc_hd__a22o_1
X_07098_ _10105_/Q VGND VGND VPWR VPWR _07098_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06049_ _10074_/Q _06046_/X _09658_/A1 _06047_/Y VGND VGND VPWR VPWR _10074_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09808_ _09572_/A1 _09808_/D _06592_/X VGND VGND VPWR VPWR _09808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09739_ _09781_/CLK _09739_/D VGND VGND VPWR VPWR _09739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10445_ _10487_/CLK _10445_/D _05034_/A VGND VGND VPWR VPWR _10445_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10376_ _10404_/CLK _10376_/D hold41/X VGND VGND VPWR VPWR _10376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _10509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05420_ _05421_/A VGND VGND VPWR VPWR _05420_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_181 input79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _07781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05351_ _05351_/A _05359_/B VGND VGND VPWR VPWR _06493_/A sky130_fd_sc_hd__or2_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05282_ _10496_/Q VGND VGND VPWR VPWR _05282_/Y sky130_fd_sc_hd__inv_2
X_08070_ _08189_/A VGND VGND VPWR VPWR _08070_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07021_ _10016_/Q VGND VGND VPWR VPWR _07021_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08972_ _08972_/A _08974_/B _09005_/A VGND VGND VPWR VPWR _09405_/B sky130_fd_sc_hd__nor3_1
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold29 hold29/A VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _10339_/Q VGND VGND VPWR VPWR _07923_/Y sky130_fd_sc_hd__inv_2
X_07854_ _07854_/A _07932_/B VGND VGND VPWR VPWR _07854_/X sky130_fd_sc_hd__or2_1
XFILLER_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06805_ _10173_/Q VGND VGND VPWR VPWR _06805_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07785_ _06796_/Y _07779_/X _07780_/Y _07781_/X _07784_/X VGND VGND VPWR VPWR _07785_/X
+ sky130_fd_sc_hd__o221a_1
X_04997_ _10450_/Q _04994_/X _09581_/X _04996_/X VGND VGND VPWR VPWR _10450_/D sky130_fd_sc_hd__a22o_1
X_09524_ _09524_/A VGND VGND VPWR VPWR _09524_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06736_ _10192_/Q VGND VGND VPWR VPWR _06736_/Y sky130_fd_sc_hd__clkinv_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06667_ _06667_/A VGND VGND VPWR VPWR _06667_/X sky130_fd_sc_hd__clkbuf_1
X_09455_ _09455_/A VGND VGND VPWR VPWR _09456_/A sky130_fd_sc_hd__clkbuf_1
X_08406_ _08426_/A _08406_/B _08406_/C _08406_/D VGND VGND VPWR VPWR _08641_/C sky130_fd_sc_hd__or4_1
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05618_ _10328_/Q _05616_/X _09545_/A1 _05617_/Y VGND VGND VPWR VPWR _10328_/D sky130_fd_sc_hd__a22o_1
X_09386_ _09386_/A _09386_/B VGND VGND VPWR VPWR _09387_/B sky130_fd_sc_hd__or2_1
X_06598_ _06593_/A _06593_/B _06593_/Y VGND VGND VPWR VPWR _09807_/D sky130_fd_sc_hd__a21oi_1
XFILLER_177_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05549_ _05549_/A VGND VGND VPWR VPWR _05550_/B sky130_fd_sc_hd__buf_4
X_08337_ _08338_/B _08337_/B VGND VGND VPWR VPWR _08337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08268_ _07368_/Y _08199_/X _07397_/Y _08200_/X _08267_/X VGND VGND VPWR VPWR _08273_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07219_ _09949_/Q VGND VGND VPWR VPWR _07219_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _10355_/CLK _10230_/D repeater406/X VGND VGND VPWR VPWR _10230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08199_ _08199_/A VGND VGND VPWR VPWR _08199_/X sky130_fd_sc_hd__buf_2
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput380 _09738_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_2
X_10161_ _10353_/CLK _10161_/D repeater403/X VGND VGND VPWR VPWR _10161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10092_ _10289_/CLK _10092_/D repeater402/X VGND VGND VPWR VPWR _10092_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput391 _09743_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10428_ net399_2/A _10428_/D _05045_/X VGND VGND VPWR VPWR _10428_/Q sky130_fd_sc_hd__dfrtn_1
X_10359_ _10364_/CLK _10359_/D repeater410/X VGND VGND VPWR VPWR _10359_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_04920_ _09788_/Q _09789_/Q _09790_/Q VGND VGND VPWR VPWR _08356_/A sky130_fd_sc_hd__or3_4
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04851_ _04851_/A VGND VGND VPWR VPWR _04851_/X sky130_fd_sc_hd__clkbuf_2
X_07570_ _07585_/C _07612_/A _07601_/A VGND VGND VPWR VPWR _07777_/A sky130_fd_sc_hd__or3_4
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06521_ _09839_/Q _06517_/X _09580_/X _06519_/X VGND VGND VPWR VPWR _09839_/D sky130_fd_sc_hd__a22o_1
X_09240_ _09319_/A _09240_/B _09446_/D _09326_/D VGND VGND VPWR VPWR _09244_/A sky130_fd_sc_hd__or4_1
X_06452_ _06452_/A VGND VGND VPWR VPWR _06452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05403_ _05406_/A VGND VGND VPWR VPWR _05404_/A sky130_fd_sc_hd__clkbuf_1
X_09171_ _09171_/A _09397_/A VGND VGND VPWR VPWR _09172_/D sky130_fd_sc_hd__or2_1
X_06383_ _06380_/X _09599_/X _09650_/X _09912_/Q VGND VGND VPWR VPWR _09912_/D sky130_fd_sc_hd__o22a_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05334_ _05334_/A VGND VGND VPWR VPWR _05567_/B sky130_fd_sc_hd__clkbuf_4
X_08122_ _09513_/A _08065_/X _09483_/A _06188_/X VGND VGND VPWR VPWR _08122_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08053_ _08220_/A VGND VGND VPWR VPWR _08053_/X sky130_fd_sc_hd__clkbuf_2
X_07004_ _09932_/Q VGND VGND VPWR VPWR _07004_/Y sky130_fd_sc_hd__clkinv_4
X_05265_ _10037_/Q VGND VGND VPWR VPWR _05265_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_162_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05196_ _05184_/Y _05927_/A _05186_/Y _05785_/B _05195_/X VGND VGND VPWR VPWR _05236_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _08972_/A _08959_/B VGND VGND VPWR VPWR _09073_/B sky130_fd_sc_hd__nor2_1
Xinput108 sram_ro_data[23] VGND VGND VPWR VPWR input108/X sky130_fd_sc_hd__buf_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07906_ _07345_/Y _07816_/X _07337_/Y _07817_/X _07905_/X VGND VGND VPWR VPWR _07911_/B
+ sky130_fd_sc_hd__o221a_1
Xinput119 sram_ro_data[4] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08886_ _09051_/A VGND VGND VPWR VPWR _09295_/B sky130_fd_sc_hd__inv_2
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07837_ _06719_/Y _07777_/X _06745_/Y _07778_/X _07836_/X VGND VGND VPWR VPWR _07860_/A
+ sky130_fd_sc_hd__o221a_1
X_07768_ _07768_/A VGND VGND VPWR VPWR _07768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09507_ _09507_/A VGND VGND VPWR VPWR _09508_/A sky130_fd_sc_hd__clkbuf_1
X_06719_ _10244_/Q VGND VGND VPWR VPWR _06719_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07699_ _09457_/A _07533_/C _09463_/A _07629_/X VGND VGND VPWR VPWR _07699_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09438_ _08766_/A _08581_/B _08939_/A _09018_/X _09212_/C VGND VGND VPWR VPWR _09439_/B
+ sky130_fd_sc_hd__o2111ai_4
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _09369_/A _09369_/B _09369_/C _09369_/D VGND VGND VPWR VPWR _09408_/C sky130_fd_sc_hd__or4_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_92 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 _09555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_81 _07502_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10213_ _10244_/CLK _10213_/D repeater402/X VGND VGND VPWR VPWR _10213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10144_ _10491_/CLK _10144_/D repeater403/X VGND VGND VPWR VPWR _10144_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10075_ _10512_/CLK _10075_/D _07492_/B VGND VGND VPWR VPWR _10075_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05050_ _05053_/A VGND VGND VPWR VPWR _05051_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _05993_/A _05952_/B VGND VGND VPWR VPWR _05954_/A sky130_fd_sc_hd__or2_1
X_08740_ _08862_/A VGND VGND VPWR VPWR _08860_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05883_ _05896_/A _05883_/B VGND VGND VPWR VPWR _05885_/A sky130_fd_sc_hd__or2_2
X_08671_ _08836_/B VGND VGND VPWR VPWR _09260_/A sky130_fd_sc_hd__clkbuf_2
X_04903_ _04903_/A VGND VGND VPWR VPWR _04904_/A sky130_fd_sc_hd__inv_2
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07622_ _07782_/A VGND VGND VPWR VPWR _07622_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_04834_ _05149_/A _05178_/A VGND VGND VPWR VPWR _04836_/B sky130_fd_sc_hd__or2_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07553_ _07642_/A _07639_/A _07629_/A _07600_/A VGND VGND VPWR VPWR _07567_/B sky130_fd_sc_hd__and4_1
X_06504_ _06505_/A VGND VGND VPWR VPWR _06504_/X sky130_fd_sc_hd__clkbuf_2
X_07484_ _05395_/A _07489_/A _07489_/B _05390_/X _07483_/X VGND VGND VPWR VPWR _07485_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06435_ _09878_/Q _06431_/X _06683_/B1 _06432_/Y VGND VGND VPWR VPWR _09878_/D sky130_fd_sc_hd__a22o_1
X_09223_ _09223_/A _09223_/B VGND VGND VPWR VPWR _09415_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09154_ _09010_/A _09012_/A _08693_/X _09153_/X _08697_/X VGND VGND VPWR VPWR _09156_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_182_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06366_ _09925_/Q _06361_/X _09579_/X _06363_/X VGND VGND VPWR VPWR _09925_/D sky130_fd_sc_hd__a22o_1
X_08105_ _07201_/Y _08069_/X _07226_/Y _08070_/X VGND VGND VPWR VPWR _08105_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09085_ _08897_/A _09085_/B _09085_/C _09085_/D VGND VGND VPWR VPWR _09297_/A sky130_fd_sc_hd__and4b_1
X_06297_ _09965_/Q _06292_/X _09579_/X _06294_/X VGND VGND VPWR VPWR _09965_/D sky130_fd_sc_hd__a22o_1
X_05317_ _10201_/Q VGND VGND VPWR VPWR _05317_/Y sky130_fd_sc_hd__clkinv_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_2
XFILLER_135_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ _05225_/Y _08199_/A _05134_/Y _08200_/A _08035_/X VGND VGND VPWR VPWR _08049_/B
+ sky130_fd_sc_hd__o221a_1
X_05248_ _09820_/Q VGND VGND VPWR VPWR _05248_/Y sky130_fd_sc_hd__inv_4
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05179_ _05179_/A VGND VGND VPWR VPWR _05179_/Y sky130_fd_sc_hd__inv_2
X_09987_ _10288_/CLK _09987_/D repeater406/X VGND VGND VPWR VPWR _09987_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08938_ _08938_/A _08942_/B VGND VGND VPWR VPWR _08939_/A sky130_fd_sc_hd__or2_2
X_08869_ _08869_/A _08869_/B VGND VGND VPWR VPWR _08869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10127_ _10127_/CLK _10127_/D _07492_/B VGND VGND VPWR VPWR _10127_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10058_ _10110_/CLK _10058_/D repeater405/X VGND VGND VPWR VPWR _10058_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06220_ _09989_/Q VGND VGND VPWR VPWR _06243_/A sky130_fd_sc_hd__inv_2
XFILLER_191_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06151_ _06137_/A _06150_/A _10020_/Q _06150_/Y _06142_/X VGND VGND VPWR VPWR _10020_/D
+ sky130_fd_sc_hd__o221a_1
X_05102_ _10133_/Q VGND VGND VPWR VPWR _05102_/Y sky130_fd_sc_hd__clkinv_2
X_06082_ _10054_/Q _06080_/X _09545_/A1 _06081_/Y VGND VGND VPWR VPWR _10054_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09910_ _10006_/CLK _09910_/D repeater409/X VGND VGND VPWR VPWR _09910_/Q sky130_fd_sc_hd__dfrtp_1
X_05033_ _09678_/X _05030_/Y _09536_/A3 _10430_/Q _05031_/X VGND VGND VPWR VPWR _10430_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_171_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09841_ _10350_/CLK _09841_/D repeater404/X VGND VGND VPWR VPWR _09841_/Q sky130_fd_sc_hd__dfstp_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06984_ _06979_/Y _06438_/A _06980_/Y _06312_/A _06983_/X VGND VGND VPWR VPWR _06985_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09572_/A1 _09772_/D _06674_/X VGND VGND VPWR VPWR _09772_/Q sky130_fd_sc_hd__dfrtp_4
X_05935_ _10145_/Q _05929_/X _09547_/A1 _05931_/X VGND VGND VPWR VPWR _10145_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08723_ _09253_/A _08665_/Y _08722_/Y VGND VGND VPWR VPWR _08725_/A sky130_fd_sc_hd__a21oi_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _08668_/A VGND VGND VPWR VPWR _08788_/A sky130_fd_sc_hd__clkbuf_2
X_05866_ _05867_/A VGND VGND VPWR VPWR _05866_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08585_/A _08951_/B VGND VGND VPWR VPWR _09200_/A sky130_fd_sc_hd__or2_1
X_04817_ _09672_/X VGND VGND VPWR VPWR _05201_/C sky130_fd_sc_hd__inv_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07605_ _05324_/Y _07816_/A _05265_/Y _07817_/A _07604_/X VGND VGND VPWR VPWR _07615_/B
+ sky130_fd_sc_hd__o221a_1
X_05797_ _05797_/A VGND VGND VPWR VPWR _05797_/X sky130_fd_sc_hd__clkbuf_2
X_07536_ _07602_/C VGND VGND VPWR VPWR _07612_/B sky130_fd_sc_hd__clkbuf_1
X_07467_ _09535_/A _09531_/A _07425_/B VGND VGND VPWR VPWR _09790_/D sky130_fd_sc_hd__o21ai_1
X_09206_ _09206_/A _09206_/B VGND VGND VPWR VPWR _09407_/A sky130_fd_sc_hd__nor2_1
X_07398_ _07396_/Y _05761_/A _07397_/Y _05993_/B VGND VGND VPWR VPWR _07398_/X sky130_fd_sc_hd__o22a_1
X_06418_ _06417_/X _09631_/X _09650_/X _09890_/Q VGND VGND VPWR VPWR _09890_/D sky130_fd_sc_hd__o22a_1
X_09137_ _09137_/A _09297_/B VGND VGND VPWR VPWR _09271_/B sky130_fd_sc_hd__or2_1
X_06349_ _09934_/Q _06341_/A _09661_/A1 _06342_/A VGND VGND VPWR VPWR _09934_/D sky130_fd_sc_hd__a22o_1
X_09068_ _09068_/A _09068_/B VGND VGND VPWR VPWR _09287_/C sky130_fd_sc_hd__or2_1
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08019_ _08037_/B _08019_/B _08019_/C VGND VGND VPWR VPWR _08187_/A sky130_fd_sc_hd__or3_4
XFILLER_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput209 _09474_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_114_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05720_ _10272_/Q _05717_/X _09587_/X _05718_/X VGND VGND VPWR VPWR _10272_/D sky130_fd_sc_hd__o22a_1
XFILLER_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05651_ _05651_/A _05651_/B _09677_/S VGND VGND VPWR VPWR _05652_/A sky130_fd_sc_hd__or3_4
X_08370_ _09790_/Q input188/X _09789_/Q input170/X _08369_/X VGND VGND VPWR VPWR _08370_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ _10194_/Q VGND VGND VPWR VPWR _07321_/Y sky130_fd_sc_hd__clkinv_4
X_05582_ _10348_/Q _05577_/X _09579_/X _05579_/X VGND VGND VPWR VPWR _10348_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07252_ _09896_/Q VGND VGND VPWR VPWR _07252_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_117_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06203_ _06203_/A VGND VGND VPWR VPWR _06203_/Y sky130_fd_sc_hd__inv_2
X_07183_ _10221_/Q VGND VGND VPWR VPWR _07183_/Y sky130_fd_sc_hd__inv_2
X_06134_ _09777_/Q VGND VGND VPWR VPWR _06227_/B sky130_fd_sc_hd__clkinv_2
XFILLER_144_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06065_ _10063_/Q _06056_/A _09659_/A1 _06057_/A VGND VGND VPWR VPWR _10063_/D sky130_fd_sc_hd__a22o_1
X_05016_ _10437_/Q _05009_/A _09536_/A3 _05010_/A VGND VGND VPWR VPWR _10437_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09824_ _10405_/CLK _09824_/D hold41/X VGND VGND VPWR VPWR _09824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09755_ _09781_/CLK _09755_/D VGND VGND VPWR VPWR _09755_/Q sky130_fd_sc_hd__dfxtp_1
X_06967_ _10171_/Q VGND VGND VPWR VPWR _06967_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_104_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09686_ _08362_/X input187/X _09698_/S VGND VGND VPWR VPWR _09686_/X sky130_fd_sc_hd__mux2_1
X_06898_ _10198_/Q VGND VGND VPWR VPWR _06898_/Y sky130_fd_sc_hd__inv_4
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05918_ _05993_/A _05918_/B VGND VGND VPWR VPWR _05920_/A sky130_fd_sc_hd__or2_1
XFILLER_104_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08706_ _08717_/A _08824_/B VGND VGND VPWR VPWR _09111_/A sky130_fd_sc_hd__or2_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08637_ _09236_/A _08635_/Y _08556_/D _08888_/B VGND VGND VPWR VPWR _08675_/B sky130_fd_sc_hd__o22a_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ _10194_/Q _05841_/A _09661_/A1 _05842_/A VGND VGND VPWR VPWR _10194_/D sky130_fd_sc_hd__a22o_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08568_ _08568_/A _09236_/B VGND VGND VPWR VPWR _09225_/A sky130_fd_sc_hd__or2b_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _10350_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08499_ _08585_/A VGND VGND VPWR VPWR _08620_/A sky130_fd_sc_hd__buf_2
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07519_ _07519_/A VGND VGND VPWR VPWR _07533_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10461_ _10486_/CLK _10461_/D repeater409/X VGND VGND VPWR VPWR _10461_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10512_/CLK sky130_fd_sc_hd__clkbuf_16
X_10392_ _04811_/A1 _10392_/D _05468_/X VGND VGND VPWR VPWR _10392_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_77_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07870_ _05287_/Y _07755_/X _05232_/Y _07802_/X VGND VGND VPWR VPWR _07870_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06821_ _10147_/Q VGND VGND VPWR VPWR _06821_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09540_ input66/X VGND VGND VPWR VPWR _09540_/X sky130_fd_sc_hd__clkbuf_1
X_06752_ _10174_/Q VGND VGND VPWR VPWR _06752_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09471_ _09471_/A VGND VGND VPWR VPWR _09472_/A sky130_fd_sc_hd__clkbuf_1
X_05703_ _10282_/Q _05701_/X _09543_/X _05702_/X VGND VGND VPWR VPWR _10282_/D sky130_fd_sc_hd__o22a_1
X_08422_ _08424_/B VGND VGND VPWR VPWR _08476_/A sky130_fd_sc_hd__inv_2
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06683_ _09768_/Q _06681_/A _06683_/B1 _06681_/Y VGND VGND VPWR VPWR _09768_/D sky130_fd_sc_hd__a22o_1
X_05634_ _10319_/Q _05627_/X _09658_/A1 _05629_/X VGND VGND VPWR VPWR _10319_/D sky130_fd_sc_hd__a22o_1
X_08353_ _08353_/A _08354_/A _09788_/Q VGND VGND VPWR VPWR _08353_/X sky130_fd_sc_hd__and3_1
X_05565_ _10356_/Q _05564_/X _04923_/Y VGND VGND VPWR VPWR _10356_/D sky130_fd_sc_hd__o21a_1
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08284_ _07258_/Y _08193_/X _07265_/Y _08194_/X _08283_/X VGND VGND VPWR VPWR _08291_/A
+ sky130_fd_sc_hd__o221a_1
X_07304_ _10509_/Q _04822_/Y _10468_/Q _04959_/Y VGND VGND VPWR VPWR _07304_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05496_ _05496_/A VGND VGND VPWR VPWR _10385_/D sky130_fd_sc_hd__clkbuf_1
X_07235_ _07233_/Y _06205_/A _07234_/Y _06529_/B VGND VGND VPWR VPWR _07235_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07166_ input102/X _05153_/X _10331_/Q _05151_/X _07165_/X VGND VGND VPWR VPWR _07167_/C
+ sky130_fd_sc_hd__a221o_1
X_06117_ _10031_/Q _06110_/A _06683_/B1 _06111_/A VGND VGND VPWR VPWR _10031_/D sky130_fd_sc_hd__a22o_1
X_07097_ _10204_/Q VGND VGND VPWR VPWR _07097_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06048_ _10075_/Q _06046_/X _09545_/A1 _06047_/Y VGND VGND VPWR VPWR _10075_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07999_ _08032_/A _08044_/B _10006_/Q VGND VGND VPWR VPWR _08220_/A sky130_fd_sc_hd__or3_4
X_09807_ _10406_/CLK _09807_/D _06597_/X VGND VGND VPWR VPWR _09807_/Q sky130_fd_sc_hd__dfrtp_2
X_09738_ _09781_/CLK _09738_/D VGND VGND VPWR VPWR _09738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09669_ _09802_/Q _09801_/Q _09773_/Q VGND VGND VPWR VPWR _09669_/X sky130_fd_sc_hd__mux2_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ _10513_/CLK _10513_/D _07492_/B VGND VGND VPWR VPWR _10513_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10444_ _10486_/CLK _10444_/D _05034_/A VGND VGND VPWR VPWR _10444_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10375_ _10404_/CLK _10375_/D repeater410/X VGND VGND VPWR VPWR _10375_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _07098_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _04807_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _07781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05350_ _09849_/Q VGND VGND VPWR VPWR _05350_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05281_ _05281_/A _05281_/B _05281_/C _05281_/D VGND VGND VPWR VPWR _05365_/B sky130_fd_sc_hd__and4_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07020_ _07015_/Y _06393_/B _07016_/Y _05434_/B _07019_/X VGND VGND VPWR VPWR _07027_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08971_ _08971_/A _09427_/B VGND VGND VPWR VPWR _08973_/A sky130_fd_sc_hd__or2_1
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07922_ _07176_/Y _07799_/X _07275_/Y _07801_/X _07921_/X VGND VGND VPWR VPWR _07926_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold19 hold19/A VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _06741_/Y _07816_/X _06717_/Y _07817_/X _07852_/X VGND VGND VPWR VPWR _07859_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06804_ _09847_/Q VGND VGND VPWR VPWR _06804_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07784_ _06823_/Y _07782_/X _06817_/Y _07783_/X VGND VGND VPWR VPWR _07784_/X sky130_fd_sc_hd__o22a_1
X_04996_ _04996_/A VGND VGND VPWR VPWR _04996_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09523_ input63/X input79/X VGND VGND VPWR VPWR _09524_/A sky130_fd_sc_hd__and2_1
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06735_ _09927_/Q VGND VGND VPWR VPWR _06735_/Y sky130_fd_sc_hd__clkinv_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09454_ _09441_/Y _09435_/Y _09443_/X _09453_/X VGND VGND VPWR VPWR _09454_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06666_ _06666_/A VGND VGND VPWR VPWR _06667_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08405_ _08634_/A _08417_/A _08405_/C _08405_/D VGND VGND VPWR VPWR _08406_/D sky130_fd_sc_hd__nand4bb_1
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09385_ _09385_/A _09418_/A _09385_/C _09419_/B VGND VGND VPWR VPWR _09385_/X sky130_fd_sc_hd__or4_1
X_05617_ _05617_/A VGND VGND VPWR VPWR _05617_/Y sky130_fd_sc_hd__inv_2
X_06597_ _06597_/A VGND VGND VPWR VPWR _06597_/X sky130_fd_sc_hd__clkbuf_1
X_08336_ _09801_/Q _08335_/B _09802_/Q VGND VGND VPWR VPWR _08337_/B sky130_fd_sc_hd__a21oi_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05548_ _10365_/Q _05542_/X _09536_/A3 _05543_/Y VGND VGND VPWR VPWR _10365_/D sky130_fd_sc_hd__a22o_1
XFILLER_165_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08267_ _07318_/Y _08201_/X _07898_/Y _08202_/X VGND VGND VPWR VPWR _08267_/X sky130_fd_sc_hd__o22a_1
X_05479_ _10388_/Q _05475_/X _06683_/B1 _05476_/Y VGND VGND VPWR VPWR _10388_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08198_ _06799_/Y _08193_/X _06818_/Y _08194_/X _08197_/X VGND VGND VPWR VPWR _08217_/A
+ sky130_fd_sc_hd__o221a_1
X_07218_ _07218_/A _07218_/B _07218_/C _07218_/D VGND VGND VPWR VPWR _07288_/A sky130_fd_sc_hd__and4_1
X_07149_ _09455_/A _05527_/A _09461_/A _06538_/B _07148_/X VGND VGND VPWR VPWR _07156_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _10353_/CLK _10160_/D repeater403/X VGND VGND VPWR VPWR _10160_/Q sky130_fd_sc_hd__dfstp_1
Xoutput370 _09753_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10091_ _10289_/CLK _10091_/D repeater402/X VGND VGND VPWR VPWR _10091_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput381 _09739_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10427_ net399_2/A _10427_/D _05048_/X VGND VGND VPWR VPWR _10427_/Q sky130_fd_sc_hd__dfrtn_1
X_10358_ _10364_/CLK _10358_/D repeater410/X VGND VGND VPWR VPWR _10358_/Q sky130_fd_sc_hd__dfstp_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10289_/CLK _10289_/D repeater402/X VGND VGND VPWR VPWR _10289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04850_ _04852_/A VGND VGND VPWR VPWR _04851_/A sky130_fd_sc_hd__inv_2
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06520_ _09840_/Q _06517_/X _09581_/X _06519_/X VGND VGND VPWR VPWR _09840_/D sky130_fd_sc_hd__a22o_1
X_06451_ _06644_/A VGND VGND VPWR VPWR _06452_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05402_ _10417_/Q _05396_/X _10416_/Q _05398_/X VGND VGND VPWR VPWR _10417_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06382_ _06380_/X _09601_/X _09650_/X _09913_/Q VGND VGND VPWR VPWR _09913_/D sky130_fd_sc_hd__o22a_1
X_09170_ _08491_/B _08999_/B _08527_/Y _09253_/A _08665_/Y VGND VGND VPWR VPWR _09380_/A
+ sky130_fd_sc_hd__a32o_1
X_05333_ _05333_/A _05359_/B VGND VGND VPWR VPWR _05334_/A sky130_fd_sc_hd__or2_1
X_08121_ _09473_/A _08058_/X _09461_/A _08059_/X _08120_/X VGND VGND VPWR VPWR _08135_/B
+ sky130_fd_sc_hd__o221a_1
X_05264_ _05305_/A _05284_/B VGND VGND VPWR VPWR _05727_/A sky130_fd_sc_hd__or2_4
X_08052_ _08219_/A VGND VGND VPWR VPWR _08052_/X sky130_fd_sc_hd__clkbuf_2
X_07003_ _10197_/Q VGND VGND VPWR VPWR _07003_/Y sky130_fd_sc_hd__inv_4
X_05195_ _05189_/Y _05851_/A _05192_/Y _06036_/A VGND VGND VPWR VPWR _05195_/X sky130_fd_sc_hd__o22a_1
XFILLER_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput109 sram_ro_data[24] VGND VGND VPWR VPWR input109/X sky130_fd_sc_hd__buf_2
X_08954_ _08954_/A _09386_/B VGND VGND VPWR VPWR _08956_/A sky130_fd_sc_hd__or2_1
XFILLER_69_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07905_ _07358_/Y _07818_/X _07904_/Y _07819_/X VGND VGND VPWR VPWR _07905_/X sky130_fd_sc_hd__o22a_1
X_08885_ _08884_/A _08908_/A _08884_/Y VGND VGND VPWR VPWR _09051_/A sky130_fd_sc_hd__a21oi_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07836_ _06748_/Y _07779_/X _07834_/Y _07781_/X _07835_/X VGND VGND VPWR VPWR _07836_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04979_ _04993_/A _05088_/A VGND VGND VPWR VPWR _04981_/A sky130_fd_sc_hd__or2_2
X_07767_ _06852_/Y _07656_/X _06891_/Y _07657_/X _07766_/X VGND VGND VPWR VPWR _07775_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09506_ _09506_/A VGND VGND VPWR VPWR _09506_/X sky130_fd_sc_hd__clkbuf_1
X_06718_ _10122_/Q VGND VGND VPWR VPWR _06718_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07698_ _09509_/A _07618_/X _09511_/A _07619_/X _07697_/X VGND VGND VPWR VPWR _07717_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06649_ _06655_/A VGND VGND VPWR VPWR _06650_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09437_ _09414_/Y _09445_/A _09424_/Y _09451_/A _09436_/Y VGND VGND VPWR VPWR _09437_/Y
+ sky130_fd_sc_hd__o221ai_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _08491_/B _08527_/Y _09226_/A _09073_/B VGND VGND VPWR VPWR _09369_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09299_ _09299_/A _09318_/B VGND VGND VPWR VPWR _09393_/A sky130_fd_sc_hd__or2_1
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08319_ _07006_/Y _08195_/A _06986_/Y _08196_/A VGND VGND VPWR VPWR _08319_/X sky130_fd_sc_hd__o22a_1
XANTENNA_60 input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _07502_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_71 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10212_ _10491_/CLK _10212_/D repeater403/X VGND VGND VPWR VPWR _10212_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10143_ _10238_/CLK _10143_/D repeater403/X VGND VGND VPWR VPWR _10143_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10074_ _10512_/CLK _10074_/D _07492_/B VGND VGND VPWR VPWR _10074_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05951_ _10133_/Q _05942_/A _09536_/A3 _05943_/A VGND VGND VPWR VPWR _10133_/D sky130_fd_sc_hd__a22o_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05882_ _05882_/A VGND VGND VPWR VPWR _05883_/B sky130_fd_sc_hd__clkbuf_4
X_08670_ _08835_/A VGND VGND VPWR VPWR _08836_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_04902_ _04903_/A VGND VGND VPWR VPWR _04902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_9_0_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_9_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_07621_ _07781_/A VGND VGND VPWR VPWR _07621_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04833_ _09674_/X _09676_/X _05027_/A _05109_/D VGND VGND VPWR VPWR _05178_/A sky130_fd_sc_hd__or4_2
XFILLER_81_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07552_ _07564_/C _07575_/B VGND VGND VPWR VPWR _07600_/A sky130_fd_sc_hd__or2_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06503_ _06538_/A _06503_/B VGND VGND VPWR VPWR _06505_/A sky130_fd_sc_hd__or2_2
XFILLER_179_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07483_ _05671_/B _05389_/Y _07483_/C _09681_/X VGND VGND VPWR VPWR _07483_/X sky130_fd_sc_hd__and4bb_1
X_09222_ _09222_/A _09222_/B _09222_/C VGND VGND VPWR VPWR _09317_/B sky130_fd_sc_hd__or3_1
X_06434_ _09879_/Q _06431_/X _09577_/X _06432_/Y VGND VGND VPWR VPWR _09879_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09153_ _08970_/A _08586_/A _08851_/A _09233_/C _08775_/A VGND VGND VPWR VPWR _09153_/X
+ sky130_fd_sc_hd__a311o_1
X_06365_ _09926_/Q _06361_/X _09580_/X _06363_/X VGND VGND VPWR VPWR _09926_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05316_ _05351_/A _05316_/B VGND VGND VPWR VPWR _05864_/A sky130_fd_sc_hd__or2_1
X_08104_ _07225_/Y _08065_/X _07233_/Y _06188_/X VGND VGND VPWR VPWR _08104_/X sky130_fd_sc_hd__o22a_1
X_09084_ _09276_/A _09084_/B VGND VGND VPWR VPWR _09432_/C sky130_fd_sc_hd__nor2_1
X_06296_ _09966_/Q _06292_/X _09580_/X _06294_/X VGND VGND VPWR VPWR _09966_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_4
X_05247_ _05237_/Y _06338_/A _05239_/Y _05575_/A _05246_/X VGND VGND VPWR VPWR _05281_/A
+ sky130_fd_sc_hd__o221a_2
X_08035_ _05241_/Y _08201_/A _05239_/Y _08202_/A VGND VGND VPWR VPWR _08035_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05178_ _05178_/A VGND VGND VPWR VPWR _05336_/A sky130_fd_sc_hd__buf_2
XFILLER_103_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09986_ _10288_/CLK _09986_/D repeater406/X VGND VGND VPWR VPWR _09986_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08937_ _08937_/A _09286_/B _09067_/B _09442_/B VGND VGND VPWR VPWR _08941_/A sky130_fd_sc_hd__or4_1
X_08868_ _09082_/A _08868_/B VGND VGND VPWR VPWR _08869_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07819_ _07819_/A VGND VGND VPWR VPWR _07819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08799_ _08913_/A _08895_/B _08913_/C VGND VGND VPWR VPWR _09057_/A sky130_fd_sc_hd__or3_4
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10126_ _10127_/CLK _10126_/D _07492_/B VGND VGND VPWR VPWR _10126_/Q sky130_fd_sc_hd__dfrtp_1
X_10057_ _10482_/CLK _10057_/D repeater405/X VGND VGND VPWR VPWR _10057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06150_ _06150_/A VGND VGND VPWR VPWR _06150_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05101_ _05101_/A VGND VGND VPWR VPWR _05101_/X sky130_fd_sc_hd__clkbuf_2
X_06081_ _06081_/A VGND VGND VPWR VPWR _06081_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05032_ _09678_/X _05030_/Y _06684_/B1 _10431_/Q _05031_/X VGND VGND VPWR VPWR _10431_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _10364_/CLK _09840_/D repeater410/X VGND VGND VPWR VPWR _09840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06983_ _06981_/Y _05748_/A _06982_/Y _05347_/A VGND VGND VPWR VPWR _06983_/X sky130_fd_sc_hd__o22a_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _10406_/CLK _09771_/D _06676_/X VGND VGND VPWR VPWR _09771_/Q sky130_fd_sc_hd__dfrtp_1
X_05934_ _10146_/Q _05929_/X _09579_/X _05931_/X VGND VGND VPWR VPWR _10146_/D sky130_fd_sc_hd__a22o_1
X_08722_ _08743_/A _09262_/A _08721_/X VGND VGND VPWR VPWR _08722_/Y sky130_fd_sc_hd__o21ai_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _08781_/B _08667_/A VGND VGND VPWR VPWR _08786_/A sky130_fd_sc_hd__nand2_4
X_05865_ _05874_/A _05865_/B VGND VGND VPWR VPWR _05867_/A sky130_fd_sc_hd__or2_1
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _09446_/A _08584_/B _09021_/A _09309_/A VGND VGND VPWR VPWR _08584_/Y sky130_fd_sc_hd__nor4_1
X_04816_ _04991_/A _09668_/X _05005_/C _04963_/B VGND VGND VPWR VPWR _05318_/A sky130_fd_sc_hd__or4_2
X_07604_ _05294_/Y _07818_/A _07603_/Y _07659_/A VGND VGND VPWR VPWR _07604_/X sky130_fd_sc_hd__o22a_1
X_05796_ _05796_/A VGND VGND VPWR VPWR _05797_/A sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07535_ _07606_/B VGND VGND VPWR VPWR _07983_/B sky130_fd_sc_hd__clkbuf_2
X_07466_ _09534_/A _09531_/A _06761_/B VGND VGND VPWR VPWR _09789_/D sky130_fd_sc_hd__o21ai_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09205_ _09205_/A _09103_/X VGND VGND VPWR VPWR _09209_/C sky130_fd_sc_hd__or2b_1
X_06417_ _06417_/A VGND VGND VPWR VPWR _06417_/X sky130_fd_sc_hd__clkbuf_2
X_07397_ _10103_/Q VGND VGND VPWR VPWR _07397_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06348_ _09935_/Q _06341_/A _09660_/A1 _06342_/A VGND VGND VPWR VPWR _09935_/D sky130_fd_sc_hd__a22o_1
X_09136_ _09399_/B _09136_/B VGND VGND VPWR VPWR _09138_/A sky130_fd_sc_hd__or2_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06279_ _06279_/A VGND VGND VPWR VPWR _06280_/B sky130_fd_sc_hd__clkbuf_4
X_09067_ _09067_/A _09067_/B VGND VGND VPWR VPWR _09442_/C sky130_fd_sc_hd__or2_1
XFILLER_190_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08018_ _08026_/A _10002_/Q _08032_/B _10006_/Q VGND VGND VPWR VPWR _08186_/A sky130_fd_sc_hd__or4_4
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09969_ _10283_/CLK _09969_/D repeater406/X VGND VGND VPWR VPWR _09969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10109_ _10482_/CLK _10109_/D _07492_/B VGND VGND VPWR VPWR _10109_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05650_ _10308_/Q _05641_/A _09659_/A1 _05642_/A VGND VGND VPWR VPWR _10308_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05581_ _10349_/Q _05577_/X _09580_/X _05579_/X VGND VGND VPWR VPWR _10349_/D sky130_fd_sc_hd__a22o_1
X_07320_ _10150_/Q VGND VGND VPWR VPWR _07320_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07251_ _10117_/Q VGND VGND VPWR VPWR _07251_/Y sky130_fd_sc_hd__inv_2
X_07182_ _10409_/Q VGND VGND VPWR VPWR _07182_/Y sky130_fd_sc_hd__clkinv_4
X_06202_ _06147_/X _06193_/Y _06200_/Y _10003_/Q _06203_/A VGND VGND VPWR VPWR _10003_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06133_ _09778_/Q VGND VGND VPWR VPWR _06133_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06064_ _10064_/Q _06056_/A _09661_/A1 _06057_/A VGND VGND VPWR VPWR _10064_/D sky130_fd_sc_hd__a22o_1
X_05015_ _10438_/Q _05008_/X _06684_/B1 _05010_/X VGND VGND VPWR VPWR _10438_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09823_ _10405_/CLK _09823_/D repeater410/X VGND VGND VPWR VPWR _09823_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09754_ _09781_/CLK _09754_/D VGND VGND VPWR VPWR _09754_/Q sky130_fd_sc_hd__dfxtp_1
X_06966_ _06961_/Y _04885_/A _06962_/Y _05927_/A _06965_/X VGND VGND VPWR VPWR _06985_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09685_ _08360_/X input176/X _09698_/S VGND VGND VPWR VPWR _09685_/X sky130_fd_sc_hd__mux2_1
X_05917_ _10154_/Q _05911_/X _09574_/X _05912_/Y VGND VGND VPWR VPWR _10154_/D sky130_fd_sc_hd__a22o_1
X_06897_ _10242_/Q VGND VGND VPWR VPWR _06897_/Y sky130_fd_sc_hd__inv_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08705_ _09109_/A _08650_/A _08684_/A _09109_/A _08704_/X VGND VGND VPWR VPWR _08705_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08636_ _08634_/A _08890_/B _08635_/Y VGND VGND VPWR VPWR _08656_/A sky130_fd_sc_hd__a21oi_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ _10195_/Q _05841_/A _09660_/A1 _05842_/A VGND VGND VPWR VPWR _10195_/D sky130_fd_sc_hd__a22o_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08567_ _08567_/A _09233_/C VGND VGND VPWR VPWR _09180_/A sky130_fd_sc_hd__or2_2
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05779_ _10235_/Q _05776_/X _09577_/X _05777_/Y VGND VGND VPWR VPWR _10235_/D sky130_fd_sc_hd__a22o_1
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ _08552_/A VGND VGND VPWR VPWR _08585_/A sky130_fd_sc_hd__buf_2
X_07518_ _07769_/A VGND VGND VPWR VPWR _07519_/A sky130_fd_sc_hd__buf_2
XFILLER_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07449_ _05367_/X _07440_/A _09742_/Q _07441_/A VGND VGND VPWR VPWR _09742_/D sky130_fd_sc_hd__o22a_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10460_ _10486_/CLK _10460_/D _05034_/A VGND VGND VPWR VPWR _10460_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_108_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09119_ _09446_/B _09286_/A VGND VGND VPWR VPWR _09119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10391_ _04811_/A1 _10391_/D _05471_/X VGND VGND VPWR VPWR _10391_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _04807_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_186_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06820_ _06815_/Y _04886_/B _06816_/Y _06154_/B _06819_/X VGND VGND VPWR VPWR _06833_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06751_ _10148_/Q VGND VGND VPWR VPWR _06751_/Y sky130_fd_sc_hd__clkinv_2
X_09470_ _09470_/A VGND VGND VPWR VPWR _09470_/X sky130_fd_sc_hd__clkbuf_1
X_06682_ _09769_/Q _06681_/A _09658_/A1 _06681_/Y VGND VGND VPWR VPWR _09769_/D sky130_fd_sc_hd__a22o_1
X_05702_ _05702_/A VGND VGND VPWR VPWR _05702_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08421_ _08695_/A _08530_/D _08430_/B VGND VGND VPWR VPWR _08424_/B sky130_fd_sc_hd__or3_1
XFILLER_91_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05633_ _10320_/Q _05627_/X _09545_/A1 _05629_/X VGND VGND VPWR VPWR _10320_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05564_ _09787_/D _09783_/Q _09785_/Q _09784_/Q VGND VGND VPWR VPWR _05564_/X sky130_fd_sc_hd__or4_1
X_08352_ _08349_/Y _08348_/Y _09814_/Q _08351_/Y VGND VGND VPWR VPWR _08352_/Y sky130_fd_sc_hd__a31oi_1
X_05495_ _09691_/X _10385_/Q _05512_/S VGND VGND VPWR VPWR _05496_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08283_ _07277_/Y _08195_/X _07228_/Y _08196_/X VGND VGND VPWR VPWR _08283_/X sky130_fd_sc_hd__o22a_1
X_07303_ _07303_/A _07303_/B _07303_/C _07302_/X VGND VGND VPWR VPWR _07420_/A sky130_fd_sc_hd__or4b_1
XFILLER_177_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07234_ _09830_/Q VGND VGND VPWR VPWR _07234_/Y sky130_fd_sc_hd__inv_2
X_07165_ input111/X _05112_/X _10326_/Q _05156_/Y VGND VGND VPWR VPWR _07165_/X sky130_fd_sc_hd__a22o_1
X_07096_ _10214_/Q VGND VGND VPWR VPWR _09511_/A sky130_fd_sc_hd__inv_4
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06116_ _10032_/Q _06109_/X _09658_/A1 _06111_/X VGND VGND VPWR VPWR _10032_/D sky130_fd_sc_hd__a22o_1
XFILLER_182_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06047_ _06047_/A VGND VGND VPWR VPWR _06047_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09806_ net399_2/A _09806_/D _06600_/X VGND VGND VPWR VPWR _09806_/Q sky130_fd_sc_hd__dfrtp_1
X_07998_ _08046_/C VGND VGND VPWR VPWR _08044_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09737_ _09781_/CLK _09737_/D VGND VGND VPWR VPWR _09737_/Q sky130_fd_sc_hd__dfxtp_1
X_06949_ _09796_/Q VGND VGND VPWR VPWR _06949_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09668_ _09667_/X _10393_/Q _10299_/Q VGND VGND VPWR VPWR _09668_/X sky130_fd_sc_hd__mux2_4
X_08619_ _08771_/A _09084_/B VGND VGND VPWR VPWR _08879_/A sky130_fd_sc_hd__or2_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09598_/X _09911_/Q _09776_/Q VGND VGND VPWR VPWR _09599_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10512_ _10512_/CLK _10512_/D _07492_/B VGND VGND VPWR VPWR _10512_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10443_ _10487_/CLK _10443_/D _05034_/A VGND VGND VPWR VPWR _10443_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10374_ _10374_/CLK _10374_/D hold41/X VGND VGND VPWR VPWR _10374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _05406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 _07098_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 _07799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 _10406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05280_ _05271_/Y _05895_/A _05273_/Y _04885_/A _05279_/X VGND VGND VPWR VPWR _05281_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08970_ _08970_/A _08974_/B _09005_/A VGND VGND VPWR VPWR _09427_/B sky130_fd_sc_hd__nor3_2
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07921_ _07240_/Y _07512_/A _07269_/Y _07802_/X VGND VGND VPWR VPWR _07921_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_30_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10349_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07852_ _06754_/Y _07818_/X _07851_/Y _07819_/X VGND VGND VPWR VPWR _07852_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06803_ _10264_/Q VGND VGND VPWR VPWR _06803_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
X_07783_ _07783_/A VGND VGND VPWR VPWR _07783_/X sky130_fd_sc_hd__buf_2
X_09522_ _09522_/A VGND VGND VPWR VPWR _09522_/X sky130_fd_sc_hd__clkbuf_1
X_04995_ _04995_/A VGND VGND VPWR VPWR _04996_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_45_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10341_/CLK sky130_fd_sc_hd__clkbuf_16
X_06734_ _09827_/Q VGND VGND VPWR VPWR _06734_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09453_ _09444_/Y _09445_/Y _09447_/X _09452_/X VGND VGND VPWR VPWR _09453_/X sky130_fd_sc_hd__a31o_1
XFILLER_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08404_ _09233_/A VGND VGND VPWR VPWR _08417_/A sky130_fd_sc_hd__inv_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09384_ _09415_/B _09384_/B _09384_/C VGND VGND VPWR VPWR _09385_/C sky130_fd_sc_hd__or3_1
X_05616_ _05617_/A VGND VGND VPWR VPWR _05616_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08335_ _09801_/Q _08335_/B _09802_/Q VGND VGND VPWR VPWR _08338_/B sky130_fd_sc_hd__and3_1
X_06596_ _06614_/A VGND VGND VPWR VPWR _06597_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_177_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05547_ _10366_/Q _05542_/X _06684_/B1 _05543_/Y VGND VGND VPWR VPWR _10366_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08266_ _07390_/Y _08193_/X _07371_/Y _08194_/X _08265_/X VGND VGND VPWR VPWR _08273_/A
+ sky130_fd_sc_hd__o221a_1
X_05478_ _10389_/Q _05475_/X _09658_/A1 _05476_/Y VGND VGND VPWR VPWR _10389_/D sky130_fd_sc_hd__a22o_1
X_08197_ _06817_/Y _08195_/X _06822_/Y _08196_/X VGND VGND VPWR VPWR _08197_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07217_ _07212_/Y _05865_/B _07213_/Y _05821_/B _07216_/X VGND VGND VPWR VPWR _07218_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07148_ _07146_/Y _06167_/B _09501_/A _05793_/A VGND VGND VPWR VPWR _07148_/X sky130_fd_sc_hd__o22a_1
X_07079_ _10170_/Q VGND VGND VPWR VPWR _09497_/A sky130_fd_sc_hd__inv_6
Xoutput371 _09759_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput360 _09758_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10090_ _10119_/CLK _10090_/D repeater403/X VGND VGND VPWR VPWR _10090_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_160_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput382 _09760_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10426_ net399_2/A _10426_/D _05051_/X VGND VGND VPWR VPWR _10426_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10357_ _10364_/CLK _10357_/D repeater410/X VGND VGND VPWR VPWR _10357_/Q sky130_fd_sc_hd__dfstp_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/CLK _10288_/D repeater406/X VGND VGND VPWR VPWR _10288_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06450_ _09868_/Q _06441_/A _09659_/A1 _06442_/A VGND VGND VPWR VPWR _09868_/D sky130_fd_sc_hd__a22o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05401_ _05401_/A VGND VGND VPWR VPWR _05401_/X sky130_fd_sc_hd__clkbuf_1
X_06381_ _06380_/X _09603_/X _09650_/X _09914_/Q VGND VGND VPWR VPWR _09914_/D sky130_fd_sc_hd__o22a_1
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05332_ _10351_/Q VGND VGND VPWR VPWR _05332_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08120_ _09457_/A _08060_/X _09501_/A _08061_/X VGND VGND VPWR VPWR _08120_/X sky130_fd_sc_hd__o22a_1
X_05263_ _10258_/Q VGND VGND VPWR VPWR _05263_/Y sky130_fd_sc_hd__inv_4
X_08051_ _08051_/A VGND VGND VPWR VPWR _08051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07002_ _06986_/Y _06079_/B _06989_/X _06995_/X _07001_/X VGND VGND VPWR VPWR _07028_/C
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_opt_5_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_5_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05194_ _05340_/A _05316_/B VGND VGND VPWR VPWR _06036_/A sky130_fd_sc_hd__or2_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08953_ _08957_/A _08961_/B VGND VGND VPWR VPWR _09386_/B sky130_fd_sc_hd__nor2_1
X_07904_ _10124_/Q VGND VGND VPWR VPWR _07904_/Y sky130_fd_sc_hd__clkinv_2
X_08884_ _08884_/A _08908_/A VGND VGND VPWR VPWR _08884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07835_ _06718_/Y _07782_/X _06731_/Y _07783_/X VGND VGND VPWR VPWR _07835_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04978_ _04992_/A _05148_/A VGND VGND VPWR VPWR _05088_/A sky130_fd_sc_hd__or2_1
XFILLER_44_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07766_ _06898_/Y _07658_/X _07765_/Y _07659_/X VGND VGND VPWR VPWR _07766_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09505_ _09505_/A VGND VGND VPWR VPWR _09506_/A sky130_fd_sc_hd__clkbuf_1
X_06717_ _10044_/Q VGND VGND VPWR VPWR _06717_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09436_ _09441_/A _09443_/C _09435_/Y VGND VGND VPWR VPWR _09436_/Y sky130_fd_sc_hd__o21ai_1
X_07697_ _09477_/A _07620_/X _07050_/Y _07621_/X _07696_/X VGND VGND VPWR VPWR _07697_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06648_ _06648_/A VGND VGND VPWR VPWR _06648_/X sky130_fd_sc_hd__clkbuf_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A VGND VGND VPWR VPWR _09367_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06579_ _09808_/Q _06579_/B _09809_/Q _06579_/D VGND VGND VPWR VPWR _06580_/A sky130_fd_sc_hd__or4_1
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09298_ _09298_/A _09358_/B _09390_/B _09433_/B VGND VGND VPWR VPWR _09300_/B sky130_fd_sc_hd__or4_1
XANTENNA_50 _04807_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08318_ _06951_/Y _08183_/A _08315_/X _08317_/X VGND VGND VPWR VPWR _08328_/C sky130_fd_sc_hd__o211a_1
XANTENNA_83 _07502_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08249_ _05337_/Y _08201_/X _07872_/Y _08202_/X VGND VGND VPWR VPWR _08249_/X sky130_fd_sc_hd__o22a_1
XANTENNA_61 _10482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10211_ _10491_/CLK _10211_/D repeater402/X VGND VGND VPWR VPWR _10211_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10142_ _10238_/CLK _10142_/D repeater403/X VGND VGND VPWR VPWR _10142_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10073_ _10512_/CLK _10073_/D _07492_/B VGND VGND VPWR VPWR _10073_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10409_ _10409_/CLK _10409_/D repeater406/X VGND VGND VPWR VPWR _10409_/Q sky130_fd_sc_hd__dfstp_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _09752_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05950_ _10134_/Q _05942_/A _06684_/B1 _05943_/A VGND VGND VPWR VPWR _10134_/D sky130_fd_sc_hd__a22o_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05881_ _10175_/Q _05875_/X _09574_/X _05876_/Y VGND VGND VPWR VPWR _10175_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04901_ _06538_/A _05124_/A VGND VGND VPWR VPWR _04903_/A sky130_fd_sc_hd__or2_1
X_07620_ _07779_/A VGND VGND VPWR VPWR _07620_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04832_ _04991_/B VGND VGND VPWR VPWR _05109_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_07551_ _09991_/Q _07551_/B _09989_/Q _09988_/Q VGND VGND VPWR VPWR _07575_/B sky130_fd_sc_hd__or4_1
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06502_ _06502_/A VGND VGND VPWR VPWR _06503_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07482_ _07482_/A VGND VGND VPWR VPWR _09781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09221_ _09221_/A VGND VGND VPWR VPWR _09221_/X sky130_fd_sc_hd__clkbuf_1
X_06433_ _09880_/Q _06431_/X _09578_/X _06432_/Y VGND VGND VPWR VPWR _09880_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09152_ _09152_/A _09152_/B VGND VGND VPWR VPWR _09156_/B sky130_fd_sc_hd__or2_1
X_06364_ _09927_/Q _06361_/X _09581_/X _06363_/X VGND VGND VPWR VPWR _09927_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05315_ _10180_/Q VGND VGND VPWR VPWR _05315_/Y sky130_fd_sc_hd__inv_2
X_08103_ _07207_/Y _08058_/X _07259_/Y _08059_/X _08102_/X VGND VGND VPWR VPWR _08117_/B
+ sky130_fd_sc_hd__o221a_1
X_09083_ _09295_/C _09083_/B _09083_/C VGND VGND VPWR VPWR _09276_/A sky130_fd_sc_hd__or3_1
X_06295_ _09967_/Q _06292_/X _09581_/X _06294_/X VGND VGND VPWR VPWR _09967_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_4
X_05246_ _05241_/Y _06153_/A _05244_/Y _05540_/A VGND VGND VPWR VPWR _05246_/X sky130_fd_sc_hd__o22a_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__buf_4
X_08034_ _08034_/A _08040_/A _10006_/Q VGND VGND VPWR VPWR _08202_/A sky130_fd_sc_hd__or3_4
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__buf_2
X_05177_ _05177_/A VGND VGND VPWR VPWR _06045_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09985_ _10283_/CLK _09985_/D repeater406/X VGND VGND VPWR VPWR _09985_/Q sky130_fd_sc_hd__dfstp_1
X_08936_ _08936_/A _08943_/A VGND VGND VPWR VPWR _09442_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08867_ _09400_/A _08867_/B VGND VGND VPWR VPWR _08868_/B sky130_fd_sc_hd__or2_1
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07818_ _07818_/A VGND VGND VPWR VPWR _07818_/X sky130_fd_sc_hd__clkbuf_2
X_08798_ _08895_/C VGND VGND VPWR VPWR _08913_/C sky130_fd_sc_hd__inv_2
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07749_ _07749_/A VGND VGND VPWR VPWR _07749_/X sky130_fd_sc_hd__buf_4
X_09419_ _09419_/A _09419_/B _09419_/C VGND VGND VPWR VPWR _09445_/A sky130_fd_sc_hd__or3_2
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10125_ _10127_/CLK _10125_/D _07492_/B VGND VGND VPWR VPWR _10125_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10056_ _10482_/CLK _10056_/D repeater405/X VGND VGND VPWR VPWR _10056_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05100_ _05157_/A _05100_/B VGND VGND VPWR VPWR _05101_/A sky130_fd_sc_hd__nor2_2
X_06080_ _06081_/A VGND VGND VPWR VPWR _06080_/X sky130_fd_sc_hd__clkbuf_2
X_05031_ _05031_/A _05031_/B VGND VGND VPWR VPWR _05031_/X sky130_fd_sc_hd__or2_1
XFILLER_112_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _10411_/Q VGND VGND VPWR VPWR _06982_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09770_ _10406_/CLK _09770_/D _06678_/X VGND VGND VPWR VPWR _09770_/Q sky130_fd_sc_hd__dfstp_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05933_ _10147_/Q _05929_/X _09580_/X _05931_/X VGND VGND VPWR VPWR _10147_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08721_ _08721_/A _09168_/A VGND VGND VPWR VPWR _08721_/X sky130_fd_sc_hd__and2_1
XFILLER_66_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _08640_/A _08641_/B _08890_/B VGND VGND VPWR VPWR _08667_/A sky130_fd_sc_hd__a21bo_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05864_ _05864_/A VGND VGND VPWR VPWR _05865_/B sky130_fd_sc_hd__buf_2
X_07603_ _10107_/Q VGND VGND VPWR VPWR _07603_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05795_ _05796_/A VGND VGND VPWR VPWR _05795_/X sky130_fd_sc_hd__clkbuf_2
X_08583_ _08583_/A _08951_/B VGND VGND VPWR VPWR _09309_/A sky130_fd_sc_hd__nor2_1
X_04815_ _09676_/X VGND VGND VPWR VPWR _04963_/B sky130_fd_sc_hd__inv_2
XFILLER_179_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07534_ _07534_/A _07549_/B VGND VGND VPWR VPWR _07606_/B sky130_fd_sc_hd__or2_1
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07465_ _09532_/A _09531_/A _07438_/B VGND VGND VPWR VPWR _09788_/D sky130_fd_sc_hd__o21ai_1
XFILLER_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09204_ _09204_/A _09204_/B VGND VGND VPWR VPWR _09407_/C sky130_fd_sc_hd__nor2_1
X_06416_ _06386_/X _09633_/X _09650_/X _09891_/Q VGND VGND VPWR VPWR _09891_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07396_ _10238_/Q VGND VGND VPWR VPWR _07396_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06347_ _09936_/Q _06340_/X _09550_/A0 _06342_/X VGND VGND VPWR VPWR _09936_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09135_ _09135_/A _09313_/D VGND VGND VPWR VPWR _09136_/B sky130_fd_sc_hd__or2_1
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09066_ _09066_/A _09285_/C _09354_/C _09286_/C VGND VGND VPWR VPWR _09070_/A sky130_fd_sc_hd__or4_2
X_06278_ _09974_/Q _06269_/A _09659_/A1 _06270_/A VGND VGND VPWR VPWR _09974_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05229_ _05229_/A VGND VGND VPWR VPWR _06351_/B sky130_fd_sc_hd__clkbuf_2
X_08017_ _05189_/Y _08184_/A _05221_/Y _08158_/A VGND VGND VPWR VPWR _08017_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09968_ _10023_/CLK _09968_/D _05034_/A VGND VGND VPWR VPWR _09968_/Q sky130_fd_sc_hd__dfrtp_1
X_08919_ _09307_/C _08919_/B _08919_/C _08918_/X VGND VGND VPWR VPWR _08922_/B sky130_fd_sc_hd__or4b_2
X_09899_ _10268_/CLK _09899_/D repeater404/X VGND VGND VPWR VPWR _09899_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10108_ _10482_/CLK _10108_/D repeater405/X VGND VGND VPWR VPWR _10108_/Q sky130_fd_sc_hd__dfstp_1
X_10039_ _10404_/CLK _10039_/D repeater410/X VGND VGND VPWR VPWR _10039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05580_ _10350_/Q _05577_/X _09581_/X _05579_/X VGND VGND VPWR VPWR _10350_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07250_ _09971_/Q VGND VGND VPWR VPWR _07932_/A sky130_fd_sc_hd__inv_4
XFILLER_176_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07181_ _07181_/A _07181_/B _07181_/C _07180_/X VGND VGND VPWR VPWR _07193_/B sky130_fd_sc_hd__or4b_2
X_06201_ _09775_/Q _09777_/Q VGND VGND VPWR VPWR _06203_/A sky130_fd_sc_hd__or2_4
X_06132_ _09776_/Q VGND VGND VPWR VPWR _07477_/A sky130_fd_sc_hd__clkinv_2
XFILLER_144_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06063_ _10065_/Q _06056_/A _09660_/A1 _06057_/A VGND VGND VPWR VPWR _10065_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05014_ _10439_/Q _05008_/X _06683_/B1 _05010_/X VGND VGND VPWR VPWR _10439_/D sky130_fd_sc_hd__a22o_1
X_09822_ _10364_/CLK _09822_/D repeater410/X VGND VGND VPWR VPWR _09822_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09753_ _09781_/CLK _09753_/D VGND VGND VPWR VPWR _09753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06965_ _06963_/Y _06053_/A _06964_/Y _05775_/B VGND VGND VPWR VPWR _06965_/X sky130_fd_sc_hd__o22a_1
X_08704_ _09324_/A _08700_/X _08704_/C _09149_/B VGND VGND VPWR VPWR _08704_/X sky130_fd_sc_hd__and4bb_1
XFILLER_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09684_ _08358_/X input165/X _09698_/S VGND VGND VPWR VPWR _09684_/X sky130_fd_sc_hd__mux2_1
X_05916_ _10155_/Q _05911_/X hold46/X _05912_/Y VGND VGND VPWR VPWR _10155_/D sky130_fd_sc_hd__a22o_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06896_ _06894_/Y _05883_/B _06895_/Y _06154_/B VGND VGND VPWR VPWR _06896_/X sky130_fd_sc_hd__o22a_1
X_08635_ _08888_/B VGND VGND VPWR VPWR _08635_/Y sky130_fd_sc_hd__clkinvlp_2
X_05847_ _10196_/Q _05840_/X _09550_/A0 _05842_/X VGND VGND VPWR VPWR _10196_/D sky130_fd_sc_hd__a22o_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08566_ _08695_/C VGND VGND VPWR VPWR _09233_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05778_ _10236_/Q _05776_/X _09578_/X _05777_/Y VGND VGND VPWR VPWR _10236_/D sky130_fd_sc_hd__a22o_1
X_07517_ _07564_/C _07608_/B VGND VGND VPWR VPWR _07769_/A sky130_fd_sc_hd__or2_1
XFILLER_167_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08497_ _09085_/D _09102_/B _09102_/C _08624_/A VGND VGND VPWR VPWR _08552_/A sky130_fd_sc_hd__or4_4
X_07448_ _07421_/X _07440_/A _09743_/Q _07441_/A VGND VGND VPWR VPWR _09743_/D sky130_fd_sc_hd__o22a_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ _07377_/Y _05851_/A _07378_/Y _05910_/B VGND VGND VPWR VPWR _07379_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09118_ _09118_/A VGND VGND VPWR VPWR _09446_/B sky130_fd_sc_hd__inv_2
XFILLER_135_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10390_ _10500_/CLK _10390_/D repeater407/X VGND VGND VPWR VPWR _10390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09049_ _08553_/B _08686_/Y _08801_/C VGND VGND VPWR VPWR _09049_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06750_ _06745_/Y _05808_/B _06746_/Y _06893_/B _06749_/X VGND VGND VPWR VPWR _06750_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06681_ _06681_/A VGND VGND VPWR VPWR _06681_/Y sky130_fd_sc_hd__inv_2
X_05701_ _05701_/A VGND VGND VPWR VPWR _05701_/X sky130_fd_sc_hd__clkbuf_2
X_08420_ _08556_/B VGND VGND VPWR VPWR _08530_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_05632_ _10321_/Q _05627_/X _09579_/X _05629_/X VGND VGND VPWR VPWR _10321_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05563_ _05563_/A VGND VGND VPWR VPWR _05563_/X sky130_fd_sc_hd__clkbuf_1
X_08351_ _08349_/Y _08348_/Y _09814_/Q VGND VGND VPWR VPWR _08351_/Y sky130_fd_sc_hd__a21oi_1
X_05494_ _05525_/S VGND VGND VPWR VPWR _05512_/S sky130_fd_sc_hd__clkbuf_2
X_08282_ _07196_/Y _08183_/X _08279_/X _08281_/X VGND VGND VPWR VPWR _08292_/C sky130_fd_sc_hd__o211a_1
X_07302_ _07298_/Y _05980_/B _07299_/Y _06066_/B _07301_/X VGND VGND VPWR VPWR _07302_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07233_ _09996_/Q VGND VGND VPWR VPWR _07233_/Y sky130_fd_sc_hd__clkinv_4
X_07164_ input115/X _06696_/X _10339_/Q _05126_/Y _07163_/X VGND VGND VPWR VPWR _07167_/B
+ sky130_fd_sc_hd__a221o_1
X_07095_ _09491_/A _06010_/A _09505_/A _04885_/A _07094_/X VGND VGND VPWR VPWR _07114_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06115_ _10033_/Q _06109_/X _09545_/A1 _06111_/X VGND VGND VPWR VPWR _10033_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06046_ _06047_/A VGND VGND VPWR VPWR _06046_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09805_ net399_2/A _09805_/D _06609_/X VGND VGND VPWR VPWR _09805_/Q sky130_fd_sc_hd__dfrtp_2
X_07997_ _08006_/A _08000_/B VGND VGND VPWR VPWR _08046_/C sky130_fd_sc_hd__or2_1
XFILLER_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06948_ _10262_/Q VGND VGND VPWR VPWR _06948_/Y sky130_fd_sc_hd__inv_2
X_09736_ _09781_/CLK _09736_/D VGND VGND VPWR VPWR _09736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09667_ _09801_/Q _09800_/Q _09773_/Q VGND VGND VPWR VPWR _09667_/X sky130_fd_sc_hd__mux2_1
X_08618_ _09057_/B VGND VGND VPWR VPWR _09084_/B sky130_fd_sc_hd__buf_4
X_06879_ _06874_/Y _05576_/B _06875_/Y _05550_/B _06878_/X VGND VGND VPWR VPWR _06880_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _08172_/Y _10334_/Q _09700_/S VGND VGND VPWR VPWR _09598_/X sky130_fd_sc_hd__mux2_1
X_08549_ _08687_/A _08697_/A VGND VGND VPWR VPWR _08813_/A sky130_fd_sc_hd__or2_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10511_ _10512_/CLK _10511_/D _07492_/B VGND VGND VPWR VPWR _10511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10442_ _10487_/CLK _10442_/D repeater409/X VGND VGND VPWR VPWR _10442_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10373_ _10374_/CLK _10373_/D hold41/X VGND VGND VPWR VPWR _10373_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _05406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _07440_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _09521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_195 _09487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07920_ _07206_/Y _07792_/X _07258_/Y _07793_/X _07919_/X VGND VGND VPWR VPWR _07926_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07851_ _10114_/Q VGND VGND VPWR VPWR _07851_/Y sky130_fd_sc_hd__clkinv_2
X_06802_ _09966_/Q VGND VGND VPWR VPWR _06802_/Y sky130_fd_sc_hd__clkinv_2
X_07782_ _07782_/A VGND VGND VPWR VPWR _07782_/X sky130_fd_sc_hd__buf_2
XFILLER_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_2
X_06733_ _06728_/Y _04886_/B _06729_/Y _05749_/B _06732_/X VGND VGND VPWR VPWR _06740_/C
+ sky130_fd_sc_hd__o221a_1
X_09521_ input68/X _09521_/B VGND VGND VPWR VPWR _09522_/A sky130_fd_sc_hd__and2_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_2_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
X_04994_ _04995_/A VGND VGND VPWR VPWR _04994_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06664_ _06664_/A VGND VGND VPWR VPWR _06664_/X sky130_fd_sc_hd__clkbuf_1
X_09452_ _09424_/B _09449_/Y _09401_/A _09450_/Y _09451_/Y VGND VGND VPWR VPWR _09452_/X
+ sky130_fd_sc_hd__o311a_1
X_08403_ _08571_/C VGND VGND VPWR VPWR _08634_/A sky130_fd_sc_hd__inv_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09383_ _09447_/D _09411_/D _09383_/C _09415_/A VGND VGND VPWR VPWR _09383_/Y sky130_fd_sc_hd__nor4_1
X_05615_ _05775_/A _05615_/B VGND VGND VPWR VPWR _05617_/A sky130_fd_sc_hd__or2_1
X_06595_ _06668_/A VGND VGND VPWR VPWR _06614_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05546_ _10367_/Q _05542_/X _06683_/B1 _05543_/Y VGND VGND VPWR VPWR _10367_/D sky130_fd_sc_hd__a22o_1
X_08334_ _09801_/Q _08335_/B _09801_/Q _08335_/B VGND VGND VPWR VPWR _08334_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08265_ _07340_/Y _08195_/X _07383_/Y _08196_/X VGND VGND VPWR VPWR _08265_/X sky130_fd_sc_hd__o22a_1
X_05477_ _10390_/Q _05475_/X _09545_/A1 _05476_/Y VGND VGND VPWR VPWR _10390_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07216_ _07214_/Y _05993_/B _07215_/Y _05262_/A VGND VGND VPWR VPWR _07216_/X sky130_fd_sc_hd__o22a_1
X_08196_ _08196_/A VGND VGND VPWR VPWR _08196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07147_ _10222_/Q VGND VGND VPWR VPWR _09501_/A sky130_fd_sc_hd__inv_6
XFILLER_105_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07078_ _09936_/Q VGND VGND VPWR VPWR _09475_/A sky130_fd_sc_hd__clkinv_4
XFILLER_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput361 _09744_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput350 _10473_/Q VGND VGND VPWR VPWR sram_ro_addr[1] sky130_fd_sc_hd__buf_2
Xoutput383 _09740_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput372 _09754_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_2
X_06029_ _10087_/Q _06025_/X _09580_/X _06027_/X VGND VGND VPWR VPWR _10087_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09719_ _10505_/Q _09491_/A VGND VGND VPWR VPWR _09719_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10425_ net399_2/A _10425_/D _05054_/X VGND VGND VPWR VPWR _10425_/Q sky130_fd_sc_hd__dfrtn_1
X_10356_ _10382_/CLK _10356_/D _05563_/X VGND VGND VPWR VPWR _10356_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10288_/CLK _10287_/D repeater406/X VGND VGND VPWR VPWR _10287_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05400_ _05406_/A VGND VGND VPWR VPWR _05401_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06380_ _06417_/A VGND VGND VPWR VPWR _06380_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05331_ _05322_/Y _06359_/A _05324_/Y _05433_/A _05330_/X VGND VGND VPWR VPWR _05364_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_186_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05262_ _05262_/A VGND VGND VPWR VPWR _06635_/B sky130_fd_sc_hd__clkbuf_2
X_08050_ _08050_/A _08050_/B _08050_/C _08050_/D VGND VGND VPWR VPWR _08051_/A sky130_fd_sc_hd__and4_1
XFILLER_162_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07001_ _06996_/Y _05993_/B _06997_/Y _06708_/B _07000_/X VGND VGND VPWR VPWR _07001_/X
+ sky130_fd_sc_hd__o221a_1
X_05193_ _05299_/B VGND VGND VPWR VPWR _05316_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08952_ _08952_/A _09201_/B VGND VGND VPWR VPWR _08954_/A sky130_fd_sc_hd__or2_1
X_08883_ _08883_/A _08883_/B VGND VGND VPWR VPWR _09318_/B sky130_fd_sc_hd__nor2_2
X_07903_ _07352_/Y _07762_/X _07318_/Y _07811_/X _07902_/X VGND VGND VPWR VPWR _07911_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07834_ _10088_/Q VGND VGND VPWR VPWR _07834_/Y sky130_fd_sc_hd__inv_2
X_07765_ _10112_/Q VGND VGND VPWR VPWR _07765_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04977_ _05027_/A _04991_/B _09674_/X _05109_/B VGND VGND VPWR VPWR _05148_/A sky130_fd_sc_hd__or4_1
X_09504_ _09504_/A VGND VGND VPWR VPWR _09504_/X sky130_fd_sc_hd__clkbuf_1
X_07696_ _09493_/A _07622_/X _09491_/A _07623_/X VGND VGND VPWR VPWR _07696_/X sky130_fd_sc_hd__o22a_1
X_06716_ _10019_/Q VGND VGND VPWR VPWR _06716_/Y sky130_fd_sc_hd__clkinv_2
X_06647_ _06655_/A VGND VGND VPWR VPWR _06648_/A sky130_fd_sc_hd__clkbuf_1
X_09435_ _09435_/A _09435_/B _09435_/C VGND VGND VPWR VPWR _09435_/Y sky130_fd_sc_hd__nor3_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _09417_/A _09419_/B _09332_/Y _09349_/X _09365_/X VGND VGND VPWR VPWR _09367_/A
+ sky130_fd_sc_hd__o311a_1
X_06578_ _06578_/A VGND VGND VPWR VPWR _06578_/X sky130_fd_sc_hd__clkbuf_1
X_09297_ _09297_/A _09297_/B VGND VGND VPWR VPWR _09433_/B sky130_fd_sc_hd__or2_1
XFILLER_138_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08317_ _06999_/Y _08186_/A _06957_/Y _08187_/A _08316_/X VGND VGND VPWR VPWR _08317_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_40 _07650_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05529_ _05530_/A VGND VGND VPWR VPWR _05529_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08248_ _05227_/Y _08193_/X _05186_/Y _08194_/X _08247_/X VGND VGND VPWR VPWR _08255_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA_51 _10342_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _09867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 input22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_95 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _10409_/CLK _10210_/D repeater406/X VGND VGND VPWR VPWR _10210_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08179_ _08179_/A VGND VGND VPWR VPWR _08179_/X sky130_fd_sc_hd__buf_2
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ _10238_/CLK _10141_/D repeater403/X VGND VGND VPWR VPWR _10141_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ _10512_/CLK _10072_/D _07492_/B VGND VGND VPWR VPWR _10072_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10513_/CLK sky130_fd_sc_hd__clkbuf_16
X_10408_ _10409_/CLK _10408_/D repeater406/X VGND VGND VPWR VPWR _10408_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10341_/CLK _10339_/D repeater409/X VGND VGND VPWR VPWR _10339_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04900_ _05157_/A _05327_/A VGND VGND VPWR VPWR _05124_/A sky130_fd_sc_hd__or2_2
X_05880_ _10176_/Q _05875_/X _09661_/A1 _05876_/Y VGND VGND VPWR VPWR _10176_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04831_ _09668_/X VGND VGND VPWR VPWR _04991_/B sky130_fd_sc_hd__inv_2
X_07550_ _07789_/A VGND VGND VPWR VPWR _07629_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06501_ _09849_/Q _06495_/X _09574_/X _06496_/Y VGND VGND VPWR VPWR _09849_/D sky130_fd_sc_hd__a22o_1
X_07481_ _09787_/Q _07481_/B VGND VGND VPWR VPWR _07482_/A sky130_fd_sc_hd__or2_1
X_09220_ _09315_/A _09220_/B _09315_/C _09220_/D VGND VGND VPWR VPWR _09221_/A sky130_fd_sc_hd__or4_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06432_ _06432_/A VGND VGND VPWR VPWR _06432_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09151_ _08570_/B _08710_/A _08563_/X VGND VGND VPWR VPWR _09152_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06363_ _06363_/A VGND VGND VPWR VPWR _06363_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09082_ _09082_/A _09248_/A VGND VGND VPWR VPWR _09086_/B sky130_fd_sc_hd__or2_1
X_05314_ _05314_/A VGND VGND VPWR VPWR _05740_/B sky130_fd_sc_hd__clkbuf_4
X_08102_ _07195_/Y _08060_/X _07183_/Y _08061_/X VGND VGND VPWR VPWR _08102_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06294_ _06294_/A VGND VGND VPWR VPWR _06294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08033_ _08034_/A _08040_/A _08045_/D VGND VGND VPWR VPWR _08201_/A sky130_fd_sc_hd__or3_4
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_6
XFILLER_162_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_2
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_4
X_05245_ _05245_/A _05277_/A VGND VGND VPWR VPWR _05540_/A sky130_fd_sc_hd__or2_2
Xinput93 sram_ro_data[0] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_2
X_05176_ _06630_/A _05261_/B VGND VGND VPWR VPWR _05177_/A sky130_fd_sc_hd__or2_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09984_ _10355_/CLK _09984_/D repeater406/X VGND VGND VPWR VPWR _09984_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08935_ _08951_/A _08935_/B VGND VGND VPWR VPWR _09067_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08866_ _08866_/A _09079_/A _08865_/X VGND VGND VPWR VPWR _08867_/B sky130_fd_sc_hd__or3b_1
XFILLER_111_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08797_ _08379_/B _08795_/Y _08492_/B _08795_/A VGND VGND VPWR VPWR _08895_/C sky130_fd_sc_hd__o22a_1
XFILLER_123_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07817_ _07817_/A VGND VGND VPWR VPWR _07817_/X sky130_fd_sc_hd__clkbuf_2
X_07748_ _06897_/Y _07618_/X _06863_/Y _07619_/X _07747_/X VGND VGND VPWR VPWR _07776_/A
+ sky130_fd_sc_hd__o221a_1
X_07679_ _07227_/Y _07632_/X _07257_/Y _07633_/X _07678_/X VGND VGND VPWR VPWR _07684_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09418_ _09418_/A _09418_/B _09418_/C _09418_/D VGND VGND VPWR VPWR _09419_/C sky130_fd_sc_hd__or4_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09349_ _09333_/Y _09345_/Y _09347_/Y _09426_/C VGND VGND VPWR VPWR _09349_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10124_ _10127_/CLK _10124_/D _07492_/B VGND VGND VPWR VPWR _10124_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10055_ _10110_/CLK _10055_/D repeater405/X VGND VGND VPWR VPWR _10055_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05030_ _05031_/B VGND VGND VPWR VPWR _05030_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _10249_/Q VGND VGND VPWR VPWR _06981_/Y sky130_fd_sc_hd__inv_4
XFILLER_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05932_ _10148_/Q _05929_/X _09581_/X _05931_/X VGND VGND VPWR VPWR _10148_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08720_ _08732_/A _08841_/B VGND VGND VPWR VPWR _09168_/A sky130_fd_sc_hd__or2_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _09095_/A VGND VGND VPWR VPWR _08743_/A sky130_fd_sc_hd__buf_2
X_05863_ _10185_/Q _05854_/A _09659_/A1 _05855_/A VGND VGND VPWR VPWR _10185_/D sky130_fd_sc_hd__a22o_1
X_07602_ _09989_/Q _09988_/Q _07602_/C _07602_/D VGND VGND VPWR VPWR _07818_/A sky130_fd_sc_hd__or4_4
X_04814_ _09674_/X VGND VGND VPWR VPWR _05005_/C sky130_fd_sc_hd__inv_2
X_08582_ _08582_/A _08582_/B VGND VGND VPWR VPWR _08951_/B sky130_fd_sc_hd__or2_1
X_05794_ _05794_/A _05794_/B VGND VGND VPWR VPWR _05796_/A sky130_fd_sc_hd__or2_2
XFILLER_81_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07533_ _07533_/A _07533_/B _07533_/C _07533_/D VGND VGND VPWR VPWR _07568_/C sky130_fd_sc_hd__and4_1
X_07464_ _09533_/A _09531_/A _06469_/X VGND VGND VPWR VPWR _09786_/D sky130_fd_sc_hd__o21ai_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09203_ _08461_/X _09206_/A _08483_/D _08552_/X VGND VGND VPWR VPWR _09204_/B sky130_fd_sc_hd__o22a_1
X_06415_ _06386_/X _09635_/X _09650_/X _09892_/Q VGND VGND VPWR VPWR _09892_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07395_ _10212_/Q VGND VGND VPWR VPWR _07395_/Y sky130_fd_sc_hd__inv_2
X_09134_ _09184_/A _09248_/A VGND VGND VPWR VPWR _09313_/D sky130_fd_sc_hd__or2_2
X_06346_ _09937_/Q _06340_/X _09547_/A1 _06342_/X VGND VGND VPWR VPWR _09937_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09065_ _09065_/A _09065_/B VGND VGND VPWR VPWR _09286_/C sky130_fd_sc_hd__or2_1
X_06277_ _09975_/Q _06269_/A _09661_/A1 _06270_/A VGND VGND VPWR VPWR _09975_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05228_ _05261_/B _05275_/B VGND VGND VPWR VPWR _05229_/A sky130_fd_sc_hd__or2_1
X_08016_ _08016_/A VGND VGND VPWR VPWR _08158_/A sky130_fd_sc_hd__buf_2
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05159_ input93/X _06696_/A input11/X _06698_/A VGND VGND VPWR VPWR _05159_/X sky130_fd_sc_hd__a22o_1
X_09967_ _10244_/CLK _09967_/D repeater403/X VGND VGND VPWR VPWR _09967_/Q sky130_fd_sc_hd__dfrtp_1
X_08918_ _08918_/A _08918_/B VGND VGND VPWR VPWR _08918_/X sky130_fd_sc_hd__and2_1
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09898_ _10268_/CLK _09898_/D repeater404/X VGND VGND VPWR VPWR _09898_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _08849_/A _08849_/B VGND VGND VPWR VPWR _09290_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10107_ _10482_/CLK _10107_/D repeater405/X VGND VGND VPWR VPWR _10107_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10038_ _10062_/CLK _10038_/D repeater410/X VGND VGND VPWR VPWR _10038_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06200_ _08019_/B VGND VGND VPWR VPWR _06200_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07180_ _07176_/Y _06087_/B _07177_/Y _06024_/B _07179_/X VGND VGND VPWR VPWR _07180_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06131_ _10020_/Q VGND VGND VPWR VPWR _06137_/A sky130_fd_sc_hd__inv_2
XFILLER_160_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06062_ _10066_/Q _06055_/X _09550_/A0 _06057_/X VGND VGND VPWR VPWR _10066_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05013_ _10440_/Q _05008_/X _09658_/A1 _05010_/X VGND VGND VPWR VPWR _10440_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09821_ _10364_/CLK _09821_/D repeater410/X VGND VGND VPWR VPWR _09821_/Q sky130_fd_sc_hd__dfstp_1
X_09752_ _09752_/CLK _09752_/D VGND VGND VPWR VPWR _09752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06964_ _10236_/Q VGND VGND VPWR VPWR _06964_/Y sky130_fd_sc_hd__inv_2
X_08703_ _08703_/A _08819_/B VGND VGND VPWR VPWR _09149_/B sky130_fd_sc_hd__or2_1
XFILLER_100_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09683_ _08355_/X _05491_/X _09683_/S VGND VGND VPWR VPWR _09683_/X sky130_fd_sc_hd__mux2_1
X_05915_ _10156_/Q _05911_/X _09660_/A1 _05912_/Y VGND VGND VPWR VPWR _10156_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06895_ _10017_/Q VGND VGND VPWR VPWR _06895_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08634_ _08634_/A _08634_/B _08641_/B VGND VGND VPWR VPWR _08888_/B sky130_fd_sc_hd__or3_2
X_05846_ _10197_/Q _05840_/X _09547_/A1 _05842_/X VGND VGND VPWR VPWR _10197_/D sky130_fd_sc_hd__a22o_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08565_ _08692_/C _08565_/B VGND VGND VPWR VPWR _08695_/C sky130_fd_sc_hd__or2_1
X_05777_ _05777_/A VGND VGND VPWR VPWR _05777_/Y sky130_fd_sc_hd__inv_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07516_ _07592_/A _07597_/C VGND VGND VPWR VPWR _07608_/B sky130_fd_sc_hd__or2_1
X_08496_ _08890_/A VGND VGND VPWR VPWR _08624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07447_ _07290_/X _07440_/A _09744_/Q _07441_/A VGND VGND VPWR VPWR _09744_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07378_ _10155_/Q VGND VGND VPWR VPWR _07378_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06329_ _06472_/A _06329_/B VGND VGND VPWR VPWR _06331_/A sky130_fd_sc_hd__or2_1
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09117_ _08674_/X _09109_/B _09114_/X _09116_/Y VGND VGND VPWR VPWR _09117_/X sky130_fd_sc_hd__o211a_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _09048_/A VGND VGND VPWR VPWR _09048_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06680_ _06680_/A VGND VGND VPWR VPWR _06681_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05700_ _05702_/A VGND VGND VPWR VPWR _05701_/A sky130_fd_sc_hd__inv_2
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05631_ _10322_/Q _05627_/X _09580_/X _05629_/X VGND VGND VPWR VPWR _10322_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08350_ _08349_/Y _08348_/Y _09813_/Q _09812_/Q VGND VGND VPWR VPWR _08350_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05562_ _06644_/A VGND VGND VPWR VPWR _05563_/A sky130_fd_sc_hd__clkbuf_1
X_07301_ input72/X _09699_/S _07300_/Y _06045_/B VGND VGND VPWR VPWR _07301_/X sky130_fd_sc_hd__o2bb2a_1
X_05493_ _05493_/A _05493_/B _05493_/C _05493_/D VGND VGND VPWR VPWR _05525_/S sky130_fd_sc_hd__or4_2
X_08281_ _07234_/Y _08186_/X _07244_/Y _08187_/X _08280_/X VGND VGND VPWR VPWR _08281_/X
+ sky130_fd_sc_hd__o221a_1
X_07232_ _10014_/Q VGND VGND VPWR VPWR _07232_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07163_ _10439_/Q _05091_/X _10434_/Q _05121_/Y VGND VGND VPWR VPWR _07163_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_06114_ _10034_/Q _06109_/X _09579_/X _06111_/X VGND VGND VPWR VPWR _10034_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _07092_/Y _06122_/B _07093_/Y _05775_/B VGND VGND VPWR VPWR _07094_/X sky130_fd_sc_hd__o22a_1
XFILLER_160_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06045_ _06087_/A _06045_/B VGND VGND VPWR VPWR _06047_/A sky130_fd_sc_hd__or2_1
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ net399_2/A _09804_/D _06612_/X VGND VGND VPWR VPWR _09804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07996_ _10005_/Q VGND VGND VPWR VPWR _08006_/A sky130_fd_sc_hd__inv_2
X_09735_ _09781_/CLK _09735_/D VGND VGND VPWR VPWR _09735_/Q sky130_fd_sc_hd__dfxtp_1
X_06947_ _06942_/Y _06205_/A _06943_/Y _05761_/A _06946_/X VGND VGND VPWR VPWR _06960_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09666_ _09806_/Q _09805_/Q _09773_/Q VGND VGND VPWR VPWR _09666_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08617_ _08847_/B VGND VGND VPWR VPWR _09057_/B sky130_fd_sc_hd__clkbuf_4
X_06878_ _06876_/Y _06206_/B _06877_/Y _06538_/B VGND VGND VPWR VPWR _06878_/X sky130_fd_sc_hd__o22a_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05829_ _05829_/A VGND VGND VPWR VPWR _05830_/B sky130_fd_sc_hd__buf_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09596_/X _09910_/Q _09776_/Q VGND VGND VPWR VPWR _09597_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08548_ _08548_/A VGND VGND VPWR VPWR _09278_/A sky130_fd_sc_hd__inv_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _08869_/A VGND VGND VPWR VPWR _09184_/A sky130_fd_sc_hd__inv_2
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10510_ _10510_/CLK _10510_/D repeater409/X VGND VGND VPWR VPWR _10510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10441_ _10478_/CLK _10441_/D repeater409/X VGND VGND VPWR VPWR _10441_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10372_ _10404_/CLK _10372_/D repeater410/X VGND VGND VPWR VPWR _10372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 _05406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _08679_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 input130/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _09487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07850_ _06710_/Y _07762_/X _06716_/Y _07811_/X _07849_/X VGND VGND VPWR VPWR _07859_/A
+ sky130_fd_sc_hd__o221a_1
X_07781_ _07781_/A VGND VGND VPWR VPWR _07781_/X sky130_fd_sc_hd__clkbuf_2
X_06801_ _06796_/Y _06313_/B _06797_/Y _06402_/B _06800_/X VGND VGND VPWR VPWR _06814_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04993_ _04993_/A _05130_/A VGND VGND VPWR VPWR _04995_/A sky130_fd_sc_hd__or2_2
X_09520_ _09520_/A VGND VGND VPWR VPWR _09520_/X sky130_fd_sc_hd__clkbuf_1
X_06732_ _06730_/Y _05896_/B _06731_/Y _06011_/B VGND VGND VPWR VPWR _06732_/X sky130_fd_sc_hd__o22a_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_8
X_06663_ _06663_/A VGND VGND VPWR VPWR _06664_/A sky130_fd_sc_hd__clkbuf_1
X_09451_ _09451_/A VGND VGND VPWR VPWR _09451_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08402_ _08402_/A _08402_/B _08402_/C _08402_/D VGND VGND VPWR VPWR _08406_/C sky130_fd_sc_hd__nand4_1
X_09382_ _09415_/C _09417_/D _09382_/C _09419_/A VGND VGND VPWR VPWR _09383_/C sky130_fd_sc_hd__or4_1
XFILLER_101_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06594_ _09808_/Q _06593_/Y _06589_/X VGND VGND VPWR VPWR _09808_/D sky130_fd_sc_hd__o21ba_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05614_ _10329_/Q _05605_/A _09536_/A3 _05606_/A VGND VGND VPWR VPWR _10329_/D sky130_fd_sc_hd__a22o_1
X_05545_ _10368_/Q _05542_/X _09658_/A1 _05543_/Y VGND VGND VPWR VPWR _10368_/D sky130_fd_sc_hd__a22o_1
X_08333_ _08333_/A VGND VGND VPWR VPWR _08335_/B sky130_fd_sc_hd__inv_2
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08264_ _07345_/Y _08183_/X _08261_/X _08263_/X VGND VGND VPWR VPWR _08274_/C sky130_fd_sc_hd__o211a_1
X_05476_ _05476_/A VGND VGND VPWR VPWR _05476_/Y sky130_fd_sc_hd__inv_2
X_07215_ _09794_/Q VGND VGND VPWR VPWR _07215_/Y sky130_fd_sc_hd__clkinv_2
X_08195_ _08195_/A VGND VGND VPWR VPWR _08195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07146_ _10010_/Q VGND VGND VPWR VPWR _07146_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07077_ _09836_/Q VGND VGND VPWR VPWR _09463_/A sky130_fd_sc_hd__inv_6
Xoutput362 _09745_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_126_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput340 _09557_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_2
Xoutput351 _10474_/Q VGND VGND VPWR VPWR sram_ro_addr[2] sky130_fd_sc_hd__buf_2
X_06028_ _10088_/Q _06025_/X _09581_/X _06027_/X VGND VGND VPWR VPWR _10088_/D sky130_fd_sc_hd__a22o_1
Xoutput384 _09741_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_160_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput373 _09755_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_113_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09718_ _10504_/Q _09489_/A VGND VGND VPWR VPWR _09718_/Z sky130_fd_sc_hd__ebufn_1
X_07979_ _07018_/Y _07532_/A _06992_/Y _07811_/A _07978_/X VGND VGND VPWR VPWR _07987_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_142_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ _08342_/X _09803_/Q _09773_/Q VGND VGND VPWR VPWR _09649_/X sky130_fd_sc_hd__mux2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10424_ _10406_/CLK _10424_/D _05059_/X VGND VGND VPWR VPWR _10424_/Q sky130_fd_sc_hd__dfrtn_1
X_10355_ _10355_/CLK _10355_/D repeater406/X VGND VGND VPWR VPWR _10355_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10288_/CLK _10286_/D repeater406/X VGND VGND VPWR VPWR _10286_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05330_ _05326_/Y _06392_/A _05328_/Y _06480_/A VGND VGND VPWR VPWR _05330_/X sky130_fd_sc_hd__o22a_1
XFILLER_186_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05261_ _05286_/B _05261_/B VGND VGND VPWR VPWR _05262_/A sky130_fd_sc_hd__or2_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05192_ _10076_/Q VGND VGND VPWR VPWR _05192_/Y sky130_fd_sc_hd__clkinv_2
X_07000_ _06998_/Y _05910_/B _06999_/Y _06529_/B VGND VGND VPWR VPWR _07000_/X sky130_fd_sc_hd__o22a_1
XFILLER_127_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08951_ _08951_/A _08951_/B VGND VGND VPWR VPWR _09201_/B sky130_fd_sc_hd__nor2_1
X_08882_ _08882_/A VGND VGND VPWR VPWR _09362_/B sky130_fd_sc_hd__inv_2
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07902_ _07362_/Y _07812_/X _07328_/Y _07813_/X VGND VGND VPWR VPWR _07902_/X sky130_fd_sc_hd__o22a_1
X_07833_ _07833_/A _07833_/B _07833_/C VGND VGND VPWR VPWR _07833_/Y sky130_fd_sc_hd__nand3_4
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07764_ _06881_/Y _07762_/X _06895_/Y _07651_/X _07763_/X VGND VGND VPWR VPWR _07775_/A
+ sky130_fd_sc_hd__o221a_1
X_04976_ _10459_/Q _04967_/A _09536_/A3 _04968_/A VGND VGND VPWR VPWR _10459_/D sky130_fd_sc_hd__a22o_1
X_09503_ _09503_/A VGND VGND VPWR VPWR _09504_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07695_ _07695_/A _07695_/B _07695_/C VGND VGND VPWR VPWR _07695_/Y sky130_fd_sc_hd__nand3_2
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06715_ _06715_/A _06715_/B _06708_/X _06714_/X VGND VGND VPWR VPWR _06758_/B sky130_fd_sc_hd__or4bb_1
X_06646_ _06646_/A VGND VGND VPWR VPWR _06655_/A sky130_fd_sc_hd__clkbuf_2
X_09434_ _09434_/A _09434_/B _09434_/C VGND VGND VPWR VPWR _09435_/B sky130_fd_sc_hd__or3_1
XFILLER_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _09350_/Y _09359_/Y _09361_/Y _09364_/X VGND VGND VPWR VPWR _09365_/X sky130_fd_sc_hd__a31o_1
X_06577_ _06591_/A VGND VGND VPWR VPWR _06578_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09296_ _09045_/C _09253_/B _09295_/Y _09035_/B _09086_/B VGND VGND VPWR VPWR _09390_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_138_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_30 _07278_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08316_ _06956_/Y _08188_/A _06998_/Y _08189_/A VGND VGND VPWR VPWR _08316_/X sky130_fd_sc_hd__o22a_1
X_05528_ _05603_/A _06708_/B VGND VGND VPWR VPWR _05530_/A sky130_fd_sc_hd__or2_2
XANTENNA_41 _07643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _09568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _09731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08247_ _05192_/Y _08195_/X _05254_/Y _08196_/X VGND VGND VPWR VPWR _08247_/X sky130_fd_sc_hd__o22a_1
X_05459_ _05459_/A VGND VGND VPWR VPWR _05460_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_74 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_96 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 input36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08178_ _08178_/A VGND VGND VPWR VPWR _08178_/X sky130_fd_sc_hd__buf_2
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _09467_/A _06480_/A _07128_/Y _05567_/B VGND VGND VPWR VPWR _07129_/X sky130_fd_sc_hd__o22a_1
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10140_ _10371_/CLK _10140_/D repeater410/X VGND VGND VPWR VPWR _10140_/Q sky130_fd_sc_hd__dfrtp_1
X_10071_ _10512_/CLK _10071_/D _07492_/B VGND VGND VPWR VPWR _10071_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10407_ _10411_/CLK _10407_/D repeater407/X VGND VGND VPWR VPWR _10407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _10510_/CLK _10338_/D repeater409/X VGND VGND VPWR VPWR _10338_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10504_/CLK _10269_/D repeater404/X VGND VGND VPWR VPWR _10269_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04830_ _04991_/A VGND VGND VPWR VPWR _05027_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06500_ _09850_/Q _06495_/X hold46/X _06496_/Y VGND VGND VPWR VPWR _09850_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07480_ _09778_/Q _06262_/B _07476_/Y _07479_/Y VGND VGND VPWR VPWR _09778_/D sky130_fd_sc_hd__a22o_1
X_06431_ _06432_/A VGND VGND VPWR VPWR _06431_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09150_ _08563_/A _09206_/A _08710_/A _08697_/B VGND VGND VPWR VPWR _09152_/A sky130_fd_sc_hd__o22ai_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06362_ _06362_/A VGND VGND VPWR VPWR _06363_/A sky130_fd_sc_hd__inv_2
X_09081_ _09081_/A _09294_/A _09390_/A _09358_/A VGND VGND VPWR VPWR _09086_/A sky130_fd_sc_hd__or4_1
X_06293_ _06293_/A VGND VGND VPWR VPWR _06294_/A sky130_fd_sc_hd__inv_2
X_05313_ _05313_/A _05349_/A VGND VGND VPWR VPWR _05314_/A sky130_fd_sc_hd__or2_1
X_08101_ _07264_/Y _08052_/X _07219_/Y _08053_/X _08100_/X VGND VGND VPWR VPWR _08117_/A
+ sky130_fd_sc_hd__o221a_1
X_05244_ _10365_/Q VGND VGND VPWR VPWR _05244_/Y sky130_fd_sc_hd__clkinv_2
X_08032_ _08032_/A _08032_/B _08038_/C VGND VGND VPWR VPWR _08200_/A sky130_fd_sc_hd__or3_4
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_6
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_6
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_4
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_6
Xinput94 sram_ro_data[10] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__clkbuf_2
X_05175_ _10071_/Q VGND VGND VPWR VPWR _05175_/Y sky130_fd_sc_hd__inv_2
X_09983_ _10288_/CLK _09983_/D repeater406/X VGND VGND VPWR VPWR _09983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08934_ _08934_/A _08957_/B VGND VGND VPWR VPWR _09286_/B sky130_fd_sc_hd__nor2_1
X_08865_ _09104_/A _09105_/B VGND VGND VPWR VPWR _08865_/X sky130_fd_sc_hd__or2_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08796_ _08485_/A _08795_/A _08644_/A _08795_/Y VGND VGND VPWR VPWR _08895_/B sky130_fd_sc_hd__a22o_1
XFILLER_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07816_ _07816_/A VGND VGND VPWR VPWR _07816_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07747_ _06868_/Y _07620_/X _07745_/Y _07621_/X _07746_/X VGND VGND VPWR VPWR _07747_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04959_ _04960_/B VGND VGND VPWR VPWR _04959_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07678_ _07226_/Y _07634_/X _07184_/Y _07635_/X VGND VGND VPWR VPWR _07678_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09417_ _09417_/A _09417_/B _09417_/C _09417_/D VGND VGND VPWR VPWR _09418_/D sky130_fd_sc_hd__or4_1
X_06629_ _09799_/Q _06605_/A _09644_/X _06606_/A VGND VGND VPWR VPWR _09799_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09348_ _09348_/A _09348_/B _09348_/C _09348_/D VGND VGND VPWR VPWR _09426_/C sky130_fd_sc_hd__or4_2
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09279_ _09352_/A _09278_/Y _09058_/A VGND VGND VPWR VPWR _09353_/B sky130_fd_sc_hd__o21ai_4
XFILLER_138_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10123_ _10127_/CLK _10123_/D _07492_/B VGND VGND VPWR VPWR _10123_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10054_ _10482_/CLK _10054_/D repeater405/X VGND VGND VPWR VPWR _10054_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _09951_/Q VGND VGND VPWR VPWR _06980_/Y sky130_fd_sc_hd__inv_2
X_05931_ _05931_/A VGND VGND VPWR VPWR _05931_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _08650_/A VGND VGND VPWR VPWR _09095_/A sky130_fd_sc_hd__buf_2
XFILLER_39_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05862_ _10186_/Q _05854_/A _09661_/A1 _05855_/A VGND VGND VPWR VPWR _10186_/D sky130_fd_sc_hd__a22o_1
X_07601_ _07601_/A _07601_/B VGND VGND VPWR VPWR _07817_/A sky130_fd_sc_hd__or2_4
X_04813_ _09670_/X VGND VGND VPWR VPWR _04991_/A sky130_fd_sc_hd__inv_2
X_05793_ _05793_/A VGND VGND VPWR VPWR _05794_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08581_ _08586_/A _08581_/B VGND VGND VPWR VPWR _09021_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07532_ _07532_/A VGND VGND VPWR VPWR _07533_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07463_ _10421_/Q _10274_/Q _05651_/B VGND VGND VPWR VPWR _09531_/A sky130_fd_sc_hd__o21ai_4
XFILLER_179_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09202_ _08620_/A _08761_/A _09372_/A _09204_/A _09046_/B VGND VGND VPWR VPWR _09306_/A
+ sky130_fd_sc_hd__a311oi_4
X_06414_ _06386_/X _09637_/X _09650_/X _09893_/Q VGND VGND VPWR VPWR _09893_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09133_ _09400_/A _09343_/A _09133_/C VGND VGND VPWR VPWR _09135_/A sky130_fd_sc_hd__or3_1
X_07394_ _10358_/Q VGND VGND VPWR VPWR _07394_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_175_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06345_ _09938_/Q _06340_/X _09579_/X _06342_/X VGND VGND VPWR VPWR _09938_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09064_ _09064_/A _09064_/B VGND VGND VPWR VPWR _09354_/C sky130_fd_sc_hd__or2_1
X_06276_ _09976_/Q _06269_/A _09660_/A1 _06270_/A VGND VGND VPWR VPWR _09976_/D sky130_fd_sc_hd__a22o_1
X_05227_ _09928_/Q VGND VGND VPWR VPWR _05227_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08015_ _08019_/B _08044_/B _08019_/C VGND VGND VPWR VPWR _08184_/A sky130_fd_sc_hd__or3_4
XFILLER_190_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05158_ _05163_/B _05261_/B VGND VGND VPWR VPWR _06698_/A sky130_fd_sc_hd__nor2_2
XFILLER_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09966_ _10244_/CLK _09966_/D repeater403/X VGND VGND VPWR VPWR _09966_/Q sky130_fd_sc_hd__dfrtp_1
X_05089_ _05089_/A VGND VGND VPWR VPWR _05089_/X sky130_fd_sc_hd__buf_2
X_08917_ _08927_/A _09011_/A _09057_/A VGND VGND VPWR VPWR _08918_/B sky130_fd_sc_hd__or3_1
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09897_ _10310_/CLK _09897_/D repeater404/X VGND VGND VPWR VPWR _09897_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _08848_/A _09073_/A VGND VGND VPWR VPWR _08850_/A sky130_fd_sc_hd__or2_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08779_ _08913_/B _08492_/A _08794_/B VGND VGND VPWR VPWR _08814_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10110_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10106_ _10283_/CLK _10106_/D repeater406/X VGND VGND VPWR VPWR _10106_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10037_ _10062_/CLK _10037_/D repeater410/X VGND VGND VPWR VPWR _10037_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06130_ _10022_/Q VGND VGND VPWR VPWR _06140_/B sky130_fd_sc_hd__inv_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06061_ _10067_/Q _06055_/X _09547_/A1 _06057_/X VGND VGND VPWR VPWR _10067_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05012_ _10441_/Q _05008_/X _09545_/A1 _05010_/X VGND VGND VPWR VPWR _10441_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09820_ _10405_/CLK _09820_/D repeater410/X VGND VGND VPWR VPWR _09820_/Q sky130_fd_sc_hd__dfstp_1
X_09751_ _09752_/CLK _09751_/D VGND VGND VPWR VPWR _09751_/Q sky130_fd_sc_hd__dfxtp_1
X_06963_ _10067_/Q VGND VGND VPWR VPWR _06963_/Y sky130_fd_sc_hd__inv_2
X_05914_ _10157_/Q _05911_/X _09550_/A0 _05912_/Y VGND VGND VPWR VPWR _10157_/D sky130_fd_sc_hd__a22o_1
X_08702_ _08717_/A _08819_/B VGND VGND VPWR VPWR _08704_/C sky130_fd_sc_hd__or2_1
XFILLER_100_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06894_ _10172_/Q VGND VGND VPWR VPWR _06894_/Y sky130_fd_sc_hd__inv_4
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09682_ _07617_/X _07506_/Y _09682_/S VGND VGND VPWR VPWR _09682_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08633_ _08633_/A _08789_/B VGND VGND VPWR VPWR _08641_/B sky130_fd_sc_hd__or2_1
X_05845_ _10198_/Q _05840_/X _09579_/X _05842_/X VGND VGND VPWR VPWR _10198_/D sky130_fd_sc_hd__a22o_1
X_08564_ _08564_/A VGND VGND VPWR VPWR _08692_/C sky130_fd_sc_hd__inv_2
X_05776_ _05777_/A VGND VGND VPWR VPWR _05776_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07515_ _07549_/B VGND VGND VPWR VPWR _07564_/C sky130_fd_sc_hd__clkbuf_1
X_08495_ _08794_/A VGND VGND VPWR VPWR _08890_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07446_ _07159_/X _07439_/X _09745_/Q _07441_/X VGND VGND VPWR VPWR _09745_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07377_ _10186_/Q VGND VGND VPWR VPWR _07377_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09116_ _09319_/B _09285_/A VGND VGND VPWR VPWR _09116_/Y sky130_fd_sc_hd__nor2_1
X_06328_ _06328_/A VGND VGND VPWR VPWR _06329_/B sky130_fd_sc_hd__buf_2
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09047_ _08806_/Y _08808_/X _09306_/B VGND VGND VPWR VPWR _09062_/A sky130_fd_sc_hd__a21o_1
XFILLER_190_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06259_ _09778_/Q _09554_/X VGND VGND VPWR VPWR _06259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09949_ _10062_/CLK _09949_/D repeater405/X VGND VGND VPWR VPWR _09949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05630_ _10323_/Q _05627_/X _09581_/X _05629_/X VGND VGND VPWR VPWR _10323_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05561_ _10357_/Q _05552_/A _09659_/A1 _05553_/A VGND VGND VPWR VPWR _10357_/D sky130_fd_sc_hd__a22o_1
X_07300_ _10072_/Q VGND VGND VPWR VPWR _07300_/Y sky130_fd_sc_hd__inv_2
X_05492_ _09534_/A _05489_/X _09533_/A _05491_/X VGND VGND VPWR VPWR _05493_/C sky130_fd_sc_hd__o22ai_1
X_08280_ _07212_/Y _08188_/X _07231_/Y _08189_/X VGND VGND VPWR VPWR _08280_/X sky130_fd_sc_hd__o22a_1
X_07231_ _10156_/Q VGND VGND VPWR VPWR _07231_/Y sky130_fd_sc_hd__inv_2
X_07162_ input94/X _05101_/X _10474_/Q _06933_/B _07161_/X VGND VGND VPWR VPWR _07167_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06113_ _10035_/Q _06109_/X _09580_/X _06111_/X VGND VGND VPWR VPWR _10035_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07093_ _10235_/Q VGND VGND VPWR VPWR _07093_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06044_ _10076_/Q _06038_/X _09574_/X _06039_/Y VGND VGND VPWR VPWR _10076_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09803_ _10406_/CLK _09803_/D _06615_/X VGND VGND VPWR VPWR _09803_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07995_ _08040_/A VGND VGND VPWR VPWR _08032_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09734_ _09781_/CLK _09734_/D VGND VGND VPWR VPWR _09734_/Q sky130_fd_sc_hd__dfxtp_1
X_06946_ _06944_/Y _06251_/B _06945_/Y _05541_/B VGND VGND VPWR VPWR _06946_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06877_ _09825_/Q VGND VGND VPWR VPWR _06877_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09665_ _09664_/X _10397_/Q _10299_/Q VGND VGND VPWR VPWR _09665_/X sky130_fd_sc_hd__mux2_1
X_05828_ _10206_/Q _05822_/X _09574_/X _05823_/Y VGND VGND VPWR VPWR _10206_/D sky130_fd_sc_hd__a22o_1
X_08616_ _08823_/B VGND VGND VPWR VPWR _08847_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _08153_/Y _10333_/Q _09700_/S VGND VGND VPWR VPWR _09596_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05759_ _10246_/Q _05751_/A _09661_/A1 _05752_/A VGND VGND VPWR VPWR _10246_/D sky130_fd_sc_hd__a22o_1
X_08547_ _09102_/D _08970_/A VGND VGND VPWR VPWR _08548_/A sky130_fd_sc_hd__or2_2
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08478_ _08757_/A _08970_/A VGND VGND VPWR VPWR _08869_/A sky130_fd_sc_hd__or2_1
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07429_ _06759_/X _07426_/X _09757_/Q _07428_/X VGND VGND VPWR VPWR _09757_/D sky130_fd_sc_hd__o22a_1
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10440_ _10478_/CLK _10440_/D _05034_/A VGND VGND VPWR VPWR _10440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10371_ _10371_/CLK _10371_/D repeater410/X VGND VGND VPWR VPWR _10371_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_191_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_120 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _05406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _09353_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_175 input131/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_186 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _07498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06800_ _06798_/Y _05576_/B _06799_/Y _06339_/B VGND VGND VPWR VPWR _06800_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07780_ _10087_/Q VGND VGND VPWR VPWR _07780_/Y sky130_fd_sc_hd__inv_2
X_04992_ _04992_/A _05155_/B VGND VGND VPWR VPWR _05130_/A sky130_fd_sc_hd__or2_1
X_06731_ _10096_/Q VGND VGND VPWR VPWR _06731_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09450_ _09450_/A VGND VGND VPWR VPWR _09450_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08401_ _08401_/A _08401_/B VGND VGND VPWR VPWR _08406_/B sky130_fd_sc_hd__nand2_1
X_06662_ _06662_/A VGND VGND VPWR VPWR _06662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09381_ _09425_/A _09415_/D _09418_/B VGND VGND VPWR VPWR _09382_/C sky130_fd_sc_hd__or3_1
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06593_ _06593_/A _06593_/B VGND VGND VPWR VPWR _06593_/Y sky130_fd_sc_hd__nor2_1
X_05613_ _10330_/Q _05605_/A _06684_/B1 _05606_/A VGND VGND VPWR VPWR _10330_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05544_ _10369_/Q _05542_/X _09545_/A1 _05543_/Y VGND VGND VPWR VPWR _10369_/D sky130_fd_sc_hd__a22o_1
X_08332_ _09800_/Q _09799_/Q _08333_/A VGND VGND VPWR VPWR _08332_/X sky130_fd_sc_hd__o21a_1
X_08263_ _07353_/Y _08186_/X _07414_/Y _08187_/X _08262_/X VGND VGND VPWR VPWR _08263_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07214_ _10104_/Q VGND VGND VPWR VPWR _07214_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05475_ _05476_/A VGND VGND VPWR VPWR _05475_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08194_ _08194_/A VGND VGND VPWR VPWR _08194_/X sky130_fd_sc_hd__clkbuf_2
X_07145_ _09823_/Q VGND VGND VPWR VPWR _09461_/A sky130_fd_sc_hd__inv_4
XFILLER_173_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07076_ _07071_/Y _05952_/B _09471_/A _06402_/B _07075_/X VGND VGND VPWR VPWR _07089_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput341 _09558_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_2
X_06027_ _06027_/A VGND VGND VPWR VPWR _06027_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput330 _10450_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_2
Xoutput352 _10475_/Q VGND VGND VPWR VPWR sram_ro_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_160_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput374 _09756_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput363 _09746_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput385 _09761_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07978_ _06944_/Y _07812_/A _06982_/Y _07653_/A VGND VGND VPWR VPWR _07978_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09717_ _10503_/Q _09487_/A VGND VGND VPWR VPWR _09717_/Z sky130_fd_sc_hd__ebufn_1
X_06929_ _10153_/Q VGND VGND VPWR VPWR _06929_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09648_ _08339_/X _09802_/Q _09773_/Q VGND VGND VPWR VPWR _09648_/X sky130_fd_sc_hd__mux2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10416_/Q _10383_/Q _10299_/Q VGND VGND VPWR VPWR _09579_/X sky130_fd_sc_hd__mux2_8
XFILLER_70_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10423_ _10406_/CLK _10423_/D _05062_/X VGND VGND VPWR VPWR _10423_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_167_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10354_ _10354_/CLK _10354_/D repeater406/X VGND VGND VPWR VPWR _10354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10285_ _10288_/CLK _10285_/D repeater406/X VGND VGND VPWR VPWR _10285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05260_ _09792_/Q VGND VGND VPWR VPWR _05260_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05191_ _05336_/A _05286_/B VGND VGND VPWR VPWR _05851_/A sky130_fd_sc_hd__or2_4
XFILLER_155_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08950_ _08950_/A _09289_/B VGND VGND VPWR VPWR _08952_/A sky130_fd_sc_hd__or2_1
X_08881_ _09044_/B VGND VGND VPWR VPWR _09384_/C sky130_fd_sc_hd__clkbuf_2
X_07901_ _07901_/A _07901_/B _07901_/C _07901_/D VGND VGND VPWR VPWR _07912_/B sky130_fd_sc_hd__and4_1
X_07832_ _07832_/A _07832_/B _07832_/C _07832_/D VGND VGND VPWR VPWR _07833_/C sky130_fd_sc_hd__and4_1
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09502_ _09502_/A VGND VGND VPWR VPWR _09502_/X sky130_fd_sc_hd__clkbuf_1
X_07763_ _06876_/Y _07652_/X _06865_/Y _07653_/X VGND VGND VPWR VPWR _07763_/X sky130_fd_sc_hd__o22a_1
X_04975_ _10460_/Q _04967_/A _06684_/B1 _04968_/A VGND VGND VPWR VPWR _10460_/D sky130_fd_sc_hd__a22o_1
X_06714_ _06709_/Y _06291_/B _06710_/Y _06481_/B _06713_/X VGND VGND VPWR VPWR _06714_/X
+ sky130_fd_sc_hd__o221a_2
X_07694_ _07694_/A _07694_/B _07694_/C _07694_/D VGND VGND VPWR VPWR _07695_/C sky130_fd_sc_hd__and4_1
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06645_ _06645_/A VGND VGND VPWR VPWR _06645_/X sky130_fd_sc_hd__clkbuf_1
X_09433_ _09433_/A _09433_/B _09433_/C _09433_/D VGND VGND VPWR VPWR _09434_/C sky130_fd_sc_hd__or4_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09364_ _09393_/A _09434_/B _09393_/C VGND VGND VPWR VPWR _09364_/X sky130_fd_sc_hd__or3_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08315_ _07011_/Y _08184_/A _06944_/Y _08158_/A VGND VGND VPWR VPWR _08315_/X sky130_fd_sc_hd__o22a_1
X_06576_ _06576_/A VGND VGND VPWR VPWR _09812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09295_ _09295_/A _09295_/B _09295_/C VGND VGND VPWR VPWR _09295_/Y sky130_fd_sc_hd__nor3_1
XANTENNA_31 _07278_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05527_ _05527_/A VGND VGND VPWR VPWR _06708_/B sky130_fd_sc_hd__buf_4
XANTENNA_20 _06997_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _09563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _09732_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05458_ _09696_/X _05449_/X _10395_/Q _05451_/X VGND VGND VPWR VPWR _10395_/D sky130_fd_sc_hd__a22o_1
X_08246_ _05339_/Y _08183_/X _08243_/X _08245_/X VGND VGND VPWR VPWR _08256_/C sky130_fd_sc_hd__o211a_1
XANTENNA_75 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_42 _07703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08177_ _08177_/A VGND VGND VPWR VPWR _08177_/X sky130_fd_sc_hd__buf_2
XANTENNA_97 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07128_ _10354_/Q VGND VGND VPWR VPWR _07128_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05389_ _09808_/Q _06593_/A VGND VGND VPWR VPWR _05389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07059_ _09931_/Q VGND VGND VPWR VPWR _07059_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10070_ _10350_/CLK _10070_/D repeater405/X VGND VGND VPWR VPWR _10070_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10406_ _10406_/CLK _10406_/D _05428_/X VGND VGND VPWR VPWR _10406_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10337_ _10341_/CLK _10337_/D repeater409/X VGND VGND VPWR VPWR _10337_/Q sky130_fd_sc_hd__dfrtp_1
X_10268_ _10268_/CLK _10268_/D repeater404/X VGND VGND VPWR VPWR _10268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10199_ _10289_/CLK _10199_/D repeater402/X VGND VGND VPWR VPWR _10199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06430_ _06472_/A _06430_/B VGND VGND VPWR VPWR _06432_/A sky130_fd_sc_hd__or2_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06361_ _06362_/A VGND VGND VPWR VPWR _06361_/X sky130_fd_sc_hd__clkbuf_2
X_09080_ _08900_/A _08977_/C _08978_/C VGND VGND VPWR VPWR _09358_/A sky130_fd_sc_hd__o21ai_1
X_06292_ _06293_/A VGND VGND VPWR VPWR _06292_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05312_ _10253_/Q VGND VGND VPWR VPWR _05312_/Y sky130_fd_sc_hd__inv_2
X_08100_ _07227_/Y _08054_/X _07202_/Y _08055_/X VGND VGND VPWR VPWR _08100_/X sky130_fd_sc_hd__o22a_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_6
X_05243_ _05305_/B _05307_/B VGND VGND VPWR VPWR _06153_/A sky130_fd_sc_hd__or2_4
X_08031_ _08037_/B _08032_/A _10006_/Q VGND VGND VPWR VPWR _08199_/A sky130_fd_sc_hd__or3_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_6
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_6
XFILLER_162_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__clkbuf_2
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_6
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05174_ _06692_/A VGND VGND VPWR VPWR _06024_/B sky130_fd_sc_hd__buf_2
Xinput95 sram_ro_data[11] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09982_ _10023_/CLK _09982_/D _05034_/A VGND VGND VPWR VPWR _09982_/Q sky130_fd_sc_hd__dfrtp_1
X_08933_ _08933_/A VGND VGND VPWR VPWR _08957_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08864_ _08864_/A _09095_/A VGND VGND VPWR VPWR _09104_/A sky130_fd_sc_hd__or2_1
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08795_ _08795_/A VGND VGND VPWR VPWR _08795_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07815_ _06791_/Y _07762_/X _06816_/Y _07811_/X _07814_/X VGND VGND VPWR VPWR _07832_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07746_ _06871_/Y _07622_/X _06869_/Y _07623_/X VGND VGND VPWR VPWR _07746_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04958_ _05118_/A _05305_/B VGND VGND VPWR VPWR _04960_/B sky130_fd_sc_hd__or2_1
X_09416_ _09416_/A _09416_/B VGND VGND VPWR VPWR _09417_/C sky130_fd_sc_hd__or2_1
X_04889_ _04889_/A VGND VGND VPWR VPWR _04889_/X sky130_fd_sc_hd__clkbuf_2
X_07677_ _07197_/Y _07627_/X _07259_/Y _07628_/X _07676_/X VGND VGND VPWR VPWR _07684_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06628_ _06628_/A VGND VGND VPWR VPWR _06628_/X sky130_fd_sc_hd__clkbuf_1
X_09347_ _09425_/B _09426_/A VGND VGND VPWR VPWR _09347_/Y sky130_fd_sc_hd__nor2_1
X_06559_ _06568_/A VGND VGND VPWR VPWR _06560_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09278_ _09278_/A _09278_/B VGND VGND VPWR VPWR _09278_/Y sky130_fd_sc_hd__nor2_1
X_08229_ _06731_/Y _08195_/X _06746_/Y _08196_/X VGND VGND VPWR VPWR _08229_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10122_ _10289_/CLK _10122_/D repeater402/X VGND VGND VPWR VPWR _10122_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10053_ _10110_/CLK _10053_/D repeater405/X VGND VGND VPWR VPWR _10053_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _05930_/A VGND VGND VPWR VPWR _05931_/A sky130_fd_sc_hd__inv_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05861_ _10187_/Q _05854_/A _09660_/A1 _05855_/A VGND VGND VPWR VPWR _10187_/D sky130_fd_sc_hd__a22o_1
X_04812_ _10271_/Q _05179_/A _10513_/Q VGND VGND VPWR VPWR _09712_/A sky130_fd_sc_hd__mux2_1
X_07600_ _07600_/A VGND VGND VPWR VPWR _07816_/A sky130_fd_sc_hd__buf_2
X_08580_ _08583_/A _08581_/B _09010_/A _09020_/A _08579_/X VGND VGND VPWR VPWR _08584_/B
+ sky130_fd_sc_hd__o221ai_1
X_05792_ _10227_/Q _05786_/X _09574_/X _05787_/Y VGND VGND VPWR VPWR _10227_/D sky130_fd_sc_hd__a22o_1
X_07531_ _07762_/A VGND VGND VPWR VPWR _07532_/A sky130_fd_sc_hd__clkbuf_2
X_07462_ _10136_/Q VGND VGND VPWR VPWR _09517_/A sky130_fd_sc_hd__clkinv_8
XFILLER_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06413_ _09894_/Q _06404_/A _09659_/A1 _06405_/A VGND VGND VPWR VPWR _09894_/D sky130_fd_sc_hd__a22o_1
X_07393_ _07393_/A _07393_/B _07393_/C VGND VGND VPWR VPWR _07419_/C sky130_fd_sc_hd__and3_1
X_09201_ _09326_/A _09201_/B _09201_/C VGND VGND VPWR VPWR _09369_/C sky130_fd_sc_hd__or3_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06344_ _09939_/Q _06340_/X _09580_/X _06342_/X VGND VGND VPWR VPWR _09939_/D sky130_fd_sc_hd__a22o_1
X_09132_ _08860_/A _09099_/X _09131_/X VGND VGND VPWR VPWR _09133_/C sky130_fd_sc_hd__o21bai_1
XFILLER_187_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09063_ _09063_/A _09370_/B VGND VGND VPWR VPWR _09285_/C sky130_fd_sc_hd__or2_1
X_06275_ _09977_/Q _06268_/X _09550_/A0 _06270_/X VGND VGND VPWR VPWR _09977_/D sky130_fd_sc_hd__a22o_1
X_05226_ _05305_/B _05275_/B VGND VGND VPWR VPWR _06438_/A sky130_fd_sc_hd__or2_4
X_08014_ _08038_/A _08032_/B _10006_/Q VGND VGND VPWR VPWR _08183_/A sky130_fd_sc_hd__or3_4
X_05157_ _05157_/A _05292_/A VGND VGND VPWR VPWR _06696_/A sky130_fd_sc_hd__nor2_2
XFILLER_190_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09965_ _10244_/CLK _09965_/D repeater403/X VGND VGND VPWR VPWR _09965_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05088_ _05088_/A VGND VGND VPWR VPWR _05089_/A sky130_fd_sc_hd__clkinv_2
X_08916_ _08916_/A _09011_/A _09057_/A VGND VGND VPWR VPWR _08918_/A sky130_fd_sc_hd__or3_1
X_09896_ _10268_/CLK _09896_/D repeater404/X VGND VGND VPWR VPWR _09896_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08847_ _08849_/B _08847_/B VGND VGND VPWR VPWR _09073_/A sky130_fd_sc_hd__nor2_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08778_ _08883_/B _09093_/A VGND VGND VPWR VPWR _09141_/B sky130_fd_sc_hd__nor2_1
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _10397_/CLK sky130_fd_sc_hd__clkbuf_2
X_07729_ _07726_/Y _07639_/X _07727_/Y _07641_/X _07728_/X VGND VGND VPWR VPWR _07732_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10105_ _10283_/CLK _10105_/D repeater406/X VGND VGND VPWR VPWR _10105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10036_ _10135_/CLK _10036_/D _07492_/B VGND VGND VPWR VPWR _10036_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06060_ _10068_/Q _06055_/X _09579_/X _06057_/X VGND VGND VPWR VPWR _10068_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05011_ _10442_/Q _05008_/X _09579_/X _05010_/X VGND VGND VPWR VPWR _10442_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09750_ _09781_/CLK _09750_/D VGND VGND VPWR VPWR _09750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06962_ _10145_/Q VGND VGND VPWR VPWR _06962_/Y sky130_fd_sc_hd__clkinv_4
X_05913_ _10158_/Q _05911_/X _09578_/X _05912_/Y VGND VGND VPWR VPWR _10158_/D sky130_fd_sc_hd__a22o_1
X_08701_ _08701_/A VGND VGND VPWR VPWR _08717_/A sky130_fd_sc_hd__buf_2
X_09681_ _09807_/Q _09809_/Q _09808_/Q VGND VGND VPWR VPWR _09681_/X sky130_fd_sc_hd__mux2_1
X_08632_ _08634_/B _08884_/A _08789_/B VGND VGND VPWR VPWR _08890_/B sky130_fd_sc_hd__or3_1
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06893_ _06893_/A _06893_/B VGND VGND VPWR VPWR _06893_/X sky130_fd_sc_hd__or2_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05844_ _10199_/Q _05840_/X _09580_/X _05842_/X VGND VGND VPWR VPWR _10199_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05775_ _05775_/A _05775_/B VGND VGND VPWR VPWR _05777_/A sky130_fd_sc_hd__or2_1
X_08563_ _08563_/A _09012_/A VGND VGND VPWR VPWR _08563_/X sky130_fd_sc_hd__or2_1
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08494_ _08494_/A VGND VGND VPWR VPWR _08794_/A sky130_fd_sc_hd__inv_2
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07514_ _07554_/C VGND VGND VPWR VPWR _07549_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07445_ _07030_/X _07439_/X _09746_/Q _07441_/X VGND VGND VPWR VPWR _09746_/D sky130_fd_sc_hd__o22a_2
XFILLER_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07376_ _10168_/Q VGND VGND VPWR VPWR _07376_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06327_ _06327_/A VGND VGND VPWR VPWR _06472_/A sky130_fd_sc_hd__buf_2
X_09115_ _09115_/A VGND VGND VPWR VPWR _09319_/B sky130_fd_sc_hd__inv_2
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06258_ _09983_/Q _06252_/X _09574_/X _06253_/Y VGND VGND VPWR VPWR _09983_/D sky130_fd_sc_hd__a22o_1
X_09046_ _09046_/A _09046_/B _09103_/A VGND VGND VPWR VPWR _09306_/B sky130_fd_sc_hd__nor3_1
XFILLER_190_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05209_ _05313_/A _05333_/A VGND VGND VPWR VPWR _05774_/A sky130_fd_sc_hd__or2_1
XFILLER_163_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06189_ _10006_/Q _06177_/Y _06184_/Y _06147_/X _06188_/X VGND VGND VPWR VPWR _10006_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09948_ _10110_/CLK _09948_/D repeater405/X VGND VGND VPWR VPWR _09948_/Q sky130_fd_sc_hd__dfstp_1
X_09879_ _10409_/CLK _09879_/D repeater407/X VGND VGND VPWR VPWR _09879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ _10495_/CLK _10019_/D repeater404/X VGND VGND VPWR VPWR _10019_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05560_ _10358_/Q _05552_/A _09661_/A1 _05553_/A VGND VGND VPWR VPWR _10358_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05491_ _05491_/A VGND VGND VPWR VPWR _05491_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07230_ _07225_/Y _05852_/B _07226_/Y _05882_/A _07229_/X VGND VGND VPWR VPWR _07243_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07161_ input130/X _05118_/Y _10485_/Q _06633_/A VGND VGND VPWR VPWR _07161_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06112_ _10036_/Q _06109_/X _09581_/X _06111_/X VGND VGND VPWR VPWR _10036_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07092_ _10027_/Q VGND VGND VPWR VPWR _07092_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_160_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06043_ _10077_/Q _06038_/X _06684_/B1 _06039_/Y VGND VGND VPWR VPWR _10077_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_42_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09802_ net399_2/A _09802_/D _06619_/X VGND VGND VPWR VPWR _09802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07994_ _10003_/Q _07994_/B VGND VGND VPWR VPWR _08040_/A sky130_fd_sc_hd__or2_1
X_09733_ _10285_/Q _09519_/A VGND VGND VPWR VPWR _09733_/Z sky130_fd_sc_hd__ebufn_2
X_06945_ _10369_/Q VGND VGND VPWR VPWR _06945_/Y sky130_fd_sc_hd__inv_2
X_06876_ _09999_/Q VGND VGND VPWR VPWR _06876_/Y sky130_fd_sc_hd__inv_2
X_09664_ _09805_/Q _09804_/Q _09773_/Q VGND VGND VPWR VPWR _09664_/X sky130_fd_sc_hd__mux2_1
X_08615_ _09085_/D _09085_/B _08768_/C VGND VGND VPWR VPWR _08823_/B sky130_fd_sc_hd__or3_4
X_05827_ _10207_/Q _05822_/X _09661_/A1 _05823_/Y VGND VGND VPWR VPWR _10207_/D sky130_fd_sc_hd__a22o_1
X_09595_ _09594_/X _09909_/Q _09776_/Q VGND VGND VPWR VPWR _09595_/X sky130_fd_sc_hd__mux2_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05758_ _10247_/Q _05751_/A _09660_/A1 _05752_/A VGND VGND VPWR VPWR _10247_/D sky130_fd_sc_hd__a22o_1
X_08546_ _08546_/A _08546_/B VGND VGND VPWR VPWR _08546_/Y sky130_fd_sc_hd__nor2_1
X_08477_ _09247_/C _08567_/A _08774_/A VGND VGND VPWR VPWR _08757_/A sky130_fd_sc_hd__or3_2
XFILLER_145_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05689_ _06679_/A _05689_/B VGND VGND VPWR VPWR _05691_/A sky130_fd_sc_hd__or2_4
X_07428_ _07428_/A VGND VGND VPWR VPWR _07428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07359_ _10142_/Q VGND VGND VPWR VPWR _07359_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10370_ _10371_/CLK _10370_/D repeater410/X VGND VGND VPWR VPWR _10370_/Q sky130_fd_sc_hd__dfstp_1
X_09029_ _09029_/A _09206_/B VGND VGND VPWR VPWR _09214_/C sky130_fd_sc_hd__nor2_1
XFILLER_104_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 _07505_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _09481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 _10479_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 _06096_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10499_ _10500_/CLK _10499_/D repeater407/X VGND VGND VPWR VPWR _10499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04991_ _04991_/A _04991_/B _05082_/A _09676_/X VGND VGND VPWR VPWR _05155_/B sky130_fd_sc_hd__or4_2
X_06730_ _10166_/Q VGND VGND VPWR VPWR _06730_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06661_ _06663_/A VGND VGND VPWR VPWR _06662_/A sky130_fd_sc_hd__clkbuf_1
X_08400_ _09236_/A VGND VGND VPWR VPWR _08426_/A sky130_fd_sc_hd__inv_2
XFILLER_91_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05612_ _10331_/Q _05605_/A _06683_/B1 _05606_/A VGND VGND VPWR VPWR _10331_/D sky130_fd_sc_hd__a22o_1
X_09380_ _09380_/A _09380_/B _09380_/C _09380_/D VGND VGND VPWR VPWR _09411_/D sky130_fd_sc_hd__or4_4
X_06592_ _06592_/A VGND VGND VPWR VPWR _06592_/X sky130_fd_sc_hd__clkbuf_1
X_05543_ _05543_/A VGND VGND VPWR VPWR _05543_/Y sky130_fd_sc_hd__inv_2
X_08331_ _09800_/Q _09799_/Q VGND VGND VPWR VPWR _08333_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08262_ _07358_/Y _08188_/X _07378_/Y _08189_/X VGND VGND VPWR VPWR _08262_/X sky130_fd_sc_hd__o22a_1
X_05474_ _05541_/A _05474_/B VGND VGND VPWR VPWR _05476_/A sky130_fd_sc_hd__or2_1
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07213_ _10208_/Q VGND VGND VPWR VPWR _07213_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_118_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08193_ _08193_/A VGND VGND VPWR VPWR _08193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07144_ _10373_/Q VGND VGND VPWR VPWR _09455_/A sky130_fd_sc_hd__clkinv_4
XFILLER_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07075_ _07073_/Y _05865_/B _07074_/Y _05910_/B VGND VGND VPWR VPWR _07075_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput353 _10476_/Q VGND VGND VPWR VPWR sram_ro_addr[4] sky130_fd_sc_hd__buf_2
X_06026_ _06026_/A VGND VGND VPWR VPWR _06027_/A sky130_fd_sc_hd__inv_2
Xoutput342 _09555_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_2
Xoutput331 _10451_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_2
Xoutput320 _10464_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_2
Xoutput375 _09757_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput364 _09747_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput386 _09762_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07977_ _07977_/A _07977_/B _07977_/C _07977_/D VGND VGND VPWR VPWR _07988_/B sky130_fd_sc_hd__and4_1
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09716_ _10502_/Q _09485_/A VGND VGND VPWR VPWR _09716_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06928_ _10257_/Q VGND VGND VPWR VPWR _06928_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06859_ _10250_/Q VGND VGND VPWR VPWR _06859_/Y sky130_fd_sc_hd__clkinv_4
X_09647_ _08337_/Y _09801_/Q _09773_/Q VGND VGND VPWR VPWR _09647_/X sky130_fd_sc_hd__mux2_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ hold45/X _10382_/Q _10299_/Q VGND VGND VPWR VPWR _09578_/X sky130_fd_sc_hd__mux2_8
XFILLER_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08529_/A VGND VGND VPWR VPWR _09010_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10422_ _10406_/CLK _10422_/D _05065_/X VGND VGND VPWR VPWR _10422_/Q sky130_fd_sc_hd__dfrtn_1
X_10353_ _10353_/CLK _10353_/D repeater406/X VGND VGND VPWR VPWR _10353_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_151_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10284_ _10288_/CLK _10284_/D repeater406/X VGND VGND VPWR VPWR _10284_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05190_ _05318_/B VGND VGND VPWR VPWR _05286_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08880_ _08880_/A VGND VGND VPWR VPWR _09044_/B sky130_fd_sc_hd__inv_2
X_07900_ _07351_/Y _07805_/X _07898_/Y _07758_/X _07899_/X VGND VGND VPWR VPWR _07901_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07831_ _06822_/Y _07825_/X _07826_/Y _07827_/X _07830_/X VGND VGND VPWR VPWR _07832_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09501_ _09501_/A VGND VGND VPWR VPWR _09502_/A sky130_fd_sc_hd__clkbuf_1
X_07762_ _07762_/A VGND VGND VPWR VPWR _07762_/X sky130_fd_sc_hd__buf_2
X_04974_ _10461_/Q _04967_/A _06683_/B1 _04968_/A VGND VGND VPWR VPWR _10461_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06713_ _06711_/Y _06338_/A _06712_/Y _06516_/B VGND VGND VPWR VPWR _06713_/X sky130_fd_sc_hd__o22a_1
X_07693_ _07237_/Y _07665_/X _07188_/Y _07666_/X _07692_/X VGND VGND VPWR VPWR _07694_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06644_ _06644_/A VGND VGND VPWR VPWR _06645_/A sky130_fd_sc_hd__clkbuf_1
X_09432_ _09432_/A _09432_/B _09432_/C VGND VGND VPWR VPWR _09433_/D sky130_fd_sc_hd__or3_1
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09363_ _09363_/A _09363_/B VGND VGND VPWR VPWR _09393_/C sky130_fd_sc_hd__or2_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06575_ _09653_/X _09812_/Q _06575_/S VGND VGND VPWR VPWR _06576_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05526_ _05526_/A VGND VGND VPWR VPWR _10378_/D sky130_fd_sc_hd__clkbuf_1
X_08314_ _07015_/Y _08177_/A _06955_/Y _08178_/A _08313_/X VGND VGND VPWR VPWR _08328_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09294_ _09294_/A _09294_/B VGND VGND VPWR VPWR _09358_/B sky130_fd_sc_hd__or2_1
XANTENNA_32 _07278_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _07881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _07028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _09564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _05179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05457_ _05457_/A VGND VGND VPWR VPWR _05457_/X sky130_fd_sc_hd__clkbuf_1
X_08245_ _05358_/Y _08186_/X _05282_/Y _08187_/X _08244_/X VGND VGND VPWR VPWR _08245_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_43 _07728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _06784_/Y _08052_/X _06796_/Y _08053_/X _08175_/X VGND VGND VPWR VPWR _08218_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA_98 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05388_ _06579_/B VGND VGND VPWR VPWR _06593_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_87 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07127_ _09857_/Q VGND VGND VPWR VPWR _09467_/A sky130_fd_sc_hd__clkinv_4
XFILLER_4_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07058_ _10196_/Q VGND VGND VPWR VPWR _09499_/A sky130_fd_sc_hd__inv_6
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06009_ _10097_/Q _06003_/X _09536_/A3 _06004_/Y VGND VGND VPWR VPWR _10097_/D sky130_fd_sc_hd__a22o_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10405_ _10405_/CLK _10405_/D hold41/X VGND VGND VPWR VPWR _10405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ _10336_/CLK _10336_/D repeater409/X VGND VGND VPWR VPWR _10336_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10267_ _10268_/CLK _10267_/D repeater404/X VGND VGND VPWR VPWR _10267_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10198_ _10289_/CLK _10198_/D repeater402/X VGND VGND VPWR VPWR _10198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06360_ _06481_/A _06360_/B VGND VGND VPWR VPWR _06362_/A sky130_fd_sc_hd__or2_2
XFILLER_174_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06291_ _06313_/A _06291_/B VGND VGND VPWR VPWR _06293_/A sky130_fd_sc_hd__or2_2
X_05311_ _05357_/A _05311_/B VGND VGND VPWR VPWR _06053_/A sky130_fd_sc_hd__or2_2
XFILLER_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05242_ _05299_/B VGND VGND VPWR VPWR _05307_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08030_ _05237_/Y _08193_/A _05285_/Y _08194_/A _08029_/X VGND VGND VPWR VPWR _08049_/A
+ sky130_fd_sc_hd__o221a_1
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__buf_12
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_6
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_4
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_6
XFILLER_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__clkbuf_4
X_05173_ _06630_/A _05173_/B VGND VGND VPWR VPWR _06692_/A sky130_fd_sc_hd__or2_1
Xinput96 sram_ro_data[12] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09981_ _10350_/CLK _09981_/D repeater405/X VGND VGND VPWR VPWR _09981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08932_ _08932_/A _09064_/B _09354_/B _09065_/B VGND VGND VPWR VPWR _08937_/A sky130_fd_sc_hd__or4_1
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08863_ _08863_/A VGND VGND VPWR VPWR _09079_/A sky130_fd_sc_hd__inv_2
X_08794_ _08794_/A _08794_/B VGND VGND VPWR VPWR _08795_/A sky130_fd_sc_hd__or2_1
X_07814_ _06793_/Y _07812_/X _06804_/Y _07813_/X VGND VGND VPWR VPWR _07814_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07745_ _10086_/Q VGND VGND VPWR VPWR _07745_/Y sky130_fd_sc_hd__inv_2
X_04957_ _05103_/B VGND VGND VPWR VPWR _05305_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09415_ _09415_/A _09415_/B _09415_/C _09415_/D VGND VGND VPWR VPWR _09418_/C sky130_fd_sc_hd__or4_1
X_04888_ _04888_/A VGND VGND VPWR VPWR _04889_/A sky130_fd_sc_hd__inv_2
X_07676_ _07195_/Y _07533_/C _07283_/Y _07629_/X VGND VGND VPWR VPWR _07676_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06627_ _06666_/A VGND VGND VPWR VPWR _06628_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06558_ _09815_/Q _06552_/X _09659_/A1 _06553_/Y VGND VGND VPWR VPWR _09815_/D sky130_fd_sc_hd__a22o_1
X_09346_ _09253_/A _08782_/Y _09299_/A _09139_/A VGND VGND VPWR VPWR _09426_/A sky130_fd_sc_hd__a211o_2
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05509_ _05509_/A VGND VGND VPWR VPWR _10382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09277_ _09277_/A VGND VGND VPWR VPWR _09352_/A sky130_fd_sc_hd__buf_2
X_06489_ _09857_/Q _06482_/X _09550_/A0 _06484_/X VGND VGND VPWR VPWR _09857_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08228_ _06741_/Y _08183_/X _08225_/X _08227_/X VGND VGND VPWR VPWR _08238_/C sky130_fd_sc_hd__o211a_1
XFILLER_153_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08159_ _06886_/Y _08065_/X _06876_/Y _08158_/X VGND VGND VPWR VPWR _08159_/X sky130_fd_sc_hd__o22a_1
XFILLER_180_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10121_ _10289_/CLK _10121_/D repeater402/X VGND VGND VPWR VPWR _10121_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10052_ _10482_/CLK _10052_/D repeater405/X VGND VGND VPWR VPWR _10052_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10319_ _10405_/CLK _10319_/D hold41/X VGND VGND VPWR VPWR _10319_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537__412 VGND VGND VPWR VPWR _09779_/D _09537__412/LO sky130_fd_sc_hd__conb_1
XFILLER_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05860_ _10188_/Q _05853_/X _09658_/A1 _05855_/X VGND VGND VPWR VPWR _10188_/D sky130_fd_sc_hd__a22o_1
X_05791_ _10228_/Q _05786_/X _09661_/A1 _05787_/Y VGND VGND VPWR VPWR _10228_/D sky130_fd_sc_hd__a22o_1
X_04811_ _10272_/Q _04811_/A1 _10512_/Q VGND VGND VPWR VPWR _09713_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07530_ _09989_/Q _09988_/Q _07602_/C _07562_/B VGND VGND VPWR VPWR _07762_/A sky130_fd_sc_hd__or4_1
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07461_ _05367_/X _07452_/A _09734_/Q _07453_/A VGND VGND VPWR VPWR _09734_/D sky130_fd_sc_hd__o22a_1
XFILLER_179_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06412_ _09895_/Q _06404_/A _09661_/A1 _06405_/A VGND VGND VPWR VPWR _09895_/D sky130_fd_sc_hd__a22o_1
X_07392_ _07387_/Y _06516_/B _07388_/Y _06393_/B _07391_/X VGND VGND VPWR VPWR _07393_/C
+ sky130_fd_sc_hd__o221a_1
X_09200_ _09200_/A VGND VGND VPWR VPWR _09326_/A sky130_fd_sc_hd__inv_2
XFILLER_148_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06343_ _09940_/Q _06340_/X _09581_/X _06342_/X VGND VGND VPWR VPWR _09940_/D sky130_fd_sc_hd__a22o_1
X_09131_ _09420_/A _09420_/B _09130_/X VGND VGND VPWR VPWR _09131_/X sky130_fd_sc_hd__or3b_1
X_09062_ _09062_/A _09062_/B _09283_/C _09389_/A VGND VGND VPWR VPWR _09066_/A sky130_fd_sc_hd__or4_1
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06274_ _09978_/Q _06268_/X _09547_/A1 _06270_/X VGND VGND VPWR VPWR _09978_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05225_ _09868_/Q VGND VGND VPWR VPWR _05225_/Y sky130_fd_sc_hd__inv_4
X_08013_ _05322_/Y _08177_/A _05248_/Y _08178_/A _08012_/X VGND VGND VPWR VPWR _08050_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05156_ _05615_/B VGND VGND VPWR VPWR _05156_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09964_ _10244_/CLK _09964_/D repeater403/X VGND VGND VPWR VPWR _09964_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05087_ _10029_/Q _05080_/X _10472_/Q _06776_/A _05086_/X VGND VGND VPWR VPWR _05108_/B
+ sky130_fd_sc_hd__a221o_1
X_08915_ _08689_/A _08909_/Y _08912_/Y _08801_/C _08914_/Y VGND VGND VPWR VPWR _08919_/C
+ sky130_fd_sc_hd__o32a_1
X_09895_ _10495_/CLK _09895_/D repeater404/X VGND VGND VPWR VPWR _09895_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_85_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08846_ _08846_/A _09386_/A VGND VGND VPWR VPWR _08848_/A sky130_fd_sc_hd__or2_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08777_ _09222_/B _08776_/Y VGND VGND VPWR VPWR _08994_/A sky130_fd_sc_hd__or2b_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05989_ _10109_/Q _05982_/A _06683_/B1 _05983_/A VGND VGND VPWR VPWR _10109_/D sky130_fd_sc_hd__a22o_1
X_07728_ _06968_/Y _07568_/B _06932_/Y _07642_/X VGND VGND VPWR VPWR _07728_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07659_ _07659_/A VGND VGND VPWR VPWR _07659_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09329_ _09329_/A _09329_/B VGND VGND VPWR VPWR _09419_/A sky130_fd_sc_hd__or2_1
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10104_ _10283_/CLK _10104_/D repeater406/X VGND VGND VPWR VPWR _10104_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10035_ _10135_/CLK _10035_/D _07492_/B VGND VGND VPWR VPWR _10035_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05010_ _05010_/A VGND VGND VPWR VPWR _05010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06961_ _10492_/Q VGND VGND VPWR VPWR _06961_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05912_ _05912_/A VGND VGND VPWR VPWR _05912_/Y sky130_fd_sc_hd__inv_2
X_08700_ _08700_/A _08700_/B _08700_/C _08700_/D VGND VGND VPWR VPWR _08700_/X sky130_fd_sc_hd__or4_1
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
X_09680_ _06581_/S _05390_/X _09680_/S VGND VGND VPWR VPWR _09680_/X sky130_fd_sc_hd__mux2_1
X_08631_ _08631_/A _08631_/B _08631_/C VGND VGND VPWR VPWR _08789_/B sky130_fd_sc_hd__or3_2
X_06892_ _10068_/Q VGND VGND VPWR VPWR _06893_/A sky130_fd_sc_hd__inv_2
X_05843_ _10200_/Q _05840_/X _09581_/X _05842_/X VGND VGND VPWR VPWR _10200_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08562_ _08911_/B VGND VGND VPWR VPWR _09012_/A sky130_fd_sc_hd__clkbuf_2
X_05774_ _05774_/A VGND VGND VPWR VPWR _05775_/B sky130_fd_sc_hd__buf_4
XFILLER_81_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08493_ _09085_/D _08493_/B _09102_/D _08546_/A VGND VGND VPWR VPWR _08998_/A sky130_fd_sc_hd__or4_1
X_07513_ _09993_/Q _09992_/Q VGND VGND VPWR VPWR _07554_/C sky130_fd_sc_hd__or2_1
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07444_ _06906_/X _07439_/X _09747_/Q _07441_/X VGND VGND VPWR VPWR _09747_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07375_ _09995_/Q VGND VGND VPWR VPWR _07375_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09114_ _08678_/X _09109_/B _09110_/X _09113_/Y VGND VGND VPWR VPWR _09114_/X sky130_fd_sc_hd__o211a_1
X_06326_ _09797_/Q _09775_/Q _06133_/Y _06325_/X VGND VGND VPWR VPWR _09946_/D sky130_fd_sc_hd__a31o_1
XFILLER_163_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06257_ _09984_/Q _06252_/X hold46/X _06253_/Y VGND VGND VPWR VPWR _09984_/D sky130_fd_sc_hd__a22o_1
X_09045_ _08768_/C _09045_/B _09045_/C _09102_/A VGND VGND VPWR VPWR _09434_/A sky130_fd_sc_hd__and4b_1
XFILLER_163_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05208_ _10232_/Q VGND VGND VPWR VPWR _05208_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06188_ _08016_/A VGND VGND VPWR VPWR _06188_/X sky130_fd_sc_hd__buf_2
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05139_ _05327_/A _05139_/B VGND VGND VPWR VPWR _05139_/X sky130_fd_sc_hd__or2_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09947_ _10110_/CLK _09947_/D repeater405/X VGND VGND VPWR VPWR _09947_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09878_ _10409_/CLK _09878_/D repeater406/X VGND VGND VPWR VPWR _09878_/Q sky130_fd_sc_hd__dfstp_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08829_/A _08847_/B VGND VGND VPWR VPWR _09065_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10018_ _10490_/CLK _10018_/D repeater404/X VGND VGND VPWR VPWR _10018_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05490_ _08354_/A _05490_/B VGND VGND VPWR VPWR _05491_/A sky130_fd_sc_hd__and2_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07160_ _06763_/A _07159_/X _09761_/Q _06764_/X VGND VGND VPWR VPWR _09761_/D sky130_fd_sc_hd__o22a_1
X_07091_ _10491_/Q VGND VGND VPWR VPWR _09505_/A sky130_fd_sc_hd__inv_6
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06111_ _06111_/A VGND VGND VPWR VPWR _06111_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06042_ _10078_/Q _06038_/X _06683_/B1 _06039_/Y VGND VGND VPWR VPWR _10078_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09801_ net399_2/A _09801_/D _06622_/X VGND VGND VPWR VPWR _09801_/Q sky130_fd_sc_hd__dfrtp_2
X_09732_ _09732_/A _09517_/A VGND VGND VPWR VPWR _09732_/Z sky130_fd_sc_hd__ebufn_1
X_07993_ _08026_/A _10002_/Q _08010_/C _08019_/C VGND VGND VPWR VPWR _08219_/A sky130_fd_sc_hd__or4_4
X_06944_ _09987_/Q VGND VGND VPWR VPWR _06944_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06875_ _10362_/Q VGND VGND VPWR VPWR _06875_/Y sky130_fd_sc_hd__inv_2
X_09663_ _09662_/X _10396_/Q _10299_/Q VGND VGND VPWR VPWR _09663_/X sky130_fd_sc_hd__mux2_2
X_08614_ _09085_/C _08624_/A VGND VGND VPWR VPWR _08768_/C sky130_fd_sc_hd__or2_2
X_05826_ _10208_/Q _05822_/X _09576_/X _05823_/Y VGND VGND VPWR VPWR _10208_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09594_ _08135_/Y _10332_/Q _09700_/S VGND VGND VPWR VPWR _09594_/X sky130_fd_sc_hd__mux2_1
X_08545_ _08545_/A _08951_/A VGND VGND VPWR VPWR _08546_/B sky130_fd_sc_hd__or2_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05757_ _10248_/Q _05750_/X _09550_/A0 _05752_/X VGND VGND VPWR VPWR _10248_/D sky130_fd_sc_hd__a22o_1
X_05688_ _10289_/Q _05679_/A _09574_/X _05680_/A VGND VGND VPWR VPWR _10289_/D sky130_fd_sc_hd__a22o_1
X_08476_ _08476_/A _08476_/B _09247_/B VGND VGND VPWR VPWR _08567_/A sky130_fd_sc_hd__or3b_1
X_07427_ _07427_/A VGND VGND VPWR VPWR _07428_/A sky130_fd_sc_hd__inv_2
XFILLER_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07358_ _10181_/Q VGND VGND VPWR VPWR _07358_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06309_ _09957_/Q _06305_/X _09576_/X _06306_/Y VGND VGND VPWR VPWR _09957_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ _07289_/A _07289_/B _07288_/X VGND VGND VPWR VPWR _07290_/A sky130_fd_sc_hd__or3b_4
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09028_ _09171_/A _09357_/B VGND VGND VPWR VPWR _09311_/C sky130_fd_sc_hd__or2_1
XFILLER_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _09485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _05318_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_155 _06714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 input36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10498_ _10500_/CLK _10498_/D repeater407/X VGND VGND VPWR VPWR _10498_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04990_ _10451_/Q _04981_/A _09536_/A3 _04982_/A VGND VGND VPWR VPWR _10451_/D sky130_fd_sc_hd__a22o_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06660_ _06660_/A VGND VGND VPWR VPWR _06660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05611_ _10332_/Q _05604_/X _09658_/A1 _05606_/X VGND VGND VPWR VPWR _10332_/D sky130_fd_sc_hd__a22o_1
X_06591_ _06591_/A VGND VGND VPWR VPWR _06592_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05542_ _05543_/A VGND VGND VPWR VPWR _05542_/X sky130_fd_sc_hd__clkbuf_2
X_08330_ _09799_/Q VGND VGND VPWR VPWR _08330_/Y sky130_fd_sc_hd__clkinv_2
X_05473_ _05473_/A VGND VGND VPWR VPWR _05474_/B sky130_fd_sc_hd__clkbuf_2
X_08261_ _07332_/Y _08184_/X _07362_/Y _08158_/X VGND VGND VPWR VPWR _08261_/X sky130_fd_sc_hd__o22a_1
X_07212_ _10182_/Q VGND VGND VPWR VPWR _07212_/Y sky130_fd_sc_hd__inv_2
X_08192_ _06786_/Y _08183_/X _08185_/X _08191_/X VGND VGND VPWR VPWR _08218_/C sky130_fd_sc_hd__o211a_1
XFILLER_106_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07143_ _07138_/Y _06329_/B _09473_/A _06359_/A _07142_/X VGND VGND VPWR VPWR _07156_/B
+ sky130_fd_sc_hd__o221a_1
X_07074_ _10157_/Q VGND VGND VPWR VPWR _07074_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput310 _10455_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_2
XFILLER_145_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06025_ _06026_/A VGND VGND VPWR VPWR _06025_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput332 _10452_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_2
Xoutput321 _10465_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_2
Xoutput343 _09556_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_2
Xoutput376 _09734_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput365 _09748_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_126_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput387 _09763_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput354 _10477_/Q VGND VGND VPWR VPWR sram_ro_addr[5] sky130_fd_sc_hd__buf_2
X_07976_ _06993_/Y _07645_/A _07974_/Y _07523_/A _07975_/X VGND VGND VPWR VPWR _07977_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06927_ _10119_/Q VGND VGND VPWR VPWR _06927_/Y sky130_fd_sc_hd__inv_4
X_09715_ _10501_/Q _09483_/A VGND VGND VPWR VPWR _09715_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09646_ _08334_/X _09800_/Q _09773_/Q VGND VGND VPWR VPWR _09646_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06858_ _10375_/Q VGND VGND VPWR VPWR _06858_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09577_ hold50/X _10381_/Q _10299_/Q VGND VGND VPWR VPWR _09577_/X sky130_fd_sc_hd__mux2_8
X_05809_ _05810_/A VGND VGND VPWR VPWR _05809_/X sky130_fd_sc_hd__clkbuf_2
X_06789_ _06789_/A _06789_/B _06788_/X VGND VGND VPWR VPWR _06834_/B sky130_fd_sc_hd__or3b_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08528_ _08582_/A _08528_/B VGND VGND VPWR VPWR _08529_/A sky130_fd_sc_hd__or2_1
XFILLER_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _08927_/A VGND VGND VPWR VPWR _08951_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_168_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10421_ _10406_/CLK _10421_/D _05370_/X VGND VGND VPWR VPWR _10421_/Q sky130_fd_sc_hd__dfrtn_1
X_10352_ _10354_/CLK _10352_/D repeater406/X VGND VGND VPWR VPWR _10352_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10283_ _10283_/CLK _10283_/D repeater406/X VGND VGND VPWR VPWR _10283_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10135_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07830_ _06827_/Y _07828_/X _06792_/Y _07829_/X VGND VGND VPWR VPWR _07830_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07761_ _07761_/A _07761_/B _07761_/C _07761_/D VGND VGND VPWR VPWR _07776_/B sky130_fd_sc_hd__and4_1
X_09500_ _09500_/A VGND VGND VPWR VPWR _09500_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04973_ _10462_/Q _04966_/X _09658_/A1 _04968_/X VGND VGND VPWR VPWR _10462_/D sky130_fd_sc_hd__a22o_1
X_06712_ _09840_/Q VGND VGND VPWR VPWR _06712_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07692_ _07220_/Y _07667_/X _07183_/Y _07668_/X VGND VGND VPWR VPWR _07692_/X sky130_fd_sc_hd__o22a_1
X_09431_ _09431_/A _09431_/B _09431_/C VGND VGND VPWR VPWR _09443_/C sky130_fd_sc_hd__or3_4
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06643_ _09791_/Q _04903_/A _06684_/B1 _04904_/A VGND VGND VPWR VPWR _09791_/D sky130_fd_sc_hd__a22o_1
X_09362_ _09384_/C _09362_/B _09362_/C VGND VGND VPWR VPWR _09434_/B sky130_fd_sc_hd__or3_1
X_06574_ _06574_/A VGND VGND VPWR VPWR _06574_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05525_ _09684_/X _10378_/Q _05525_/S VGND VGND VPWR VPWR _05526_/A sky130_fd_sc_hd__mux2_1
X_08313_ _06990_/Y _08179_/A _07024_/Y _08180_/A VGND VGND VPWR VPWR _08313_/X sky130_fd_sc_hd__o22a_1
X_09293_ _08688_/A _08977_/C _08978_/B VGND VGND VPWR VPWR _09294_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_11 _05248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _07055_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _09565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_55 _05179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _07861_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05456_ _05459_/A VGND VGND VPWR VPWR _05457_/A sky130_fd_sc_hd__clkbuf_1
X_08244_ _05315_/Y _08188_/X _05267_/Y _08189_/X VGND VGND VPWR VPWR _08244_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 _07288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ _06821_/Y _08173_/X _06808_/Y _08174_/X VGND VGND VPWR VPWR _08175_/X sky130_fd_sc_hd__o22a_1
XANTENNA_99 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05387_ _05387_/A VGND VGND VPWR VPWR _05387_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07126_ _09818_/Q VGND VGND VPWR VPWR _07126_/Y sky130_fd_sc_hd__inv_2
X_07057_ _07052_/Y _05625_/C _09519_/A _05980_/B _07056_/X VGND VGND VPWR VPWR _07057_/X
+ sky130_fd_sc_hd__o221a_1
X_06008_ _10098_/Q _06003_/X _06684_/B1 _06004_/Y VGND VGND VPWR VPWR _10098_/D sky130_fd_sc_hd__a22o_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07959_ _07093_/Y _07828_/A _07110_/Y _07829_/A VGND VGND VPWR VPWR _07959_/X sky130_fd_sc_hd__o22a_1
XFILLER_75_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09629_ _09628_/X _09888_/Q _09776_/Q VGND VGND VPWR VPWR _09629_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10404_ _10404_/CLK _10404_/D hold41/X VGND VGND VPWR VPWR _10404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10335_ _10336_/CLK _10335_/D repeater409/X VGND VGND VPWR VPWR _10335_/Q sky130_fd_sc_hd__dfrtp_4
X_10266_ _10268_/CLK _10266_/D repeater404/X VGND VGND VPWR VPWR _10266_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10197_ _10244_/CLK _10197_/D repeater403/X VGND VGND VPWR VPWR _10197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06290_ _06290_/A VGND VGND VPWR VPWR _06291_/B sky130_fd_sc_hd__buf_6
X_05310_ _10063_/Q VGND VGND VPWR VPWR _05310_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05241_ _10012_/Q VGND VGND VPWR VPWR _05241_/Y sky130_fd_sc_hd__clkinv_2
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_2
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_6
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_6
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_6
X_05172_ _10081_/Q VGND VGND VPWR VPWR _05172_/Y sky130_fd_sc_hd__inv_2
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_6
XFILLER_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput75 hold42/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__buf_12
Xinput97 sram_ro_data[13] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_2
X_09980_ _10350_/CLK _09980_/D repeater405/X VGND VGND VPWR VPWR _09980_/Q sky130_fd_sc_hd__dfrtp_1
X_08931_ _08931_/A VGND VGND VPWR VPWR _09065_/B sky130_fd_sc_hd__inv_2
X_08862_ _08862_/A _09084_/B VGND VGND VPWR VPWR _08863_/A sky130_fd_sc_hd__or2_1
X_07813_ _07813_/A VGND VGND VPWR VPWR _07813_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08793_ _08897_/B VGND VGND VPWR VPWR _09337_/A sky130_fd_sc_hd__clkinv_2
X_07744_ _07744_/A _07744_/B _07744_/C VGND VGND VPWR VPWR _07744_/Y sky130_fd_sc_hd__nand3_2
X_04956_ _09674_/X _09676_/X _09670_/X _09668_/X VGND VGND VPWR VPWR _05103_/B sky130_fd_sc_hd__or4_1
X_07675_ _07200_/Y _07618_/X _07245_/Y _07619_/X _07674_/X VGND VGND VPWR VPWR _07695_/A
+ sky130_fd_sc_hd__o221a_2
X_04887_ _04888_/A VGND VGND VPWR VPWR _04887_/X sky130_fd_sc_hd__clkbuf_2
X_09414_ _09444_/A _09447_/C VGND VGND VPWR VPWR _09414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06626_ _09800_/Q _06605_/A _09645_/X _06606_/A VGND VGND VPWR VPWR _09800_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06557_ _09816_/Q _06552_/X hold46/X _06553_/Y VGND VGND VPWR VPWR _09816_/D sky130_fd_sc_hd__a22o_1
X_09345_ _09345_/A _09421_/C _09400_/C _09399_/C VGND VGND VPWR VPWR _09345_/Y sky130_fd_sc_hd__nor4_1
X_05508_ _09688_/X _10382_/Q _05512_/S VGND VGND VPWR VPWR _05509_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09276_ _09276_/A _09352_/B VGND VGND VPWR VPWR _09432_/B sky130_fd_sc_hd__nor2_1
X_06488_ _09858_/Q _06482_/X _09547_/A1 _06484_/X VGND VGND VPWR VPWR _09858_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08227_ _06712_/Y _08186_/X _06728_/Y _08187_/X _08226_/X VGND VGND VPWR VPWR _08227_/X
+ sky130_fd_sc_hd__o221a_1
X_05439_ _10404_/Q _05435_/X _09580_/X _05437_/X VGND VGND VPWR VPWR _10404_/D sky130_fd_sc_hd__a22o_1
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08158_ _08158_/A VGND VGND VPWR VPWR _08158_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08089_ _08208_/A VGND VGND VPWR VPWR _08089_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07109_ _09997_/Q VGND VGND VPWR VPWR _09483_/A sky130_fd_sc_hd__clkinv_8
X_10120_ _10289_/CLK _10120_/D repeater402/X VGND VGND VPWR VPWR _10120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10051_ _10513_/CLK _10051_/D repeater405/X VGND VGND VPWR VPWR _10051_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10405_/CLK _10318_/D hold41/X VGND VGND VPWR VPWR _10318_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _10504_/CLK _10249_/D repeater403/X VGND VGND VPWR VPWR _10249_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04810_ _10273_/Q input127/X _10509_/Q VGND VGND VPWR VPWR _09714_/A sky130_fd_sc_hd__mux2_1
X_05790_ _10229_/Q _05786_/X _09576_/X _05787_/Y VGND VGND VPWR VPWR _10229_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07460_ _07421_/X _07452_/A _09735_/Q _07453_/A VGND VGND VPWR VPWR _09735_/D sky130_fd_sc_hd__o22a_1
X_07391_ _07389_/Y _05727_/A _07390_/Y _06351_/B VGND VGND VPWR VPWR _07391_/X sky130_fd_sc_hd__o22a_2
X_06411_ _09896_/Q _06404_/A _09660_/A1 _06405_/A VGND VGND VPWR VPWR _09896_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06342_ _06342_/A VGND VGND VPWR VPWR _06342_/X sky130_fd_sc_hd__clkbuf_2
X_09130_ _09265_/A _09099_/X _09127_/X _09129_/Y VGND VGND VPWR VPWR _09130_/X sky130_fd_sc_hd__o211a_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09061_ _09395_/B _09207_/B VGND VGND VPWR VPWR _09389_/A sky130_fd_sc_hd__or2_1
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06273_ _09979_/Q _06268_/X _09579_/X _06270_/X VGND VGND VPWR VPWR _09979_/D sky130_fd_sc_hd__a22o_1
X_08012_ _05343_/Y _08179_/A _05304_/Y _08180_/A VGND VGND VPWR VPWR _08012_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05224_ _05212_/Y _06515_/A _07606_/A _06266_/A _05223_/X VGND VGND VPWR VPWR _05236_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05155_ _05155_/A _05155_/B VGND VGND VPWR VPWR _05615_/B sky130_fd_sc_hd__or2_1
X_09963_ _10244_/CLK _09963_/D repeater403/X VGND VGND VPWR VPWR _09963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05086_ _10045_/Q _05084_/Y _10459_/Q _06689_/A VGND VGND VPWR VPWR _05086_/X sky130_fd_sc_hd__a22o_1
X_08914_ _08977_/C _09015_/B VGND VGND VPWR VPWR _08914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09894_ _10495_/CLK _09894_/D repeater404/X VGND VGND VPWR VPWR _09894_/Q sky130_fd_sc_hd__dfstp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08845_ _08845_/A _08853_/B VGND VGND VPWR VPWR _09386_/A sky130_fd_sc_hd__nor2_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _08776_/A _08776_/B VGND VGND VPWR VPWR _08776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07727_ _10137_/Q VGND VGND VPWR VPWR _07727_/Y sky130_fd_sc_hd__inv_2
X_05988_ _10110_/Q _05981_/X _09658_/A1 _05983_/X VGND VGND VPWR VPWR _10110_/D sky130_fd_sc_hd__a22o_1
X_04939_ _10478_/Q _04935_/X _09580_/X _04937_/X VGND VGND VPWR VPWR _10478_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07658_ _07818_/A VGND VGND VPWR VPWR _07658_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07589_ _07589_/A VGND VGND VPWR VPWR _07801_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06609_ _06609_/A VGND VGND VPWR VPWR _06609_/X sky130_fd_sc_hd__clkbuf_1
X_09328_ _09447_/A _09328_/B _09380_/D _09411_/C VGND VGND VPWR VPWR _09331_/A sky130_fd_sc_hd__or4_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09259_ _08678_/X _09261_/A _08674_/X _09261_/A _09258_/X VGND VGND VPWR VPWR _09264_/A
+ sky130_fd_sc_hd__o221ai_2
XFILLER_181_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10103_ _10283_/CLK _10103_/D repeater406/X VGND VGND VPWR VPWR _10103_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10034_ _10135_/CLK _10034_/D _07492_/B VGND VGND VPWR VPWR _10034_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06960_ _06960_/A _06960_/B _06960_/C _06960_/D VGND VGND VPWR VPWR _07028_/A sky130_fd_sc_hd__and4_1
XFILLER_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05911_ _05912_/A VGND VGND VPWR VPWR _05911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06891_ _10042_/Q VGND VGND VPWR VPWR _06891_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05842_ _05842_/A VGND VGND VPWR VPWR _05842_/X sky130_fd_sc_hd__clkbuf_2
X_08630_ _08883_/A VGND VGND VPWR VPWR _08761_/A sky130_fd_sc_hd__buf_2
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08561_ _08634_/B _08561_/B _08571_/C _08888_/A VGND VGND VPWR VPWR _08911_/B sky130_fd_sc_hd__or4_2
X_05773_ _10237_/Q _05764_/A _09659_/A1 _05765_/A VGND VGND VPWR VPWR _10237_/D sky130_fd_sc_hd__a22o_1
X_08492_ _08492_/A _08492_/B _08492_/C VGND VGND VPWR VPWR _08546_/A sky130_fd_sc_hd__or3_4
X_07512_ _07512_/A VGND VGND VPWR VPWR _07568_/B sky130_fd_sc_hd__buf_4
X_07443_ _06835_/X _07439_/X _09748_/Q _07441_/X VGND VGND VPWR VPWR _09748_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07374_ _07374_/A _07374_/B _07374_/C _07374_/D VGND VGND VPWR VPWR _07419_/B sky130_fd_sc_hd__and4_1
X_09113_ _09113_/A VGND VGND VPWR VPWR _09113_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06325_ _09778_/Q _06176_/A _06133_/Y _06262_/B _09946_/Q VGND VGND VPWR VPWR _06325_/X
+ sky130_fd_sc_hd__o221a_1
X_06256_ _09985_/Q _06252_/X _09576_/X _06253_/Y VGND VGND VPWR VPWR _09985_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09044_ _09363_/A _09044_/B VGND VGND VPWR VPWR _09417_/A sky130_fd_sc_hd__or2_2
XFILLER_163_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05207_ _05333_/A _05275_/B VGND VGND VPWR VPWR _06429_/A sky130_fd_sc_hd__or2_1
XFILLER_150_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06187_ _08034_/A _08027_/A _08038_/C VGND VGND VPWR VPWR _08016_/A sky130_fd_sc_hd__or3_1
XFILLER_171_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05138_ _05138_/A VGND VGND VPWR VPWR _05968_/B sky130_fd_sc_hd__buf_6
XFILLER_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09946_ _10006_/CLK _09946_/D _05034_/A VGND VGND VPWR VPWR _09946_/Q sky130_fd_sc_hd__dfrtp_1
X_05069_ _05160_/A _05245_/A VGND VGND VPWR VPWR _06002_/B sky130_fd_sc_hd__or2_2
X_09877_ _10409_/CLK _09877_/D repeater407/X VGND VGND VPWR VPWR _09877_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08828_ _08829_/A _08853_/B VGND VGND VPWR VPWR _09354_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ _09223_/A _08761_/A _08758_/Y VGND VGND VPWR VPWR _08763_/A sky130_fd_sc_hd__o21bai_1
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10017_ _10490_/CLK _10017_/D repeater404/X VGND VGND VPWR VPWR _10017_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07090_ _10092_/Q VGND VGND VPWR VPWR _09491_/A sky130_fd_sc_hd__clkinv_4
X_06110_ _06110_/A VGND VGND VPWR VPWR _06111_/A sky130_fd_sc_hd__inv_2
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06041_ _10079_/Q _06038_/X _09577_/X _06039_/Y VGND VGND VPWR VPWR _10079_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09800_ _09572_/A1 _09800_/D _06625_/X VGND VGND VPWR VPWR _09800_/Q sky130_fd_sc_hd__dfrtp_2
X_07992_ _08040_/C VGND VGND VPWR VPWR _08019_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09731_ _09731_/A _09515_/A VGND VGND VPWR VPWR _09731_/Z sky130_fd_sc_hd__ebufn_1
X_06943_ _10241_/Q VGND VGND VPWR VPWR _06943_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06874_ _10348_/Q VGND VGND VPWR VPWR _06874_/Y sky130_fd_sc_hd__clkinv_2
X_09662_ _09804_/Q _09803_/Q _09773_/Q VGND VGND VPWR VPWR _09662_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08613_ _08766_/A _08883_/B _09790_/Q VGND VGND VPWR VPWR _09222_/B sky130_fd_sc_hd__o21ai_1
X_05825_ _10209_/Q _05822_/X _09577_/X _05823_/Y VGND VGND VPWR VPWR _10209_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09593_ _09592_/X _09908_/Q _09776_/Q VGND VGND VPWR VPWR _09593_/X sky130_fd_sc_hd__mux2_1
X_05756_ _10249_/Q _05750_/X _09547_/A1 _05752_/X VGND VGND VPWR VPWR _10249_/D sky130_fd_sc_hd__a22o_1
X_08544_ _08923_/A VGND VGND VPWR VPWR _08925_/A sky130_fd_sc_hd__buf_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05687_ _10290_/Q _05679_/A hold46/X _05680_/A VGND VGND VPWR VPWR _10290_/D sky130_fd_sc_hd__a22o_1
XFILLER_168_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08475_ _09137_/A VGND VGND VPWR VPWR _09415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07426_ _07427_/A VGND VGND VPWR VPWR _07426_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07357_ _09842_/Q VGND VGND VPWR VPWR _07357_/Y sky130_fd_sc_hd__clkinv_2
X_06308_ _09958_/Q _06305_/X _09577_/X _06306_/Y VGND VGND VPWR VPWR _09958_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07288_ _07288_/A _07288_/B _07288_/C _07288_/D VGND VGND VPWR VPWR _07288_/X sky130_fd_sc_hd__and4_2
X_09027_ _08527_/Y _09002_/Y _09022_/X _09201_/C _09369_/A VGND VGND VPWR VPWR _09032_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_163_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06239_ _09991_/Q _07551_/B _07592_/A VGND VGND VPWR VPWR _07584_/B sky130_fd_sc_hd__or3_2
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09929_ _10119_/CLK _09929_/D repeater403/X VGND VGND VPWR VPWR _09929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _09485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _05327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_156 _06714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_178 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10497_ _10500_/CLK _10497_/D repeater407/X VGND VGND VPWR VPWR _10497_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_2
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05610_ _10333_/Q _05604_/X _09545_/A1 _05606_/X VGND VGND VPWR VPWR _10333_/D sky130_fd_sc_hd__a22o_1
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06590_ _09809_/Q _06589_/X _07489_/A _06593_/B VGND VGND VPWR VPWR _09809_/D sky130_fd_sc_hd__o22a_1
X_05541_ _05541_/A _05541_/B VGND VGND VPWR VPWR _05543_/A sky130_fd_sc_hd__or2_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05472_ _09692_/X _05450_/A _10391_/Q _05493_/D VGND VGND VPWR VPWR _10391_/D sky130_fd_sc_hd__a22o_1
X_08260_ _07388_/Y _08177_/X _07401_/Y _08178_/X _08259_/X VGND VGND VPWR VPWR _08274_/B
+ sky130_fd_sc_hd__o221a_1
X_07211_ _07206_/Y _05952_/B _07207_/Y _06360_/B _07210_/X VGND VGND VPWR VPWR _07218_/C
+ sky130_fd_sc_hd__o221a_1
X_08191_ _06785_/Y _08186_/X _06815_/Y _08187_/X _08190_/X VGND VGND VPWR VPWR _08191_/X
+ sky130_fd_sc_hd__o221a_1
X_07142_ _09459_/A _05433_/A _07141_/Y _06494_/B VGND VGND VPWR VPWR _07142_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07073_ _10183_/Q VGND VGND VPWR VPWR _07073_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput300 _10434_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput344 _09524_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_2
Xoutput311 _10456_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_2
Xoutput322 _10466_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_2
Xoutput333 _09766_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_2
X_06024_ _06108_/A _06024_/B VGND VGND VPWR VPWR _06026_/A sky130_fd_sc_hd__or2_2
XFILLER_160_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput377 _09735_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput366 _09749_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_126_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput355 _10478_/Q VGND VGND VPWR VPWR sram_ro_addr[6] sky130_fd_sc_hd__buf_2
Xoutput388 _09764_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_2
X_07975_ _07015_/Y _07646_/A _06957_/Y _07807_/A VGND VGND VPWR VPWR _07975_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09714_ _09714_/A _09481_/A VGND VGND VPWR VPWR _09714_/Z sky130_fd_sc_hd__ebufn_1
X_06926_ _10179_/Q VGND VGND VPWR VPWR _06926_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06857_ _10146_/Q VGND VGND VPWR VPWR _06857_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09645_ _08332_/X _09799_/Q _09773_/Q VGND VGND VPWR VPWR _09645_/X sky130_fd_sc_hd__mux2_1
X_05808_ _05896_/A _05808_/B VGND VGND VPWR VPWR _05810_/A sky130_fd_sc_hd__or2_2
XFILLER_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09576_ hold44/X _10380_/Q _10299_/Q VGND VGND VPWR VPWR _09576_/X sky130_fd_sc_hd__mux2_8
X_06788_ _06783_/Y _06538_/B _06784_/Y _06096_/B _06787_/X VGND VGND VPWR VPWR _06788_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_42_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05739_ _10258_/Q _05730_/A _09574_/X _05731_/A VGND VGND VPWR VPWR _10258_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_08527_ _08957_/A VGND VGND VPWR VPWR _08527_/Y sky130_fd_sc_hd__inv_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _09085_/D _09085_/B _08493_/B VGND VGND VPWR VPWR _08927_/A sky130_fd_sc_hd__or3_4
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07409_ _10233_/Q VGND VGND VPWR VPWR _07409_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08389_ _08389_/A VGND VGND VPWR VPWR _08493_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10420_ _09572_/A1 _10420_/D _05379_/X VGND VGND VPWR VPWR _10420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10351_ _10354_/CLK _10351_/D repeater406/X VGND VGND VPWR VPWR _10351_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10282_ _10405_/CLK _10282_/D hold41/X VGND VGND VPWR VPWR _10282_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07760_ _06864_/Y _07645_/X _06874_/Y _07758_/X _07759_/X VGND VGND VPWR VPWR _07761_/D
+ sky130_fd_sc_hd__o221a_1
X_04972_ _10463_/Q _04966_/X _09545_/A1 _04968_/X VGND VGND VPWR VPWR _10463_/D sky130_fd_sc_hd__a22o_1
X_06711_ _09940_/Q VGND VGND VPWR VPWR _06711_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09430_ _09053_/X _09429_/X _08918_/B _09016_/D VGND VGND VPWR VPWR _09431_/B sky130_fd_sc_hd__o211ai_1
X_07691_ _07225_/Y _06232_/X _07202_/Y _07533_/A _07690_/X VGND VGND VPWR VPWR _07694_/C
+ sky130_fd_sc_hd__o221a_1
X_06642_ _09792_/Q _06636_/X _09574_/X _06637_/Y VGND VGND VPWR VPWR _09792_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09361_ _09434_/A _09393_/B _09432_/B VGND VGND VPWR VPWR _09361_/Y sky130_fd_sc_hd__nor3_1
X_06573_ _06591_/A VGND VGND VPWR VPWR _06574_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05524_ _05524_/A VGND VGND VPWR VPWR _05524_/X sky130_fd_sc_hd__clkbuf_1
X_08312_ _06939_/Y _08219_/A _07012_/Y _08220_/A _08311_/X VGND VGND VPWR VPWR _08328_/A
+ sky130_fd_sc_hd__o221a_1
X_09292_ _09292_/A _09387_/C _09357_/D _09428_/A VGND VGND VPWR VPWR _09298_/A sky130_fd_sc_hd__or4_4
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_23 _07071_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 _05265_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ _05317_/Y _08184_/X _05218_/Y _08158_/X VGND VGND VPWR VPWR _08243_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_45 _07869_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05455_ _09697_/X _05449_/X _10396_/Q _05451_/X VGND VGND VPWR VPWR _10396_/D sky130_fd_sc_hd__a22o_1
XANTENNA_56 _09521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_34 _07323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08174_ _08174_/A VGND VGND VPWR VPWR _08174_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_67 _09538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05386_ _05406_/A VGND VGND VPWR VPWR _05387_/A sky130_fd_sc_hd__clkbuf_1
X_07125_ _09977_/Q VGND VGND VPWR VPWR _09481_/A sky130_fd_sc_hd__clkinv_8
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07056_ _07054_/Y _06045_/B _07055_/Y _06002_/B VGND VGND VPWR VPWR _07056_/X sky130_fd_sc_hd__o22a_1
X_06007_ _10099_/Q _06003_/X _06683_/B1 _06004_/Y VGND VGND VPWR VPWR _10099_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ _07097_/Y _06232_/A _07152_/Y _07519_/A _07957_/X VGND VGND VPWR VPWR _07961_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07889_ _07333_/Y _07779_/X _07887_/Y _07781_/X _07888_/X VGND VGND VPWR VPWR _07889_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06909_ _10075_/Q VGND VGND VPWR VPWR _06909_/Y sky130_fd_sc_hd__inv_2
X_09628_ _07886_/Y _10324_/Q _09682_/S VGND VGND VPWR VPWR _09628_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09559_ _10275_/Q input3/X input1/X VGND VGND VPWR VPWR _09559_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10403_ _10405_/CLK _10403_/D hold41/X VGND VGND VPWR VPWR _10403_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10334_ _10336_/CLK _10334_/D repeater409/X VGND VGND VPWR VPWR _10334_/Q sky130_fd_sc_hd__dfrtp_4
X_10265_ _10290_/CLK _10265_/D repeater402/X VGND VGND VPWR VPWR _10265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ _10289_/CLK _10196_/D repeater402/X VGND VGND VPWR VPWR _10196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05240_ _05305_/B _05357_/B VGND VGND VPWR VPWR _05575_/A sky130_fd_sc_hd__or2_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_6
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_4
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
X_05171_ _10324_/Q _05156_/Y _05159_/X _05170_/X VGND VGND VPWR VPWR _05183_/C sky130_fd_sc_hd__a211o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__buf_12
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_6
Xinput76 qspi_enabled VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_6
Xinput98 sram_ro_data[14] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08930_ _08938_/A _08935_/B VGND VGND VPWR VPWR _08931_/A sky130_fd_sc_hd__or2_2
X_08861_ _08861_/A _09427_/A VGND VGND VPWR VPWR _08866_/A sky130_fd_sc_hd__or2_1
XFILLER_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07812_ _07812_/A VGND VGND VPWR VPWR _07812_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08792_ _08849_/A VGND VGND VPWR VPWR _08897_/B sky130_fd_sc_hd__clkbuf_4
X_07743_ _07743_/A _07743_/B _07743_/C _07743_/D VGND VGND VPWR VPWR _07744_/C sky130_fd_sc_hd__and4_1
X_04955_ _04955_/A VGND VGND VPWR VPWR _10469_/D sky130_fd_sc_hd__clkbuf_1
X_04886_ _04993_/A _04886_/B VGND VGND VPWR VPWR _04888_/A sky130_fd_sc_hd__or2_2
X_07674_ _07219_/Y _07620_/X _07177_/Y _07621_/X _07673_/X VGND VGND VPWR VPWR _07674_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09413_ _08753_/C _09412_/Y _08700_/C _09235_/C _09325_/B VGND VGND VPWR VPWR _09447_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06625_ _06625_/A VGND VGND VPWR VPWR _06625_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06556_ _09817_/Q _06552_/X _09576_/X _06553_/Y VGND VGND VPWR VPWR _09817_/D sky130_fd_sc_hd__a22o_1
X_09344_ _09344_/A _09344_/B VGND VGND VPWR VPWR _09399_/C sky130_fd_sc_hd__nor2_1
XFILLER_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05507_ _05507_/A VGND VGND VPWR VPWR _05507_/X sky130_fd_sc_hd__clkbuf_1
X_09275_ _09275_/A _09348_/B _09348_/C _09274_/X VGND VGND VPWR VPWR _09275_/X sky130_fd_sc_hd__or4b_1
X_06487_ _09859_/Q _06482_/X _09579_/X _06484_/X VGND VGND VPWR VPWR _09859_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08226_ _06754_/Y _08188_/X _06752_/Y _08189_/X VGND VGND VPWR VPWR _08226_/X sky130_fd_sc_hd__o22a_1
X_05438_ _10405_/Q _05435_/X _09581_/X _05437_/X VGND VGND VPWR VPWR _10405_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08157_ _06888_/Y _08058_/X _06877_/Y _08059_/X _08156_/X VGND VGND VPWR VPWR _08172_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_146_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07108_ _10015_/Q VGND VGND VPWR VPWR _09485_/A sky130_fd_sc_hd__inv_4
X_05369_ _05378_/A VGND VGND VPWR VPWR _05370_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08088_ _08207_/A VGND VGND VPWR VPWR _08088_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _10374_/CLK sky130_fd_sc_hd__clkbuf_16
X_07039_ _10058_/Q _05162_/X input38/X _09699_/S _07038_/X VGND VGND VPWR VPWR _07040_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10050_ _10513_/CLK _10050_/D repeater405/X VGND VGND VPWR VPWR _10050_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10317_ _10405_/CLK _10317_/D hold41/X VGND VGND VPWR VPWR _10317_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10296_/CLK _10248_/D repeater402/X VGND VGND VPWR VPWR _10248_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10179_ _10254_/CLK _10179_/D repeater407/X VGND VGND VPWR VPWR _10179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06410_ _09897_/Q _06403_/X _09550_/A0 _06405_/X VGND VGND VPWR VPWR _09897_/D sky130_fd_sc_hd__a22o_1
X_07390_ _09929_/Q VGND VGND VPWR VPWR _07390_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06341_ _06341_/A VGND VGND VPWR VPWR _06342_/A sky130_fd_sc_hd__inv_2
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09060_ _09060_/A _09307_/B VGND VGND VPWR VPWR _09283_/C sky130_fd_sc_hd__or2_1
X_06272_ _09980_/Q _06268_/X _09580_/X _06270_/X VGND VGND VPWR VPWR _09980_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05223_ _05218_/Y _06250_/A _05221_/Y _06205_/A VGND VGND VPWR VPWR _05223_/X sky130_fd_sc_hd__o22a_1
X_08011_ _08037_/B _08032_/A _08019_/C VGND VGND VPWR VPWR _08180_/A sky130_fd_sc_hd__or3_4
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05154_ _10329_/Q _05151_/X input100/X _05153_/X VGND VGND VPWR VPWR _05183_/B sky130_fd_sc_hd__a22o_1
X_09962_ _10244_/CLK _09962_/D repeater403/X VGND VGND VPWR VPWR _09962_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05085_ _05085_/A VGND VGND VPWR VPWR _06689_/A sky130_fd_sc_hd__clkinv_2
X_08913_ _08913_/A _08913_/B _08913_/C VGND VGND VPWR VPWR _08977_/C sky130_fd_sc_hd__or3_4
X_09893_ _10023_/CLK _09893_/D repeater409/X VGND VGND VPWR VPWR _09893_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A _09397_/B VGND VGND VPWR VPWR _08846_/A sky130_fd_sc_hd__or2_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08775_ _08775_/A _09247_/D VGND VGND VPWR VPWR _08776_/B sky130_fd_sc_hd__or2_2
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05987_ _10111_/Q _05981_/X _09545_/A1 _05983_/X VGND VGND VPWR VPWR _10111_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04938_ _10479_/Q _04935_/X _09581_/X _04937_/X VGND VGND VPWR VPWR _10479_/D sky130_fd_sc_hd__a22o_1
X_07726_ _10033_/Q VGND VGND VPWR VPWR _07726_/Y sky130_fd_sc_hd__inv_2
X_04869_ _05313_/A _05327_/A VGND VGND VPWR VPWR _04870_/A sky130_fd_sc_hd__or2_1
X_07657_ _07817_/A VGND VGND VPWR VPWR _07657_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07588_ _10029_/Q VGND VGND VPWR VPWR _07588_/Y sky130_fd_sc_hd__inv_2
X_06608_ _06614_/A VGND VGND VPWR VPWR _06609_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_159_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09327_ _09327_/A _09327_/B _09327_/C _09327_/D VGND VGND VPWR VPWR _09411_/C sky130_fd_sc_hd__or4_1
X_06539_ _06540_/A VGND VGND VPWR VPWR _06539_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09258_ _09101_/Y _09261_/A _09109_/A _09255_/A _09257_/X VGND VGND VPWR VPWR _09258_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08209_ _06797_/Y _08207_/X _06830_/Y _08208_/X VGND VGND VPWR VPWR _08209_/X sky130_fd_sc_hd__o22a_1
X_09189_ _09189_/A _09418_/A VGND VGND VPWR VPWR _09191_/A sky130_fd_sc_hd__or2_1
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10102_ _10283_/CLK _10102_/D repeater406/X VGND VGND VPWR VPWR _10102_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput200 wb_sel_i[2] VGND VGND VPWR VPWR _08353_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10033_ _10135_/CLK _10033_/D _07492_/B VGND VGND VPWR VPWR _10033_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05910_ _05993_/A _05910_/B VGND VGND VPWR VPWR _05912_/A sky130_fd_sc_hd__or2_2
X_06890_ _06885_/Y _06516_/B _06886_/Y _05852_/B _06889_/X VGND VGND VPWR VPWR _06890_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05841_ _05841_/A VGND VGND VPWR VPWR _05842_/A sky130_fd_sc_hd__inv_2
X_05772_ _10238_/Q _05764_/A _09661_/A1 _05765_/A VGND VGND VPWR VPWR _10238_/D sky130_fd_sc_hd__a22o_1
X_08560_ _08583_/A _08927_/B _09149_/A _08559_/X VGND VGND VPWR VPWR _08560_/X sky130_fd_sc_hd__o211a_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08491_ _08491_/A _08491_/B _08491_/C VGND VGND VPWR VPWR _09374_/A sky130_fd_sc_hd__and3_1
X_07511_ _07755_/A VGND VGND VPWR VPWR _07512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07442_ _06759_/X _07439_/X _09749_/Q _07441_/X VGND VGND VPWR VPWR _09749_/D sky130_fd_sc_hd__o22a_1
XFILLER_62_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07373_ _07368_/Y _06472_/B _07369_/Y _06154_/B _07372_/X VGND VGND VPWR VPWR _07374_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09112_ _09377_/B _09283_/A VGND VGND VPWR VPWR _09113_/A sky130_fd_sc_hd__or2_1
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06324_ _09947_/Q _06315_/A _09536_/A3 _06316_/A VGND VGND VPWR VPWR _09947_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06255_ _09986_/Q _06252_/X _09550_/A0 _06253_/Y VGND VGND VPWR VPWR _09986_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09043_ _09043_/A VGND VGND VPWR VPWR _09043_/X sky130_fd_sc_hd__clkbuf_1
X_05206_ _05338_/B VGND VGND VPWR VPWR _05275_/B sky130_fd_sc_hd__buf_2
X_06186_ _08045_/D VGND VGND VPWR VPWR _08038_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05137_ _05355_/A _05311_/B VGND VGND VPWR VPWR _05138_/A sky130_fd_sc_hd__or2_4
XFILLER_145_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09945_ _10257_/CLK _09945_/D repeater407/X VGND VGND VPWR VPWR _09945_/Q sky130_fd_sc_hd__dfrtp_1
X_05068_ _05164_/B VGND VGND VPWR VPWR _05160_/A sky130_fd_sc_hd__clkbuf_1
X_09876_ _10409_/CLK _09876_/D repeater406/X VGND VGND VPWR VPWR _09876_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08827_ _08827_/A VGND VGND VPWR VPWR _09064_/A sky130_fd_sc_hd__inv_2
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08758_ _08758_/A _08898_/A VGND VGND VPWR VPWR _08758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08689_ _08689_/A VGND VGND VPWR VPWR _09278_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _09467_/A _07533_/D _09485_/A _07651_/X _07708_/X VGND VGND VPWR VPWR _07716_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10016_ _10490_/CLK _10016_/D repeater404/X VGND VGND VPWR VPWR _10016_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06040_ _10080_/Q _06038_/X _09578_/X _06039_/Y VGND VGND VPWR VPWR _10080_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _10006_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07991_ _08045_/D VGND VGND VPWR VPWR _08040_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09730_ _10296_/Q _09513_/A VGND VGND VPWR VPWR _09730_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_113_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06942_ _09998_/Q VGND VGND VPWR VPWR _06942_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06873_ _06868_/Y _06313_/B _06869_/Y _06011_/B _06872_/X VGND VGND VPWR VPWR _06880_/C
+ sky130_fd_sc_hd__o221a_1
X_09661_ _10317_/Q _09661_/A1 _09679_/S VGND VGND VPWR VPWR _09661_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05824_ _10210_/Q _05822_/X _09578_/X _05823_/Y VGND VGND VPWR VPWR _10210_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08612_ _08752_/A VGND VGND VPWR VPWR _08766_/A sky130_fd_sc_hd__buf_4
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09592_ _08117_/Y _10331_/Q _09700_/S VGND VGND VPWR VPWR _09592_/X sky130_fd_sc_hd__mux2_1
X_05755_ _10250_/Q _05750_/X _09579_/X _05752_/X VGND VGND VPWR VPWR _10250_/D sky130_fd_sc_hd__a22o_1
X_08543_ _08552_/A _08927_/B VGND VGND VPWR VPWR _08543_/X sky130_fd_sc_hd__or2_1
XFILLER_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05686_ _10291_/Q _05679_/A _09576_/X _05680_/A VGND VGND VPWR VPWR _10291_/D sky130_fd_sc_hd__a22o_1
X_08474_ _08897_/A _08970_/A VGND VGND VPWR VPWR _09137_/A sky130_fd_sc_hd__nor2_1
X_07425_ _07450_/A _07425_/B VGND VGND VPWR VPWR _07427_/A sky130_fd_sc_hd__or2_4
X_07356_ _10220_/Q VGND VGND VPWR VPWR _07356_/Y sky130_fd_sc_hd__clkinv_2
X_06307_ _09959_/Q _06305_/X _09578_/X _06306_/Y VGND VGND VPWR VPWR _09959_/D sky130_fd_sc_hd__a22o_1
X_07287_ _07287_/A _07287_/B _07287_/C _07287_/D VGND VGND VPWR VPWR _07288_/D sky130_fd_sc_hd__and4_1
XFILLER_163_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06238_ _06238_/A VGND VGND VPWR VPWR _07592_/A sky130_fd_sc_hd__clkbuf_2
X_09026_ _09169_/A _09386_/B VGND VGND VPWR VPWR _09369_/A sky130_fd_sc_hd__or2_1
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06169_ _06169_/A VGND VGND VPWR VPWR _06169_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09928_ _10119_/CLK _09928_/D repeater402/X VGND VGND VPWR VPWR _09928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09859_ _10268_/CLK _09859_/D repeater404/X VGND VGND VPWR VPWR _09859_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _05340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _06880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _09487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_179 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10496_ _10500_/CLK _10496_/D repeater407/X VGND VGND VPWR VPWR _10496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05540_ _05540_/A VGND VGND VPWR VPWR _05541_/B sky130_fd_sc_hd__buf_2
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05471_ _05471_/A VGND VGND VPWR VPWR _05471_/X sky130_fd_sc_hd__clkbuf_1
X_07210_ _07208_/Y _04885_/A _07209_/Y _05740_/B VGND VGND VPWR VPWR _07210_/X sky130_fd_sc_hd__o22a_1
X_08190_ _06828_/Y _08188_/X _06805_/Y _08189_/X VGND VGND VPWR VPWR _08190_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07141_ _09852_/Q VGND VGND VPWR VPWR _07141_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07072_ _09897_/Q VGND VGND VPWR VPWR _09471_/A sky130_fd_sc_hd__inv_4
Xoutput301 _10435_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_2
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput312 _10457_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_2
Xoutput323 _10467_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_2
Xoutput334 _09767_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_2
X_06023_ _06337_/A VGND VGND VPWR VPWR _06108_/A sky130_fd_sc_hd__clkbuf_4
Xoutput345 _07500_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_2
Xoutput378 _09736_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_160_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput367 _09750_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput356 _10479_/Q VGND VGND VPWR VPWR sram_ro_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput389 _09765_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07974_ _10341_/Q VGND VGND VPWR VPWR _07974_/Y sky130_fd_sc_hd__clkinv_2
X_09713_ _09713_/A _09479_/A VGND VGND VPWR VPWR _09713_/Z sky130_fd_sc_hd__ebufn_2
X_06925_ _06925_/A _06925_/B _06925_/C _06925_/D VGND VGND VPWR VPWR _06935_/B sky130_fd_sc_hd__or4_2
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06856_ _10493_/Q VGND VGND VPWR VPWR _06856_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09644_ _08330_/Y input58/X _09773_/Q VGND VGND VPWR VPWR _09644_/X sky130_fd_sc_hd__mux2_1
X_05807_ _05807_/A VGND VGND VPWR VPWR _05808_/B sky130_fd_sc_hd__buf_2
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09575_ hold48/X _10379_/Q _10299_/Q VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__mux2_8
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06787_ _06785_/Y _06516_/B _06786_/Y _05434_/B VGND VGND VPWR VPWR _06787_/X sky130_fd_sc_hd__o22a_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05738_ _10259_/Q _05730_/A hold46/X _05731_/A VGND VGND VPWR VPWR _10259_/D sky130_fd_sc_hd__a22o_1
X_08526_ _09006_/A VGND VGND VPWR VPWR _08999_/B sky130_fd_sc_hd__inv_2
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08457_ _08897_/A VGND VGND VPWR VPWR _08457_/X sky130_fd_sc_hd__clkbuf_2
X_05669_ _06568_/A VGND VGND VPWR VPWR _05670_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07408_ _10038_/Q VGND VGND VPWR VPWR _07408_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08388_ _08631_/B VGND VGND VPWR VPWR _08505_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07339_ _10129_/Q VGND VGND VPWR VPWR _07339_/Y sky130_fd_sc_hd__inv_2
X_10350_ _10350_/CLK _10350_/D repeater404/X VGND VGND VPWR VPWR _10350_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09009_ _08491_/A _08999_/A _08491_/B _08546_/Y VGND VGND VPWR VPWR _09205_/A sky130_fd_sc_hd__a31o_1
X_10281_ _10405_/CLK _10281_/D repeater410/X VGND VGND VPWR VPWR _10281_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10479_ _10487_/CLK _10479_/D _05034_/A VGND VGND VPWR VPWR _10479_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04971_ _10464_/Q _04966_/X _09579_/X _04968_/X VGND VGND VPWR VPWR _10464_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06710_ _09861_/Q VGND VGND VPWR VPWR _06710_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07690_ _07690_/A _07770_/B VGND VGND VPWR VPWR _07690_/X sky130_fd_sc_hd__or2_1
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06641_ _09793_/Q _06636_/X hold46/X _06637_/Y VGND VGND VPWR VPWR _09793_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _09278_/B _08909_/Y _09045_/C VGND VGND VPWR VPWR _09393_/B sky130_fd_sc_hd__o21a_1
X_06572_ _06572_/A VGND VGND VPWR VPWR _06591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05523_ _06644_/A VGND VGND VPWR VPWR _05524_/A sky130_fd_sc_hd__clkbuf_1
X_09291_ _09420_/B _09291_/B _09291_/C VGND VGND VPWR VPWR _09428_/A sky130_fd_sc_hd__or3_1
X_08311_ _06969_/Y _08173_/A _06945_/Y _08174_/A VGND VGND VPWR VPWR _08311_/X sky130_fd_sc_hd__o22a_1
X_08242_ _05326_/Y _08177_/X _05276_/Y _08178_/X _08241_/X VGND VGND VPWR VPWR _08256_/B
+ sky130_fd_sc_hd__o221a_2
X_05454_ _05454_/A VGND VGND VPWR VPWR _05454_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_13 _05285_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _07895_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _07957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 input128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _07323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _07500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08173_ _08173_/A VGND VGND VPWR VPWR _08173_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_68 _09554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05385_ _06572_/A VGND VGND VPWR VPWR _05406_/A sky130_fd_sc_hd__buf_6
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07124_ _07119_/Y _06304_/B _09479_/A _06290_/A _07123_/X VGND VGND VPWR VPWR _07124_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07055_ _10100_/Q VGND VGND VPWR VPWR _07055_/Y sky130_fd_sc_hd__clkinv_4
X_06006_ _10100_/Q _06003_/X _09658_/A1 _06004_/Y VGND VGND VPWR VPWR _10100_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07957_ _07957_/A _07983_/B VGND VGND VPWR VPWR _07957_/X sky130_fd_sc_hd__or2_1
XFILLER_101_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06908_ _10328_/Q _05156_/Y input7/X _06838_/X VGND VGND VPWR VPWR _06908_/X sky130_fd_sc_hd__a22o_1
X_07888_ _07397_/Y _07782_/X _07340_/Y _07783_/X VGND VGND VPWR VPWR _07888_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09627_ _09626_/X _09887_/Q _09776_/Q VGND VGND VPWR VPWR _09627_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06839_ input8/X _06838_/X input114/X _05112_/X VGND VGND VPWR VPWR _06839_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09558_ _09893_/Q _10487_/Q _09791_/Q VGND VGND VPWR VPWR _09558_/X sky130_fd_sc_hd__mux2_4
X_08509_ _08631_/B _08631_/C _09102_/C _08890_/A VGND VGND VPWR VPWR _08685_/B sky130_fd_sc_hd__or4_4
X_09489_ _09489_/A VGND VGND VPWR VPWR _09490_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10402_ _10404_/CLK _10402_/D hold41/X VGND VGND VPWR VPWR _10402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10333_ _10510_/CLK _10333_/D repeater409/X VGND VGND VPWR VPWR _10333_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10264_ _10296_/CLK _10264_/D repeater402/X VGND VGND VPWR VPWR _10264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10195_ _10238_/CLK _10195_/D repeater403/X VGND VGND VPWR VPWR _10195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_2
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_8
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_6
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
X_05170_ _10055_/Q _05162_/X input20/X _06704_/A _05169_/X VGND VGND VPWR VPWR _05170_/X
+ sky130_fd_sc_hd__a221o_1
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__buf_12
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__buf_6
XFILLER_128_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__buf_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput99 sram_ro_data[15] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08860_ _08860_/A _09352_/B VGND VGND VPWR VPWR _09427_/A sky130_fd_sc_hd__nor2_1
X_07811_ _07811_/A VGND VGND VPWR VPWR _07811_/X sky130_fd_sc_hd__clkbuf_2
X_08791_ _08836_/A VGND VGND VPWR VPWR _08849_/A sky130_fd_sc_hd__buf_4
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07742_ _06963_/Y _07665_/X _07740_/Y _07666_/X _07741_/X VGND VGND VPWR VPWR _07743_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04954_ _09536_/A3 _10469_/Q _04954_/S VGND VGND VPWR VPWR _04955_/A sky130_fd_sc_hd__mux2_1
X_07673_ _07251_/Y _07622_/X _07256_/Y _07623_/X VGND VGND VPWR VPWR _07673_/X sky130_fd_sc_hd__o22a_1
X_04885_ _04885_/A VGND VGND VPWR VPWR _04886_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09412_ _09223_/B _08761_/A _09046_/B VGND VGND VPWR VPWR _09412_/Y sky130_fd_sc_hd__a21oi_1
X_06624_ _06666_/A VGND VGND VPWR VPWR _06625_/A sky130_fd_sc_hd__clkbuf_1
X_09343_ _09343_/A _09343_/B VGND VGND VPWR VPWR _09400_/C sky130_fd_sc_hd__or2_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06555_ _09818_/Q _06552_/X _09577_/X _06553_/Y VGND VGND VPWR VPWR _09818_/D sky130_fd_sc_hd__a22o_1
X_05506_ _05518_/A VGND VGND VPWR VPWR _05507_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_178_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06486_ _09860_/Q _06482_/X _09580_/X _06484_/X VGND VGND VPWR VPWR _09860_/D sky130_fd_sc_hd__a22o_1
X_09274_ _09274_/A _09425_/D _09425_/B _09348_/D VGND VGND VPWR VPWR _09274_/X sky130_fd_sc_hd__or4_1
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08225_ _06736_/Y _08184_/X _06724_/Y _08158_/X VGND VGND VPWR VPWR _08225_/X sky130_fd_sc_hd__o22a_1
X_05437_ _05437_/A VGND VGND VPWR VPWR _05437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08156_ _06875_/Y _08060_/X _06870_/Y _08061_/X VGND VGND VPWR VPWR _08156_/X sky130_fd_sc_hd__o22a_1
X_05368_ _05042_/A _09680_/S _05367_/X _10422_/Q _05041_/A VGND VGND VPWR VPWR _10422_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07107_ _09513_/A _05851_/A _09457_/A _05549_/A _07106_/X VGND VGND VPWR VPWR _07114_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08087_ _08206_/A VGND VGND VPWR VPWR _08087_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05299_ _06630_/B _05299_/B VGND VGND VPWR VPWR _05820_/A sky130_fd_sc_hd__or2_1
X_07038_ input55/X _05114_/A input64/X _06844_/X VGND VGND VPWR VPWR _07038_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08989_ _09384_/C _09362_/B _08989_/C VGND VGND VPWR VPWR _08990_/B sky130_fd_sc_hd__or3_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10316_ _10405_/CLK _10316_/D hold41/X VGND VGND VPWR VPWR _10316_/Q sky130_fd_sc_hd__dfrtp_1
X_10247_ _10313_/CLK _10247_/D repeater403/X VGND VGND VPWR VPWR _10247_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10178_ _10254_/CLK _10178_/D repeater406/X VGND VGND VPWR VPWR _10178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06340_ _06341_/A VGND VGND VPWR VPWR _06340_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ _09981_/Q _06268_/X _09581_/X _06270_/X VGND VGND VPWR VPWR _09981_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05222_ _05329_/A _05275_/B VGND VGND VPWR VPWR _06205_/A sky130_fd_sc_hd__or2_4
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08010_ _08026_/A _10002_/Q _08010_/C _10006_/Q VGND VGND VPWR VPWR _08179_/A sky130_fd_sc_hd__or4_4
XFILLER_190_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05153_ _05153_/A VGND VGND VPWR VPWR _05153_/X sky130_fd_sc_hd__clkbuf_2
X_09961_ _10244_/CLK _09961_/D repeater403/X VGND VGND VPWR VPWR _09961_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05084_ _06087_/B VGND VGND VPWR VPWR _05084_/Y sky130_fd_sc_hd__inv_2
X_08912_ _08927_/A _08911_/B _08693_/A _08910_/X _08911_/X VGND VGND VPWR VPWR _08912_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09892_ _10397_/CLK _09892_/D repeater409/X VGND VGND VPWR VPWR _09892_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08843_ _08851_/A _08845_/A VGND VGND VPWR VPWR _09397_/B sky130_fd_sc_hd__nor2_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _08774_/A _09229_/B VGND VGND VPWR VPWR _09247_/D sky130_fd_sc_hd__or2_1
X_05986_ _10112_/Q _05981_/X _09579_/X _05983_/X VGND VGND VPWR VPWR _10112_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07725_ _06962_/Y _07632_/X _07022_/Y _07633_/X _07724_/X VGND VGND VPWR VPWR _07732_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04937_ _04937_/A VGND VGND VPWR VPWR _04937_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04868_ _05245_/A VGND VGND VPWR VPWR _05327_/A sky130_fd_sc_hd__clkbuf_4
X_07656_ _07816_/A VGND VGND VPWR VPWR _07656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07587_ _05184_/Y _07792_/A _05237_/Y _07793_/A _07586_/X VGND VGND VPWR VPWR _07595_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06607_ _09806_/Q _06604_/X _09652_/X _06606_/X VGND VGND VPWR VPWR _09806_/D sky130_fd_sc_hd__a22o_1
X_09326_ _09326_/A _09326_/B _09326_/C _09326_/D VGND VGND VPWR VPWR _09380_/D sky130_fd_sc_hd__or4_2
X_06538_ _06538_/A _06538_/B VGND VGND VPWR VPWR _06540_/A sky130_fd_sc_hd__or2_2
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09257_ _08788_/A _09256_/Y _09106_/Y VGND VGND VPWR VPWR _09257_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06469_ _06469_/A _06469_/B VGND VGND VPWR VPWR _06469_/X sky130_fd_sc_hd__or2_1
X_08208_ _08208_/A VGND VGND VPWR VPWR _08208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09188_ _09223_/B _09145_/B _09229_/B _09145_/B VGND VGND VPWR VPWR _09418_/A sky130_fd_sc_hd__o22ai_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08139_ _07017_/Y _08058_/X _07023_/Y _08059_/X _08138_/X VGND VGND VPWR VPWR _08153_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10101_ _10127_/CLK _10101_/D _07492_/B VGND VGND VPWR VPWR _10101_/Q sky130_fd_sc_hd__dfrtp_2
Xinput201 wb_sel_i[3] VGND VGND VPWR VPWR _08354_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10032_ _10135_/CLK _10032_/D _07492_/B VGND VGND VPWR VPWR _10032_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05840_ _05841_/A VGND VGND VPWR VPWR _05840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05771_ _10239_/Q _05764_/A _09660_/A1 _05765_/A VGND VGND VPWR VPWR _10239_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07510_ _09989_/Q _09988_/Q _07597_/C _07539_/A VGND VGND VPWR VPWR _07755_/A sky130_fd_sc_hd__or4_4
X_08490_ _08490_/A VGND VGND VPWR VPWR _08491_/B sky130_fd_sc_hd__clkbuf_4
X_07441_ _07441_/A VGND VGND VPWR VPWR _07441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07372_ _07370_/Y _05334_/A _07371_/Y _05785_/B VGND VGND VPWR VPWR _07372_/X sky130_fd_sc_hd__o22a_1
X_09111_ _09111_/A VGND VGND VPWR VPWR _09377_/B sky130_fd_sc_hd__inv_2
X_06323_ _09948_/Q _06315_/A _06684_/B1 _06316_/A VGND VGND VPWR VPWR _09948_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06254_ _09987_/Q _06252_/X _09578_/X _06253_/Y VGND VGND VPWR VPWR _09987_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ _09275_/A _09362_/B _09042_/C VGND VGND VPWR VPWR _09043_/A sky130_fd_sc_hd__or3_1
X_06185_ _10006_/Q VGND VGND VPWR VPWR _08045_/D sky130_fd_sc_hd__inv_2
X_05205_ _05205_/A VGND VGND VPWR VPWR _05333_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05136_ _05299_/B VGND VGND VPWR VPWR _05311_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09944_ _10257_/CLK _09944_/D repeater407/X VGND VGND VPWR VPWR _09944_/Q sky130_fd_sc_hd__dfrtp_1
X_05067_ _07483_/C VGND VGND VPWR VPWR _09680_/S sky130_fd_sc_hd__inv_4
XFILLER_131_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09875_ _10490_/CLK _09875_/D repeater404/X VGND VGND VPWR VPWR _09875_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08826_ _08837_/A _08829_/A VGND VGND VPWR VPWR _08827_/A sky130_fd_sc_hd__or2_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05969_ _05970_/A VGND VGND VPWR VPWR _05969_/X sky130_fd_sc_hd__clkbuf_2
X_08757_ _08757_/A _08858_/A VGND VGND VPWR VPWR _08898_/A sky130_fd_sc_hd__or2_1
X_08688_ _08688_/A VGND VGND VPWR VPWR _08689_/A sky130_fd_sc_hd__inv_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _09483_/A _07652_/X _09465_/A _07653_/X VGND VGND VPWR VPWR _07708_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07639_/A VGND VGND VPWR VPWR _07639_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09309_ _09309_/A _09309_/B _09309_/C _09309_/D VGND VGND VPWR VPWR _09369_/D sky130_fd_sc_hd__or4_4
XFILLER_166_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10015_ _10490_/CLK _10015_/D repeater404/X VGND VGND VPWR VPWR _10015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07990_ _08046_/A VGND VGND VPWR VPWR _08026_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06941_ _06936_/Y _06096_/B _06937_/Y _06011_/B _06940_/X VGND VGND VPWR VPWR _06960_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09660_ _10318_/Q _09660_/A1 _09679_/S VGND VGND VPWR VPWR _09660_/X sky130_fd_sc_hd__mux2_1
X_08611_ _08611_/A VGND VGND VPWR VPWR _08611_/X sky130_fd_sc_hd__clkbuf_1
X_06872_ _06870_/Y _05794_/B _06871_/Y _05138_/A VGND VGND VPWR VPWR _06872_/X sky130_fd_sc_hd__o22a_1
XFILLER_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05823_ _05823_/A VGND VGND VPWR VPWR _05823_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09591_ _09590_/X _09907_/Q _09776_/Q VGND VGND VPWR VPWR _09591_/X sky130_fd_sc_hd__mux2_1
X_05754_ _10251_/Q _05750_/X _09580_/X _05752_/X VGND VGND VPWR VPWR _10251_/D sky130_fd_sc_hd__a22o_1
X_08542_ _08921_/C _08923_/A VGND VGND VPWR VPWR _08927_/B sky130_fd_sc_hd__or2_2
XFILLER_82_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08473_ _08902_/A VGND VGND VPWR VPWR _08970_/A sky130_fd_sc_hd__clkbuf_4
X_05685_ _10292_/Q _05678_/X _09550_/A0 _05680_/X VGND VGND VPWR VPWR _10292_/D sky130_fd_sc_hd__a22o_1
X_07424_ _09785_/Q VGND VGND VPWR VPWR _07425_/B sky130_fd_sc_hd__inv_2
XFILLER_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07355_ _07350_/Y _06439_/B _07351_/Y _06430_/B _07354_/X VGND VGND VPWR VPWR _07374_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06306_ _06306_/A VGND VGND VPWR VPWR _06306_/Y sky130_fd_sc_hd__inv_2
X_07286_ _07690_/A _06266_/A _07282_/Y _06502_/A _07285_/X VGND VGND VPWR VPWR _07287_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06237_ _06237_/A VGND VGND VPWR VPWR _07551_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09025_ _09025_/A VGND VGND VPWR VPWR _09169_/A sky130_fd_sc_hd__inv_2
XFILLER_191_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06168_ _06169_/A VGND VGND VPWR VPWR _06168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06099_ _06099_/A VGND VGND VPWR VPWR _06099_/X sky130_fd_sc_hd__clkbuf_2
X_05119_ _06780_/A VGND VGND VPWR VPWR _05119_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09927_ _10000_/CLK _09927_/D repeater405/X VGND VGND VPWR VPWR _09927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09858_ _10268_/CLK _09858_/D repeater404/X VGND VGND VPWR VPWR _09858_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _10382_/CLK _09789_/D _06648_/X VGND VGND VPWR VPWR _09789_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _08809_/A _08809_/B VGND VGND VPWR VPWR _08810_/B sky130_fd_sc_hd__or2_2
XFILLER_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_125 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _05355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 _06967_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _09487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10495_ _10495_/CLK _10495_/D repeater404/X VGND VGND VPWR VPWR _10495_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05470_ _05497_/A VGND VGND VPWR VPWR _05471_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07140_ _10401_/Q VGND VGND VPWR VPWR _09459_/A sky130_fd_sc_hd__inv_6
XFILLER_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07071_ _10131_/Q VGND VGND VPWR VPWR _07071_/Y sky130_fd_sc_hd__clkinv_4
X_06022_ _10089_/Q _06013_/A _09574_/X _06014_/A VGND VGND VPWR VPWR _10089_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput313 _10458_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_2
Xoutput302 _10436_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_2
Xoutput324 _10468_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_2
Xoutput335 _09768_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_2
Xoutput346 _07502_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_2
Xoutput368 _09751_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_126_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput357 _10470_/Q VGND VGND VPWR VPWR sram_ro_clk sky130_fd_sc_hd__buf_2
Xoutput379 _09737_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09712_ _09712_/A _09477_/A VGND VGND VPWR VPWR _09712_/Z sky130_fd_sc_hd__ebufn_1
X_07973_ _07971_/Y _07639_/A _06929_/Y _07801_/A _07972_/X VGND VGND VPWR VPWR _07977_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06924_ _10059_/Q _05162_/A _10341_/Q _05126_/Y _06923_/X VGND VGND VPWR VPWR _06925_/D
+ sky130_fd_sc_hd__a221o_1
X_06855_ _06855_/A _06855_/B _06855_/C _06854_/X VGND VGND VPWR VPWR _06905_/B sky130_fd_sc_hd__or4b_2
X_09643_ _10424_/Q _07159_/X _09680_/S VGND VGND VPWR VPWR _09643_/X sky130_fd_sc_hd__mux2_1
X_09574_ input58/X _10378_/Q _10299_/Q VGND VGND VPWR VPWR _09574_/X sky130_fd_sc_hd__mux2_8
X_05806_ _05806_/A VGND VGND VPWR VPWR _05896_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08525_ _08585_/A _08959_/B VGND VGND VPWR VPWR _09379_/A sky130_fd_sc_hd__nor2_1
X_06786_ _10404_/Q VGND VGND VPWR VPWR _06786_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05737_ _10260_/Q _05730_/A _09576_/X _05731_/A VGND VGND VPWR VPWR _10260_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08456_ _08467_/A VGND VGND VPWR VPWR _08897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05668_ _06572_/A VGND VGND VPWR VPWR _06568_/A sky130_fd_sc_hd__clkbuf_2
X_08387_ _09085_/D VGND VGND VPWR VPWR _08631_/B sky130_fd_sc_hd__inv_2
X_07407_ _09921_/Q VGND VGND VPWR VPWR _07407_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07338_ _10489_/Q VGND VGND VPWR VPWR _07338_/Y sky130_fd_sc_hd__clkinv_4
X_05599_ _10340_/Q _05596_/X _09658_/A1 _05597_/Y VGND VGND VPWR VPWR _10340_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07269_ _09957_/Q VGND VGND VPWR VPWR _07269_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_191_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09008_ _09006_/B _08961_/B _09149_/A VGND VGND VPWR VPWR _09014_/B sky130_fd_sc_hd__o21ai_1
X_10280_ _10364_/CLK _10280_/D repeater410/X VGND VGND VPWR VPWR _10280_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10478_ _10478_/CLK _10478_/D _05034_/A VGND VGND VPWR VPWR _10478_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04970_ _10465_/Q _04966_/X _09580_/X _04968_/X VGND VGND VPWR VPWR _10465_/D sky130_fd_sc_hd__a22o_1
X_06640_ _09794_/Q _06636_/X _09576_/X _06637_/Y VGND VGND VPWR VPWR _09794_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06571_ _06571_/A VGND VGND VPWR VPWR _09813_/D sky130_fd_sc_hd__clkbuf_1
X_05522_ _06646_/A VGND VGND VPWR VPWR _06644_/A sky130_fd_sc_hd__clkbuf_2
X_08310_ _08310_/A _08310_/B _08310_/C _08310_/D VGND VGND VPWR VPWR _08310_/Y sky130_fd_sc_hd__nand4_2
X_09290_ _09290_/A _09290_/B _09290_/C VGND VGND VPWR VPWR _09357_/D sky130_fd_sc_hd__or3_1
X_08241_ _05332_/Y _08179_/X _05298_/Y _08180_/X VGND VGND VPWR VPWR _08241_/X sky130_fd_sc_hd__o22a_1
X_05453_ _05459_/A VGND VGND VPWR VPWR _05454_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_14 _05308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_47 _07898_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_36 _07419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _07157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _08172_/A _08172_/B _08172_/C _08172_/D VGND VGND VPWR VPWR _08172_/Y sky130_fd_sc_hd__nand4_4
XANTENNA_69 _09557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_58 input128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05384_ _09770_/Q _05671_/B input58/X _10420_/Q _05383_/X VGND VGND VPWR VPWR _10420_/D
+ sky130_fd_sc_hd__a32o_1
X_07123_ _07121_/Y _06393_/B _07122_/Y _06472_/B VGND VGND VPWR VPWR _07123_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07054_ _10074_/Q VGND VGND VPWR VPWR _07054_/Y sky130_fd_sc_hd__inv_2
X_06005_ _10101_/Q _06003_/X _09545_/A1 _06004_/Y VGND VGND VPWR VPWR _10101_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07956_ _07067_/Y _07816_/A _07092_/Y _07817_/A _07955_/X VGND VGND VPWR VPWR _07961_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06907_ _06762_/X _06906_/X _09763_/Q _06764_/X VGND VGND VPWR VPWR _09763_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07887_ _10098_/Q VGND VGND VPWR VPWR _07887_/Y sky130_fd_sc_hd__clkinv_4
X_09626_ _07860_/Y _10336_/Q _09682_/S VGND VGND VPWR VPWR _09626_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06838_ _06838_/A VGND VGND VPWR VPWR _06838_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09557_ _09919_/Q _10486_/Q _09791_/Q VGND VGND VPWR VPWR _09557_/X sky130_fd_sc_hd__mux2_4
X_06769_ input27/X _06704_/X input69/X _09679_/S _06768_/X VGND VGND VPWR VPWR _06775_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09488_ _09488_/A VGND VGND VPWR VPWR _09488_/X sky130_fd_sc_hd__clkbuf_1
X_08508_ _09006_/A VGND VGND VPWR VPWR _08883_/A sky130_fd_sc_hd__buf_2
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08439_ _08472_/B VGND VGND VPWR VPWR _09102_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10401_ _10404_/CLK _10401_/D hold41/X VGND VGND VPWR VPWR _10401_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10332_ _10336_/CLK _10332_/D repeater409/X VGND VGND VPWR VPWR _10332_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10263_ _10296_/CLK _10263_/D repeater402/X VGND VGND VPWR VPWR _10263_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10194_ _10238_/CLK _10194_/D repeater403/X VGND VGND VPWR VPWR _10194_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_132_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _10406_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_6
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_6
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_2
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_4
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08790_ _08908_/A VGND VGND VPWR VPWR _08836_/A sky130_fd_sc_hd__buf_4
X_07810_ _07810_/A _07810_/B _07810_/C _07810_/D VGND VGND VPWR VPWR _07833_/B sky130_fd_sc_hd__and4_1
X_07741_ _06981_/Y _07667_/X _07009_/Y _07668_/X VGND VGND VPWR VPWR _07741_/X sky130_fd_sc_hd__o22a_1
X_04953_ _05139_/B _05292_/A _06630_/C VGND VGND VPWR VPWR _04954_/S sky130_fd_sc_hd__or3_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_04884_ _05305_/A _05357_/A VGND VGND VPWR VPWR _04885_/A sky130_fd_sc_hd__or2_2
X_07672_ _07672_/A _07672_/B _07672_/C VGND VGND VPWR VPWR _07672_/Y sky130_fd_sc_hd__nand3_2
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09411_ _09411_/A _09411_/B _09411_/C _09411_/D VGND VGND VPWR VPWR _09444_/A sky130_fd_sc_hd__or4_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06623_ _09801_/Q _06605_/A _09646_/X _06606_/A VGND VGND VPWR VPWR _09801_/D sky130_fd_sc_hd__a22o_1
X_06554_ _09819_/Q _06552_/X _09547_/A1 _06553_/Y VGND VGND VPWR VPWR _09819_/D sky130_fd_sc_hd__a22o_1
X_09342_ _09342_/A _09342_/B _09342_/C _09342_/D VGND VGND VPWR VPWR _09421_/C sky130_fd_sc_hd__or4_2
X_05505_ _05505_/A VGND VGND VPWR VPWR _10383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ _09273_/A _09384_/C _09385_/A VGND VGND VPWR VPWR _09348_/D sky130_fd_sc_hd__or3_1
X_06485_ _09861_/Q _06482_/X _09581_/X _06484_/X VGND VGND VPWR VPWR _09861_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08224_ _06735_/Y _08177_/X _06734_/Y _08178_/X _08223_/X VGND VGND VPWR VPWR _08238_/B
+ sky130_fd_sc_hd__o221a_1
X_05436_ _05436_/A VGND VGND VPWR VPWR _05437_/A sky130_fd_sc_hd__inv_2
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08155_ _06891_/Y _08052_/X _06868_/Y _08053_/X _08154_/X VGND VGND VPWR VPWR _08172_/A
+ sky130_fd_sc_hd__o221a_1
X_05367_ _05367_/A VGND VGND VPWR VPWR _05367_/X sky130_fd_sc_hd__buf_6
X_07106_ _09515_/A _05895_/A _09469_/A _06438_/A VGND VGND VPWR VPWR _07106_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05298_ _10206_/Q VGND VGND VPWR VPWR _05298_/Y sky130_fd_sc_hd__inv_2
X_08086_ _08205_/A VGND VGND VPWR VPWR _08086_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07037_ _10446_/Q _06688_/X _10032_/Q _05080_/X _07036_/X VGND VGND VPWR VPWR _07040_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08988_ _09318_/B _08988_/B VGND VGND VPWR VPWR _08989_/C sky130_fd_sc_hd__or2_1
XFILLER_102_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07939_ _07138_/Y _07779_/A _07055_/Y _07781_/A _07938_/X VGND VGND VPWR VPWR _07939_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09609_ _09608_/X _09916_/Q _09776_/Q VGND VGND VPWR VPWR _09609_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10315_ _10504_/CLK _10315_/D repeater403/X VGND VGND VPWR VPWR _10315_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10246_ _10313_/CLK _10246_/D repeater403/X VGND VGND VPWR VPWR _10246_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10177_ _10254_/CLK _10177_/D repeater407/X VGND VGND VPWR VPWR _10177_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06270_ _06270_/A VGND VGND VPWR VPWR _06270_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05221_ _09994_/Q VGND VGND VPWR VPWR _05221_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05152_ _05157_/A _05349_/A VGND VGND VPWR VPWR _05153_/A sky130_fd_sc_hd__nor2_2
Xclkbuf_opt_8_0_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_8_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_09960_ _10238_/CLK _09960_/D repeater403/X VGND VGND VPWR VPWR _09960_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05083_ _05167_/A _05297_/B VGND VGND VPWR VPWR _06087_/B sky130_fd_sc_hd__or2_2
XFILLER_170_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08911_ _08916_/A _08911_/B VGND VGND VPWR VPWR _08911_/X sky130_fd_sc_hd__or2_2
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09891_ _10397_/CLK _09891_/D repeater409/X VGND VGND VPWR VPWR _09891_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08842_ _08842_/A _09289_/A VGND VGND VPWR VPWR _08844_/A sky130_fd_sc_hd__or2_1
Xrepeater410 hold41/A VGND VGND VPWR VPWR repeater410/X sky130_fd_sc_hd__buf_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08879_/A _08882_/A _08773_/C VGND VGND VPWR VPWR _08776_/A sky130_fd_sc_hd__and3_1
X_05985_ _10113_/Q _05981_/X _09580_/X _05983_/X VGND VGND VPWR VPWR _10113_/D sky130_fd_sc_hd__a22o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07724_ _06967_/Y _07634_/X _06948_/Y _07635_/X VGND VGND VPWR VPWR _07724_/X sky130_fd_sc_hd__o22a_1
X_04936_ _04936_/A VGND VGND VPWR VPWR _04937_/A sky130_fd_sc_hd__inv_2
XFILLER_38_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07655_ _07413_/Y _07533_/D _07369_/Y _07651_/X _07654_/X VGND VGND VPWR VPWR _07671_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06606_ _06606_/A VGND VGND VPWR VPWR _06606_/X sky130_fd_sc_hd__clkbuf_2
X_04867_ _05082_/A _05109_/B _09670_/X _09668_/X VGND VGND VPWR VPWR _05245_/A sky130_fd_sc_hd__or4_2
X_07586_ _05308_/A _07794_/A _05263_/Y _07795_/A VGND VGND VPWR VPWR _07586_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _09378_/C _09325_/B _09378_/D VGND VGND VPWR VPWR _09328_/B sky130_fd_sc_hd__or3_1
X_06537_ _06537_/A VGND VGND VPWR VPWR _06538_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06468_ _07450_/B _07481_/B VGND VGND VPWR VPWR _06468_/Y sky130_fd_sc_hd__nor2_1
X_09256_ _09256_/A _09278_/B VGND VGND VPWR VPWR _09256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08207_ _08207_/A VGND VGND VPWR VPWR _08207_/X sky130_fd_sc_hd__clkbuf_2
X_05419_ _05541_/A _05419_/B VGND VGND VPWR VPWR _05421_/A sky130_fd_sc_hd__or2_2
XFILLER_193_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06399_ _09903_/Q _06394_/X hold46/X _06395_/Y VGND VGND VPWR VPWR _09903_/D sky130_fd_sc_hd__a22o_1
X_09187_ _09416_/B _09187_/B VGND VGND VPWR VPWR _09189_/A sky130_fd_sc_hd__or2_1
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08138_ _06954_/Y _08060_/X _07009_/Y _08061_/X VGND VGND VPWR VPWR _08138_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08069_ _08188_/A VGND VGND VPWR VPWR _08069_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10100_ _10127_/CLK _10100_/D _07492_/B VGND VGND VPWR VPWR _10100_/Q sky130_fd_sc_hd__dfrtp_1
Xinput202 wb_we_i VGND VGND VPWR VPWR _08354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10031_ _10135_/CLK _10031_/D _07492_/B VGND VGND VPWR VPWR _10031_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10229_ _10355_/CLK _10229_/D repeater406/X VGND VGND VPWR VPWR _10229_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05770_ _10240_/Q _05763_/X _09550_/A0 _05765_/X VGND VGND VPWR VPWR _10240_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07440_ _07440_/A VGND VGND VPWR VPWR _07441_/A sky130_fd_sc_hd__inv_2
X_07371_ _10228_/Q VGND VGND VPWR VPWR _07371_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09110_ _08897_/B _09048_/X _08704_/C _09108_/X _09109_/X VGND VGND VPWR VPWR _09110_/X
+ sky130_fd_sc_hd__o2111a_1
X_06322_ _09949_/Q _06315_/A _06683_/B1 _06316_/A VGND VGND VPWR VPWR _09949_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09041_ _09385_/A _09041_/B VGND VGND VPWR VPWR _09042_/C sky130_fd_sc_hd__or2_1
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06253_ _06253_/A VGND VGND VPWR VPWR _06253_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05204_ _09876_/Q VGND VGND VPWR VPWR _05204_/Y sky130_fd_sc_hd__clkinv_2
X_06184_ _06184_/A _07989_/B _08010_/C VGND VGND VPWR VPWR _06184_/Y sky130_fd_sc_hd__nor3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05135_ _09663_/X _09672_/X _05135_/C VGND VGND VPWR VPWR _05299_/B sky130_fd_sc_hd__or3_4
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09943_ _10257_/CLK _09943_/D repeater407/X VGND VGND VPWR VPWR _09943_/Q sky130_fd_sc_hd__dfstp_1
X_05066_ _09808_/Q _09807_/Q _09809_/Q VGND VGND VPWR VPWR _07483_/C sky130_fd_sc_hd__or3_2
XFILLER_131_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09874_ _10490_/CLK _09874_/D repeater404/X VGND VGND VPWR VPWR _09874_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08825_ _08825_/A _09388_/A _09063_/A _09285_/A VGND VGND VPWR VPWR _08830_/A sky130_fd_sc_hd__or4_1
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08756_ _08756_/A _09248_/A VGND VGND VPWR VPWR _08758_/A sky130_fd_sc_hd__nor2_1
X_05968_ _06011_/A _05968_/B VGND VGND VPWR VPWR _05970_/A sky130_fd_sc_hd__or2_4
XFILLER_85_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04919_ _09786_/Q VGND VGND VPWR VPWR _09533_/A sky130_fd_sc_hd__inv_2
XFILLER_166_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05899_ _05899_/A VGND VGND VPWR VPWR _05899_/X sky130_fd_sc_hd__clkbuf_2
X_08687_ _08687_/A _08806_/A VGND VGND VPWR VPWR _08688_/A sky130_fd_sc_hd__or2_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _07707_/A _07707_/B _07707_/C _07707_/D VGND VGND VPWR VPWR _07717_/B sky130_fd_sc_hd__and4_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07638_ _10030_/Q VGND VGND VPWR VPWR _07638_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07569_ _07569_/A VGND VGND VPWR VPWR _09682_/S sky130_fd_sc_hd__clkbuf_8
X_09308_ _08766_/A _08578_/B _08931_/A _09004_/Y _09212_/B VGND VGND VPWR VPWR _09439_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_139_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09239_ _09180_/Y _09236_/Y _09237_/X _09167_/C VGND VGND VPWR VPWR _09326_/D sky130_fd_sc_hd__a31o_1
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10014_ _10490_/CLK _10014_/D repeater404/X VGND VGND VPWR VPWR _10014_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06940_ _06938_/Y _05785_/B _06939_/Y _06122_/B VGND VGND VPWR VPWR _06940_/X sky130_fd_sc_hd__o22a_1
X_06871_ _10120_/Q VGND VGND VPWR VPWR _06871_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08610_ _09275_/A _08610_/B VGND VGND VPWR VPWR _08611_/A sky130_fd_sc_hd__or2_1
X_05822_ _05823_/A VGND VGND VPWR VPWR _05822_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09590_ _08099_/Y _10330_/Q _09700_/S VGND VGND VPWR VPWR _09590_/X sky130_fd_sc_hd__mux2_1
X_05753_ _10252_/Q _05750_/X _09581_/X _05752_/X VGND VGND VPWR VPWR _10252_/D sky130_fd_sc_hd__a22o_1
X_08541_ _09233_/A _08561_/B _08571_/C _08556_/D VGND VGND VPWR VPWR _08923_/A sky130_fd_sc_hd__or4_4
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05684_ _10293_/Q _05678_/X _09578_/X _05680_/X VGND VGND VPWR VPWR _10293_/D sky130_fd_sc_hd__a22o_1
X_08472_ _08505_/A _08472_/B _08493_/B VGND VGND VPWR VPWR _08902_/A sky130_fd_sc_hd__or3_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07423_ _05367_/X _06762_/X _09758_/Q _06764_/A VGND VGND VPWR VPWR _09758_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07354_ _07352_/Y _06494_/B _07353_/Y _06529_/B VGND VGND VPWR VPWR _07354_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06305_ _06306_/A VGND VGND VPWR VPWR _06305_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07285_ _07283_/Y _06515_/A _07284_/Y _05541_/B VGND VGND VPWR VPWR _07285_/X sky130_fd_sc_hd__o22a_1
XFILLER_148_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06236_ _09992_/Q _06235_/Y _06227_/Y VGND VGND VPWR VPWR _09992_/D sky130_fd_sc_hd__o21ba_1
X_09024_ _09024_/A _09206_/B VGND VGND VPWR VPWR _09201_/C sky130_fd_sc_hd__nor2_1
X_06167_ _06304_/A _06167_/B VGND VGND VPWR VPWR _06169_/A sky130_fd_sc_hd__or2_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06098_ _06098_/A VGND VGND VPWR VPWR _06099_/A sky130_fd_sc_hd__inv_2
X_05118_ _05118_/A _05118_/B VGND VGND VPWR VPWR _05118_/Y sky130_fd_sc_hd__nor2_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09926_ _10000_/CLK _09926_/D repeater405/X VGND VGND VPWR VPWR _09926_/Q sky130_fd_sc_hd__dfrtp_1
X_05049_ _10427_/Q _05040_/X _09638_/X _05042_/X VGND VGND VPWR VPWR _10427_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09857_ _10268_/CLK _09857_/D repeater404/X VGND VGND VPWR VPWR _09857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _10382_/CLK _09788_/D _06650_/X VGND VGND VPWR VPWR _09788_/Q sky130_fd_sc_hd__dfrtp_4
X_08808_ _08808_/A VGND VGND VPWR VPWR _08808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08739_ _08739_/A _09100_/A VGND VGND VPWR VPWR _08742_/A sky130_fd_sc_hd__nand2_1
XANTENNA_104 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _05263_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _06967_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10494_ _10495_/CLK _10494_/D repeater404/X VGND VGND VPWR VPWR _10494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07070_ _07065_/Y _06037_/B _09509_/A _05762_/B _07069_/X VGND VGND VPWR VPWR _07089_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06021_ _10090_/Q _06013_/A hold46/X _06014_/A VGND VGND VPWR VPWR _10090_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput314 _10459_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_2
Xoutput325 _10445_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_2
Xoutput303 _10430_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_2
Xoutput347 _09539_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_2
Xoutput369 _09752_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput358 _10471_/Q VGND VGND VPWR VPWR sram_ro_csb sky130_fd_sc_hd__buf_2
Xoutput336 _09769_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_2
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07972_ _06926_/Y _07512_/A _06975_/Y _07642_/A VGND VGND VPWR VPWR _07972_/X sky130_fd_sc_hd__o22a_1
X_09711_ _10270_/Q _09475_/A VGND VGND VPWR VPWR _09711_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06923_ _10441_/Q _05091_/X input48/X _06697_/A VGND VGND VPWR VPWR _06923_/X sky130_fd_sc_hd__a22o_1
X_06854_ _06851_/Y _06705_/A _06852_/Y _05434_/B _06853_/Y VGND VGND VPWR VPWR _06854_/X
+ sky130_fd_sc_hd__o221a_1
X_09642_ _10423_/Q _07290_/X _09680_/S VGND VGND VPWR VPWR _09642_/X sky130_fd_sc_hd__mux2_1
X_09573_ input85/X input58/X _10298_/Q VGND VGND VPWR VPWR _09573_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06785_ _09839_/Q VGND VGND VPWR VPWR _06785_/Y sky130_fd_sc_hd__inv_2
X_05805_ _10219_/Q _05796_/A _09659_/A1 _05797_/A VGND VGND VPWR VPWR _10219_/D sky130_fd_sc_hd__a22o_1
X_05736_ _10261_/Q _05729_/X _09550_/A0 _05731_/X VGND VGND VPWR VPWR _10261_/D sky130_fd_sc_hd__a22o_1
X_08524_ _08746_/A _08959_/B VGND VGND VPWR VPWR _09171_/A sky130_fd_sc_hd__nor2_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05667_ _10299_/Q _06469_/A _05564_/X _04923_/A VGND VGND VPWR VPWR _10299_/D sky130_fd_sc_hd__a211o_1
X_08455_ _08621_/C _08545_/A VGND VGND VPWR VPWR _08467_/A sky130_fd_sc_hd__or2_1
X_08386_ _09348_/A VGND VGND VPWR VPWR _09275_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07406_ _10344_/Q VGND VGND VPWR VPWR _07406_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05598_ _10341_/Q _05596_/X _09545_/A1 _05597_/Y VGND VGND VPWR VPWR _10341_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07337_ _10025_/Q VGND VGND VPWR VPWR _07337_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07268_ _07263_/Y _06481_/B _07264_/Y _06095_/A _07267_/X VGND VGND VPWR VPWR _07287_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09007_ _08746_/A _08552_/B _09155_/B _08910_/X _09105_/A VGND VGND VPWR VPWR _09007_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07199_ _07194_/Y _06430_/B _07195_/Y _05550_/B _07198_/X VGND VGND VPWR VPWR _07218_/A
+ sky130_fd_sc_hd__o221a_1
X_06219_ _09992_/Q VGND VGND VPWR VPWR _06228_/B sky130_fd_sc_hd__inv_2
XFILLER_183_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09909_ _10006_/CLK _09909_/D repeater409/X VGND VGND VPWR VPWR _09909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10477_ _10478_/CLK _10477_/D _05034_/A VGND VGND VPWR VPWR _10477_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06570_ _09654_/X _09813_/Q _06575_/S VGND VGND VPWR VPWR _06571_/A sky130_fd_sc_hd__mux2_1
X_05521_ _05521_/A VGND VGND VPWR VPWR _10379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05452_ _09698_/X _05449_/X _10397_/Q _05451_/X VGND VGND VPWR VPWR _10397_/D sky130_fd_sc_hd__a22o_1
X_08240_ _05256_/Y _08219_/X _05348_/Y _08220_/X _08239_/X VGND VGND VPWR VPWR _08256_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08171_ _08171_/A _08171_/B _08171_/C _08171_/D VGND VGND VPWR VPWR _08172_/D sky130_fd_sc_hd__and4_2
XANTENNA_37 _07777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _05350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _08207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _07177_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07122_ _09865_/Q VGND VGND VPWR VPWR _07122_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 input128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05383_ _10419_/Q _05376_/X _05429_/A _06585_/A _05429_/D VGND VGND VPWR VPWR _05383_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07053_ _10110_/Q VGND VGND VPWR VPWR _09519_/A sky130_fd_sc_hd__inv_8
XFILLER_133_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06004_ _06004_/A VGND VGND VPWR VPWR _06004_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07955_ _07073_/Y _07818_/A _07954_/Y _07659_/A VGND VGND VPWR VPWR _07955_/X sky130_fd_sc_hd__o22a_1
X_06906_ _06906_/A VGND VGND VPWR VPWR _06906_/X sky130_fd_sc_hd__clkbuf_8
X_07886_ _07886_/A _07886_/B _07886_/C VGND VGND VPWR VPWR _07886_/Y sky130_fd_sc_hd__nand3_2
X_09625_ _09624_/X _09886_/Q _09776_/Q VGND VGND VPWR VPWR _09625_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06837_ _10477_/Q _06933_/B input25/X _06704_/X VGND VGND VPWR VPWR _06837_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09556_ _09779_/Q _10485_/Q _09791_/Q VGND VGND VPWR VPWR _09556_/X sky130_fd_sc_hd__mux2_4
X_06768_ input121/X _06696_/X _10335_/Q _05151_/A VGND VGND VPWR VPWR _06768_/X sky130_fd_sc_hd__a22o_2
X_09487_ _09487_/A VGND VGND VPWR VPWR _09488_/A sky130_fd_sc_hd__clkbuf_1
X_05719_ _10273_/Q _05717_/X _09588_/X _05718_/X VGND VGND VPWR VPWR _10273_/D sky130_fd_sc_hd__o22a_1
X_08507_ _08528_/B VGND VGND VPWR VPWR _09006_/A sky130_fd_sc_hd__buf_2
X_06699_ input19/X _06698_/X _10336_/Q _05151_/A VGND VGND VPWR VPWR _06699_/X sky130_fd_sc_hd__a22o_1
X_08438_ _08771_/A VGND VGND VPWR VPWR _08883_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08369_ _09788_/Q _08369_/B VGND VGND VPWR VPWR _08369_/X sky130_fd_sc_hd__and2_1
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10400_ _10405_/CLK _10400_/D hold41/X VGND VGND VPWR VPWR _10400_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10331_ _10336_/CLK _10331_/D repeater409/X VGND VGND VPWR VPWR _10331_/Q sky130_fd_sc_hd__dfrtp_2
X_10262_ _10296_/CLK _10262_/D repeater402/X VGND VGND VPWR VPWR _10262_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10193_ _10238_/CLK _10193_/D repeater403/X VGND VGND VPWR VPWR _10193_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_132_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_2
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_6
XFILLER_174_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_6
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput79 spi_enabled VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_6
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_8
XFILLER_123_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07740_ _10059_/Q VGND VGND VPWR VPWR _07740_/Y sky130_fd_sc_hd__inv_2
X_04952_ _05359_/A VGND VGND VPWR VPWR _05292_/A sky130_fd_sc_hd__buf_4
X_07671_ _07671_/A _07671_/B _07671_/C _07671_/D VGND VGND VPWR VPWR _07672_/C sky130_fd_sc_hd__and4_1
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04883_ _05173_/B VGND VGND VPWR VPWR _05357_/A sky130_fd_sc_hd__clkbuf_4
X_09410_ _09410_/A _09420_/A _08598_/A VGND VGND VPWR VPWR _09411_/B sky130_fd_sc_hd__or3b_1
XFILLER_92_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06622_ _06622_/A VGND VGND VPWR VPWR _06622_/X sky130_fd_sc_hd__clkbuf_1
X_06553_ _06553_/A VGND VGND VPWR VPWR _06553_/Y sky130_fd_sc_hd__inv_2
X_09341_ _09422_/A _09341_/B _09398_/D _09340_/X VGND VGND VPWR VPWR _09345_/A sky130_fd_sc_hd__or4b_1
Xclkbuf_opt_4_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_05504_ _09689_/X _10383_/Q _05512_/S VGND VGND VPWR VPWR _05505_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09272_ _09336_/B _09344_/B VGND VGND VPWR VPWR _09425_/B sky130_fd_sc_hd__nor2_1
X_06484_ _06484_/A VGND VGND VPWR VPWR _06484_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08223_ _06723_/Y _08179_/X _06737_/Y _08180_/X VGND VGND VPWR VPWR _08223_/X sky130_fd_sc_hd__o22a_1
X_05435_ _05436_/A VGND VGND VPWR VPWR _05435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08154_ _06857_/Y _08054_/X _06858_/Y _08055_/X VGND VGND VPWR VPWR _08154_/X sky130_fd_sc_hd__o22a_1
X_05366_ _05366_/A _05366_/B _05366_/C _05365_/X VGND VGND VPWR VPWR _05367_/A sky130_fd_sc_hd__or4b_4
XFILLER_146_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08085_ _07350_/Y _08080_/X _07319_/Y _08081_/X _08084_/X VGND VGND VPWR VPWR _08098_/B
+ sky130_fd_sc_hd__o221a_1
X_07105_ _09871_/Q VGND VGND VPWR VPWR _09469_/A sky130_fd_sc_hd__clkinv_4
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05297_ _05316_/B _05297_/B VGND VGND VPWR VPWR _05992_/A sky130_fd_sc_hd__or2_1
X_07036_ input95/X _05101_/A _09769_/Q _05146_/Y VGND VGND VPWR VPWR _07036_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08987_ _09337_/A _09045_/B _09045_/C _08986_/X VGND VGND VPWR VPWR _08988_/B sky130_fd_sc_hd__a31o_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07938_ _07098_/Y _07782_/A _07065_/Y _07783_/A VGND VGND VPWR VPWR _07938_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07869_ _10045_/Q VGND VGND VPWR VPWR _07869_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_113_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09608_ _08292_/Y _10326_/Q _09700_/S VGND VGND VPWR VPWR _09608_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09539_ input65/X VGND VGND VPWR VPWR _09539_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10314_ _10504_/CLK _10314_/D repeater404/X VGND VGND VPWR VPWR _10314_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10245_ _10313_/CLK _10245_/D repeater403/X VGND VGND VPWR VPWR _10245_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10176_ _10254_/CLK _10176_/D repeater407/X VGND VGND VPWR VPWR _10176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05220_ _05351_/A _05349_/B VGND VGND VPWR VPWR _06250_/A sky130_fd_sc_hd__or2_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05151_ _05151_/A VGND VGND VPWR VPWR _05151_/X sky130_fd_sc_hd__buf_2
XFILLER_170_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05082_ _05082_/A _05109_/B _09670_/X _05109_/D VGND VGND VPWR VPWR _05297_/B sky130_fd_sc_hd__or4_4
X_08910_ _08965_/A _09011_/A VGND VGND VPWR VPWR _08910_/X sky130_fd_sc_hd__or2_2
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09890_ _10397_/CLK _09890_/D repeater407/X VGND VGND VPWR VPWR _09890_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08849_/A _08841_/B VGND VGND VPWR VPWR _09289_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater400 _09574_/X VGND VGND VPWR VPWR _09536_/A3 sky130_fd_sc_hd__buf_12
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater411 hold41/A VGND VGND VPWR VPWR _07492_/B sky130_fd_sc_hd__buf_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08772_/A _08880_/A VGND VGND VPWR VPWR _08773_/C sky130_fd_sc_hd__and2_1
X_05984_ _10114_/Q _05981_/X _09581_/X _05983_/X VGND VGND VPWR VPWR _10114_/D sky130_fd_sc_hd__a22o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07723_ _06979_/Y _07627_/X _07023_/Y _07628_/X _07722_/X VGND VGND VPWR VPWR _07732_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04935_ _04936_/A VGND VGND VPWR VPWR _04935_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07654_ _07375_/Y _07652_/X _07357_/Y _07653_/X VGND VGND VPWR VPWR _07654_/X sky130_fd_sc_hd__o22a_1
XFILLER_65_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06605_ _06605_/A VGND VGND VPWR VPWR _06606_/A sky130_fd_sc_hd__inv_2
X_04866_ _04963_/B VGND VGND VPWR VPWR _05109_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07585_ _09989_/Q _09988_/Q _07585_/C _07602_/D VGND VGND VPWR VPWR _07795_/A sky130_fd_sc_hd__or4_4
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06536_ _09828_/Q _06530_/X _09659_/A1 _06531_/Y VGND VGND VPWR VPWR _09828_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09324_ _09324_/A _09324_/B VGND VGND VPWR VPWR _09378_/D sky130_fd_sc_hd__or2_1
XFILLER_193_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06467_ _09781_/Q _06469_/B VGND VGND VPWR VPWR _07481_/B sky130_fd_sc_hd__and2_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09255_ _09255_/A VGND VGND VPWR VPWR _09261_/A sky130_fd_sc_hd__buf_2
X_05418_ hold48/A _05397_/A input58/X _05398_/A VGND VGND VPWR VPWR _10412_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08206_ _08206_/A VGND VGND VPWR VPWR _08206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06398_ _09904_/Q _06394_/X _09576_/X _06395_/Y VGND VGND VPWR VPWR _09904_/D sky130_fd_sc_hd__a22o_1
X_09186_ _09415_/D _09186_/B VGND VGND VPWR VPWR _09187_/B sky130_fd_sc_hd__or2_1
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05349_ _05349_/A _05349_/B VGND VGND VPWR VPWR _06328_/A sky130_fd_sc_hd__or2_1
X_08137_ _06936_/Y _08052_/X _06980_/Y _08053_/X _08136_/X VGND VGND VPWR VPWR _08153_/A
+ sky130_fd_sc_hd__o221a_1
X_08068_ _08187_/A VGND VGND VPWR VPWR _08068_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07019_ _07017_/Y _06359_/A _07018_/Y _06494_/B VGND VGND VPWR VPWR _07019_/X sky130_fd_sc_hd__o22a_1
X_10030_ _10135_/CLK _10030_/D _07492_/B VGND VGND VPWR VPWR _10030_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10228_ _10355_/CLK _10228_/D repeater406/X VGND VGND VPWR VPWR _10228_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10159_ _10353_/CLK _10159_/D repeater403/X VGND VGND VPWR VPWR _10159_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2 hold2/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07370_ _10352_/Q VGND VGND VPWR VPWR _07370_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06321_ _09950_/Q _06314_/X _09658_/A1 _06316_/X VGND VGND VPWR VPWR _09950_/D sky130_fd_sc_hd__a22o_1
X_06252_ _06253_/A VGND VGND VPWR VPWR _06252_/X sky130_fd_sc_hd__clkbuf_2
X_09040_ _09040_/A _09039_/X VGND VGND VPWR VPWR _09041_/B sky130_fd_sc_hd__or2b_1
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05203_ _06780_/B _05355_/B VGND VGND VPWR VPWR _06401_/A sky130_fd_sc_hd__or2_4
XFILLER_190_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06183_ _08034_/A VGND VGND VPWR VPWR _08010_/C sky130_fd_sc_hd__clkbuf_2
X_05134_ _10115_/Q VGND VGND VPWR VPWR _05134_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09942_ _10257_/CLK _09942_/D repeater407/X VGND VGND VPWR VPWR _09942_/Q sky130_fd_sc_hd__dfrtp_1
X_05065_ _05065_/A VGND VGND VPWR VPWR _05065_/X sky130_fd_sc_hd__clkbuf_1
X_09873_ _10490_/CLK _09873_/D repeater404/X VGND VGND VPWR VPWR _09873_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08836_/A _08824_/B VGND VGND VPWR VPWR _09285_/A sky130_fd_sc_hd__nor2_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _08980_/B _09226_/A _08980_/C VGND VGND VPWR VPWR _09248_/A sky130_fd_sc_hd__and3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07706_ _09471_/A _07645_/X _07135_/Y _07533_/B _07705_/X VGND VGND VPWR VPWR _07707_/D
+ sky130_fd_sc_hd__o221a_1
X_05967_ _10123_/Q _05961_/X _09536_/A3 _05962_/Y VGND VGND VPWR VPWR _10123_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04918_ _06646_/A VGND VGND VPWR VPWR _05459_/A sky130_fd_sc_hd__clkbuf_4
X_05898_ _05898_/A VGND VGND VPWR VPWR _05899_/A sky130_fd_sc_hd__inv_2
X_08686_ _08693_/A VGND VGND VPWR VPWR _08686_/Y sky130_fd_sc_hd__inv_2
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07359_/Y _07632_/X _07325_/Y _07633_/X _07636_/X VGND VGND VPWR VPWR _07650_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_80_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04849_ _09677_/X _05715_/B VGND VGND VPWR VPWR _04852_/A sky130_fd_sc_hd__or2_4
X_07568_ _07601_/A _07568_/B _07568_/C _07568_/D VGND VGND VPWR VPWR _07569_/A sky130_fd_sc_hd__and4_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09307_ _09307_/A _09307_/B _09307_/C _08570_/X VGND VGND VPWR VPWR _09371_/C sky130_fd_sc_hd__or4b_1
X_06519_ _06519_/A VGND VGND VPWR VPWR _06519_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07499_ _10298_/Q input73/X VGND VGND VPWR VPWR _07500_/A sky130_fd_sc_hd__and2b_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09238_ _09231_/Y _09236_/Y _09237_/X _09163_/B VGND VGND VPWR VPWR _09446_/D sky130_fd_sc_hd__a31o_1
XFILLER_119_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09169_ _09169_/A _09339_/A VGND VGND VPWR VPWR _09172_/B sky130_fd_sc_hd__or2_1
XFILLER_5_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10013_ _10490_/CLK _10013_/D repeater404/X VGND VGND VPWR VPWR _10013_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06870_ _10224_/Q VGND VGND VPWR VPWR _06870_/Y sky130_fd_sc_hd__clkinv_2
X_05821_ _05874_/A _05821_/B VGND VGND VPWR VPWR _05823_/A sky130_fd_sc_hd__or2_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05752_ _05752_/A VGND VGND VPWR VPWR _05752_/X sky130_fd_sc_hd__clkbuf_2
X_08540_ _08935_/B VGND VGND VPWR VPWR _08578_/B sky130_fd_sc_hd__clkbuf_2
X_05683_ _10294_/Q _05678_/X _09579_/X _05680_/X VGND VGND VPWR VPWR _10294_/D sky130_fd_sc_hd__a22o_1
X_08471_ _08974_/B VGND VGND VPWR VPWR _08980_/B sky130_fd_sc_hd__inv_2
X_07422_ _06763_/A _07421_/X _09759_/Q _06764_/A VGND VGND VPWR VPWR _09759_/D sky130_fd_sc_hd__o22a_1
XFILLER_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07353_ _09829_/Q VGND VGND VPWR VPWR _07353_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06304_ _06304_/A _06304_/B VGND VGND VPWR VPWR _06306_/A sky130_fd_sc_hd__or2_2
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07284_ _10367_/Q VGND VGND VPWR VPWR _07284_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06235_ _09777_/Q _07534_/A _06203_/Y VGND VGND VPWR VPWR _06235_/Y sky130_fd_sc_hd__a21oi_1
X_09023_ _09023_/A VGND VGND VPWR VPWR _09206_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06166_ _06166_/A VGND VGND VPWR VPWR _06167_/B sky130_fd_sc_hd__clkbuf_4
X_06097_ _06098_/A VGND VGND VPWR VPWR _06097_/X sky130_fd_sc_hd__clkbuf_2
X_05117_ input109/X _05112_/X input52/X _05114_/X _05116_/X VGND VGND VPWR VPWR _05141_/A
+ sky130_fd_sc_hd__a221o_1
X_09925_ _10000_/CLK _09925_/D repeater405/X VGND VGND VPWR VPWR _09925_/Q sky130_fd_sc_hd__dfrtp_1
X_05048_ _05048_/A VGND VGND VPWR VPWR _05048_/X sky130_fd_sc_hd__clkbuf_1
X_09856_ _10268_/CLK _09856_/D repeater404/X VGND VGND VPWR VPWR _09856_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08807_/A VGND VGND VPWR VPWR _08808_/A sky130_fd_sc_hd__inv_2
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09787_ _10382_/CLK _09787_/D _06652_/X VGND VGND VPWR VPWR _09787_/Q sky130_fd_sc_hd__dfrtp_1
X_06999_ _09832_/Q VGND VGND VPWR VPWR _06999_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _09229_/A _08862_/A VGND VGND VPWR VPWR _09100_/A sky130_fd_sc_hd__or2_1
XANTENNA_105 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _05310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ _08737_/B _08672_/B VGND VGND VPWR VPWR _08835_/A sky130_fd_sc_hd__or2_2
XANTENNA_138 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10493_ _10495_/CLK _10493_/D repeater404/X VGND VGND VPWR VPWR _10493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06020_ _10091_/Q _06013_/A _09576_/X _06014_/A VGND VGND VPWR VPWR _10091_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput326 _10446_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_2
Xoutput304 _10437_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_2
Xoutput315 _10460_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_2
Xoutput348 _09540_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_2
XFILLER_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput359 _09867_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_2
Xoutput337 _05144_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_2
X_07971_ _10049_/Q VGND VGND VPWR VPWR _07971_/Y sky130_fd_sc_hd__inv_2
X_09710_ _10269_/Q _09473_/A VGND VGND VPWR VPWR _09710_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06922_ _10085_/Q _06692_/Y _10127_/Q _05073_/Y _06921_/X VGND VGND VPWR VPWR _06925_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06853_ _10464_/Q _06853_/B VGND VGND VPWR VPWR _06853_/Y sky130_fd_sc_hd__nand2_2
X_09641_ _10422_/Q _07421_/X _09680_/S VGND VGND VPWR VPWR _09641_/X sky130_fd_sc_hd__mux2_1
X_09572_ input83/X _09572_/A1 _10297_/Q VGND VGND VPWR VPWR _09572_/X sky130_fd_sc_hd__mux2_1
X_06784_ _10043_/Q VGND VGND VPWR VPWR _06784_/Y sky130_fd_sc_hd__clkinv_2
X_05804_ _10220_/Q _05796_/A _09661_/A1 _05797_/A VGND VGND VPWR VPWR _10220_/D sky130_fd_sc_hd__a22o_1
X_05735_ _10262_/Q _05729_/X _09547_/A1 _05731_/X VGND VGND VPWR VPWR _10262_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08523_ _08523_/A VGND VGND VPWR VPWR _08959_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05666_ _09781_/Q VGND VGND VPWR VPWR _06469_/A sky130_fd_sc_hd__inv_2
X_08454_ _08571_/C _09236_/A _09233_/A _08483_/D VGND VGND VPWR VPWR _08545_/A sky130_fd_sc_hd__or4_2
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08385_ _08999_/A _08385_/B _08491_/A VGND VGND VPWR VPWR _09348_/A sky130_fd_sc_hd__and3_1
X_07405_ _07400_/Y _05895_/A _07401_/Y _06551_/B _07404_/X VGND VGND VPWR VPWR _07418_/B
+ sky130_fd_sc_hd__o221a_2
X_05597_ _05597_/A VGND VGND VPWR VPWR _05597_/Y sky130_fd_sc_hd__inv_2
X_07336_ _07663_/A _06266_/A _07332_/Y _05830_/B _07335_/X VGND VGND VPWR VPWR _07349_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ _09006_/A _09006_/B VGND VGND VPWR VPWR _09155_/B sky130_fd_sc_hd__or2_1
X_07267_ _07265_/Y _05188_/A _07266_/Y _05775_/B VGND VGND VPWR VPWR _07267_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07198_ _07196_/Y _05474_/B _07197_/Y _06438_/A VGND VGND VPWR VPWR _07198_/X sky130_fd_sc_hd__o22a_1
X_06218_ _09993_/Q VGND VGND VPWR VPWR _07473_/A sky130_fd_sc_hd__inv_2
XFILLER_132_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06149_ _09776_/Q _09778_/Q _06147_/X _06137_/X _06148_/Y VGND VGND VPWR VPWR _10021_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09908_ _10006_/CLK _09908_/D repeater409/X VGND VGND VPWR VPWR _09908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09839_ _10364_/CLK _09839_/D repeater410/X VGND VGND VPWR VPWR _09839_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _09919_/CLK sky130_fd_sc_hd__clkbuf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10476_ _10478_/CLK _10476_/D _05034_/A VGND VGND VPWR VPWR _10476_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05520_ _09685_/X _10379_/Q _05525_/S VGND VGND VPWR VPWR _05521_/A sky130_fd_sc_hd__mux2_1
X_05451_ _05493_/D VGND VGND VPWR VPWR _05451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08170_ _06865_/Y _08092_/X _07770_/A _08093_/X _08169_/X VGND VGND VPWR VPWR _08171_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_38 _07778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _07226_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 _05365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07121_ _09905_/Q VGND VGND VPWR VPWR _07121_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_49 _09253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05382_ _06579_/D VGND VGND VPWR VPWR _06585_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07052_ input67/X VGND VGND VPWR VPWR _07052_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06003_ _06004_/A VGND VGND VPWR VPWR _06003_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07954_ _10126_/Q VGND VGND VPWR VPWR _07954_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07885_ _07885_/A _07885_/B _07885_/C _07885_/D VGND VGND VPWR VPWR _07886_/C sky130_fd_sc_hd__and4_2
XFILLER_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06905_ _06905_/A _06905_/B _06880_/X _06904_/X VGND VGND VPWR VPWR _06906_/A sky130_fd_sc_hd__or4bb_4
X_06836_ _06762_/X _06835_/X _09764_/Q _06764_/X VGND VGND VPWR VPWR _09764_/D sky130_fd_sc_hd__o22a_1
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09624_ _07833_/Y _10335_/Q _09682_/S VGND VGND VPWR VPWR _09624_/X sky130_fd_sc_hd__mux2_1
X_09555_ _09968_/Q _10484_/Q _09791_/Q VGND VGND VPWR VPWR _09555_/X sky130_fd_sc_hd__mux2_4
X_06767_ _10035_/Q _05080_/X _10087_/Q _06692_/Y _06766_/X VGND VGND VPWR VPWR _06775_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09486_ _09486_/A VGND VGND VPWR VPWR _09486_/X sky130_fd_sc_hd__clkbuf_1
X_05718_ _05718_/A VGND VGND VPWR VPWR _05718_/X sky130_fd_sc_hd__clkbuf_2
X_08506_ _09102_/A _09085_/B _09102_/C _08624_/A VGND VGND VPWR VPWR _08528_/B sky130_fd_sc_hd__or4_1
X_06698_ _06698_/A VGND VGND VPWR VPWR _06698_/X sky130_fd_sc_hd__buf_2
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08437_ _09218_/A _08771_/A VGND VGND VPWR VPWR _09363_/A sky130_fd_sc_hd__nor2_2
XFILLER_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05649_ _10309_/Q _05641_/A _09661_/A1 _05642_/A VGND VGND VPWR VPWR _10309_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08368_ _09790_/Q input186/X _09789_/Q input169/X _08367_/X VGND VGND VPWR VPWR _08368_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07319_ _10116_/Q VGND VGND VPWR VPWR _07319_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08299_ _07111_/Y _08186_/A _07153_/Y _08187_/A _08298_/X VGND VGND VPWR VPWR _08299_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_csclk clkbuf_opt_3_0_csclk/X VGND VGND VPWR VPWR _10478_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10330_ _10366_/CLK _10330_/D repeater409/X VGND VGND VPWR VPWR _10330_/Q sky130_fd_sc_hd__dfstp_2
X_10261_ _10296_/CLK _10261_/D repeater402/X VGND VGND VPWR VPWR _10261_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10192_ _10224_/CLK _10192_/D repeater405/X VGND VGND VPWR VPWR _10192_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_4
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__buf_2
XFILLER_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_2
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_12
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10459_ _10486_/CLK _10459_/D repeater409/X VGND VGND VPWR VPWR _10459_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04951_ _05027_/A _09668_/X _05082_/A _09676_/X VGND VGND VPWR VPWR _05359_/A sky130_fd_sc_hd__or4_4
X_07670_ _07326_/Y _07665_/X _07299_/Y _07666_/X _07669_/X VGND VGND VPWR VPWR _07671_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04882_ _09674_/X _09676_/X _09670_/X _05109_/D VGND VGND VPWR VPWR _05173_/B sky130_fd_sc_hd__or4_4
X_06621_ _06666_/A VGND VGND VPWR VPWR _06622_/A sky130_fd_sc_hd__clkbuf_1
X_06552_ _06553_/A VGND VGND VPWR VPWR _06552_/X sky130_fd_sc_hd__clkbuf_2
X_09340_ _08678_/X _09265_/B _09162_/B _08827_/A _09116_/Y VGND VGND VPWR VPWR _09340_/X
+ sky130_fd_sc_hd__o2111a_1
X_05503_ _05503_/A VGND VGND VPWR VPWR _05503_/X sky130_fd_sc_hd__clkbuf_1
X_09271_ _09271_/A _09271_/B VGND VGND VPWR VPWR _09425_/D sky130_fd_sc_hd__or2_2
XFILLER_21_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06483_ _06483_/A VGND VGND VPWR VPWR _06484_/A sky130_fd_sc_hd__inv_2
X_08222_ _06717_/Y _08219_/X _06748_/Y _08220_/X _08221_/X VGND VGND VPWR VPWR _08238_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05434_ _05603_/A _05434_/B VGND VGND VPWR VPWR _05436_/A sky130_fd_sc_hd__or2_2
X_05365_ _05365_/A _05365_/B _05365_/C _05365_/D VGND VGND VPWR VPWR _05365_/X sky130_fd_sc_hd__and4_4
X_08153_ _08153_/A _08153_/B _08153_/C _08153_/D VGND VGND VPWR VPWR _08153_/Y sky130_fd_sc_hd__nand4_4
X_07104_ _10162_/Q VGND VGND VPWR VPWR _09515_/A sky130_fd_sc_hd__clkinv_4
X_08084_ _07369_/Y _08082_/X _07406_/Y _08083_/X VGND VGND VPWR VPWR _08084_/X sky130_fd_sc_hd__o22a_1
X_05296_ _10102_/Q VGND VGND VPWR VPWR _05296_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07035_ _10462_/Q _06853_/B input103/X _05153_/X _07034_/X VGND VGND VPWR VPWR _07040_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08986_ _09045_/C _09096_/B _09045_/B _08985_/X VGND VGND VPWR VPWR _08986_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07937_ _07937_/A _07937_/B _07937_/C VGND VGND VPWR VPWR _07937_/Y sky130_fd_sc_hd__nand3_2
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07868_ _05291_/Y _07792_/X _05227_/Y _07793_/X _07867_/X VGND VGND VPWR VPWR _07875_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06819_ _06817_/Y _06011_/B _06818_/Y _05808_/B VGND VGND VPWR VPWR _06819_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07799_ _07799_/A VGND VGND VPWR VPWR _07799_/X sky130_fd_sc_hd__clkbuf_4
X_09607_ _09606_/X _09915_/Q _09776_/Q VGND VGND VPWR VPWR _09607_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09538_ input87/X VGND VGND VPWR VPWR _09538_/X sky130_fd_sc_hd__buf_2
XFILLER_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09469_ _09469_/A VGND VGND VPWR VPWR _09470_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10313_ _10313_/CLK _10313_/D repeater404/X VGND VGND VPWR VPWR _10313_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10244_ _10244_/CLK _10244_/D repeater402/X VGND VGND VPWR VPWR _10244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10175_ _10254_/CLK _10175_/D repeater406/X VGND VGND VPWR VPWR _10175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05150_ _05603_/B VGND VGND VPWR VPWR _05151_/A sky130_fd_sc_hd__clkinv_2
XFILLER_183_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05081_ _05081_/A VGND VGND VPWR VPWR _06776_/A sky130_fd_sc_hd__inv_2
XFILLER_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08840_ _08665_/Y _09253_/B _08839_/X VGND VGND VPWR VPWR _08842_/A sky130_fd_sc_hd__a21o_1
XFILLER_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater401 _09574_/X VGND VGND VPWR VPWR _09659_/A1 sky130_fd_sc_hd__buf_12
XFILLER_97_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08771_/A _09352_/B VGND VGND VPWR VPWR _08880_/A sky130_fd_sc_hd__or2_1
X_05983_ _05983_/A VGND VGND VPWR VPWR _05983_/X sky130_fd_sc_hd__clkbuf_2
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ _06954_/Y _07533_/C _06970_/Y _07629_/X VGND VGND VPWR VPWR _07722_/X sky130_fd_sc_hd__o22a_1
X_04934_ _04993_/A _05081_/A VGND VGND VPWR VPWR _04936_/A sky130_fd_sc_hd__or2_2
X_07653_ _07653_/A VGND VGND VPWR VPWR _07653_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04865_ _05005_/C VGND VGND VPWR VPWR _05082_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06604_ _06605_/A VGND VGND VPWR VPWR _06604_/X sky130_fd_sc_hd__clkbuf_2
X_09323_ _08753_/C _09322_/Y _08700_/A _09235_/B VGND VGND VPWR VPWR _09325_/B sky130_fd_sc_hd__a211o_1
X_07584_ _07612_/C _07584_/B VGND VGND VPWR VPWR _07794_/A sky130_fd_sc_hd__or2_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06535_ _09829_/Q _06530_/X hold46/X _06531_/Y VGND VGND VPWR VPWR _09829_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06466_ _06466_/A _06466_/B _06466_/C _06466_/D VGND VGND VPWR VPWR _06469_/B sky130_fd_sc_hd__or4_1
XFILLER_166_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09254_ _09337_/B VGND VGND VPWR VPWR _09255_/A sky130_fd_sc_hd__inv_2
X_05417_ _05417_/A VGND VGND VPWR VPWR _05417_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08205_ _08205_/A VGND VGND VPWR VPWR _08205_/X sky130_fd_sc_hd__clkbuf_2
X_09185_ _09185_/A _09433_/C VGND VGND VPWR VPWR _09186_/B sky130_fd_sc_hd__or2_1
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06397_ _09905_/Q _06394_/X _09550_/A0 _06395_/Y VGND VGND VPWR VPWR _09905_/D sky130_fd_sc_hd__a22o_1
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08136_ _06962_/Y _08054_/X _06997_/Y _08055_/X VGND VGND VPWR VPWR _08136_/X sky130_fd_sc_hd__o22a_1
X_05348_ _09941_/Q VGND VGND VPWR VPWR _05348_/Y sky130_fd_sc_hd__clkinv_2
X_05279_ _05274_/Y _06290_/A _05276_/Y _06550_/A VGND VGND VPWR VPWR _05279_/X sky130_fd_sc_hd__o22a_1
X_08067_ _08186_/A VGND VGND VPWR VPWR _08067_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07018_ _09853_/Q VGND VGND VPWR VPWR _07018_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08969_ _08969_/A _09214_/B VGND VGND VPWR VPWR _08971_/A sky130_fd_sc_hd__or2_1
XFILLER_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10227_ _10355_/CLK _10227_/D repeater406/X VGND VGND VPWR VPWR _10227_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _10283_/CLK _10158_/D repeater406/X VGND VGND VPWR VPWR _10158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3 hold3/A VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10089_ _10119_/CLK _10089_/D repeater403/X VGND VGND VPWR VPWR _10089_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06320_ _09951_/Q _06314_/X _09545_/A1 _06316_/X VGND VGND VPWR VPWR _09951_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06251_ _06304_/A _06251_/B VGND VGND VPWR VPWR _06253_/A sky130_fd_sc_hd__or2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05202_ _05338_/B VGND VGND VPWR VPWR _05355_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06182_ _10005_/Q _10004_/Q VGND VGND VPWR VPWR _08034_/A sky130_fd_sc_hd__or2_2
X_05133_ _10513_/Q VGND VGND VPWR VPWR _05133_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09941_ _10257_/CLK _09941_/D repeater407/X VGND VGND VPWR VPWR _09941_/Q sky130_fd_sc_hd__dfrtp_1
X_05064_ _05378_/A VGND VGND VPWR VPWR _05065_/A sky130_fd_sc_hd__clkbuf_1
X_09872_ _10490_/CLK _09872_/D repeater404/X VGND VGND VPWR VPWR _09872_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A _08823_/B VGND VGND VPWR VPWR _09063_/A sky130_fd_sc_hd__nor2_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08754_ _08754_/A _09415_/C VGND VGND VPWR VPWR _08756_/A sky130_fd_sc_hd__or2_1
X_05966_ _10124_/Q _05961_/X _06684_/B1 _05962_/Y VGND VGND VPWR VPWR _10124_/D sky130_fd_sc_hd__a22o_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04917_ _07450_/A VGND VGND VPWR VPWR _06646_/A sky130_fd_sc_hd__inv_2
X_07705_ _09473_/A _07646_/X _09505_/A _07647_/X VGND VGND VPWR VPWR _07705_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05897_ _05898_/A VGND VGND VPWR VPWR _05897_/X sky130_fd_sc_hd__clkbuf_2
X_08685_ _08687_/A _08685_/B VGND VGND VPWR VPWR _08693_/A sky130_fd_sc_hd__or2_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07376_/Y _07634_/X _07389_/Y _07635_/X VGND VGND VPWR VPWR _07636_/X sky130_fd_sc_hd__o22a_1
X_04848_ _05677_/B hold1/A _09678_/X VGND VGND VPWR VPWR _05715_/B sky130_fd_sc_hd__o21ai_2
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07567_ _07567_/A _07567_/B _07567_/C _07567_/D VGND VGND VPWR VPWR _07568_/D sky130_fd_sc_hd__and4_1
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09306_ _09306_/A _09306_/B _08563_/X VGND VGND VPWR VPWR _09307_/A sky130_fd_sc_hd__or3b_1
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06518_ _06518_/A VGND VGND VPWR VPWR _06519_/A sky130_fd_sc_hd__inv_2
X_09237_ _09237_/A VGND VGND VPWR VPWR _09237_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07498_ _07498_/A VGND VGND VPWR VPWR _07498_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06449_ _09869_/Q _06441_/A _09661_/A1 _06442_/A VGND VGND VPWR VPWR _09869_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09168_ _09168_/A VGND VGND VPWR VPWR _09339_/A sky130_fd_sc_hd__inv_2
X_09099_ _09109_/B VGND VGND VPWR VPWR _09099_/X sky130_fd_sc_hd__buf_2
X_08119_ _09495_/A _08054_/X _09455_/A _08055_/X _08118_/X VGND VGND VPWR VPWR _08135_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10012_ _10495_/CLK _10012_/D repeater404/X VGND VGND VPWR VPWR _10012_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05820_ _05820_/A VGND VGND VPWR VPWR _05821_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05751_ _05751_/A VGND VGND VPWR VPWR _05752_/A sky130_fd_sc_hd__inv_2
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05682_ _10295_/Q _05678_/X _09580_/X _05680_/X VGND VGND VPWR VPWR _10295_/D sky130_fd_sc_hd__a22o_1
X_08470_ _08571_/C _09236_/A _09295_/A _08561_/B VGND VGND VPWR VPWR _08974_/B sky130_fd_sc_hd__or4_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07421_ _07421_/A VGND VGND VPWR VPWR _07421_/X sky130_fd_sc_hd__buf_6
X_07352_ _09850_/Q VGND VGND VPWR VPWR _07352_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06303_ _06303_/A VGND VGND VPWR VPWR _06304_/B sky130_fd_sc_hd__buf_2
XFILLER_31_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07283_ _09835_/Q VGND VGND VPWR VPWR _07283_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06234_ _06234_/A VGND VGND VPWR VPWR _09993_/D sky130_fd_sc_hd__inv_2
X_09022_ _09022_/A _09198_/C _09309_/C VGND VGND VPWR VPWR _09022_/X sky130_fd_sc_hd__or3_1
XFILLER_163_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06165_ _10012_/Q _06156_/A _09659_/A1 _06157_/A VGND VGND VPWR VPWR _10012_/D sky130_fd_sc_hd__a22o_1
X_05116_ _10471_/Q _04947_/Y input34/X _06838_/A VGND VGND VPWR VPWR _05116_/X sky130_fd_sc_hd__a22o_1
X_06096_ _06108_/A _06096_/B VGND VGND VPWR VPWR _06098_/A sky130_fd_sc_hd__or2_2
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09924_ _10000_/CLK _09924_/D repeater405/X VGND VGND VPWR VPWR _09924_/Q sky130_fd_sc_hd__dfrtp_1
X_05047_ _05053_/A VGND VGND VPWR VPWR _05048_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09855_ _10268_/CLK _09855_/D repeater404/X VGND VGND VPWR VPWR _09855_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_112_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08806_/A VGND VGND VPWR VPWR _08806_/Y sky130_fd_sc_hd__inv_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09786_ _10382_/CLK _09786_/D _06654_/X VGND VGND VPWR VPWR _09786_/Q sky130_fd_sc_hd__dfrtp_1
X_06998_ _10158_/Q VGND VGND VPWR VPWR _06998_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08737_ _08786_/B _08737_/B VGND VGND VPWR VPWR _08862_/A sky130_fd_sc_hd__or2_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05949_ _10135_/Q _05942_/A _06683_/B1 _05943_/A VGND VGND VPWR VPWR _10135_/D sky130_fd_sc_hd__a22o_1
XANTENNA_106 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 input88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ _08668_/A _09092_/B VGND VGND VPWR VPWR _08737_/B sky130_fd_sc_hd__or2_4
XFILLER_121_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _07778_/A VGND VGND VPWR VPWR _07619_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08599_ _09102_/B _08998_/A _08598_/X VGND VGND VPWR VPWR _08600_/B sky130_fd_sc_hd__o21ai_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10492_ _10495_/CLK _10492_/D repeater404/X VGND VGND VPWR VPWR _10492_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput305 _10438_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_2
Xoutput316 _10461_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput338 _09522_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput327 _10447_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_2
Xoutput349 _10472_/Q VGND VGND VPWR VPWR sram_ro_addr[0] sky130_fd_sc_hd__buf_2
X_07970_ _06969_/Y _07792_/A _07004_/Y _07793_/A _07969_/X VGND VGND VPWR VPWR _07977_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_141_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06921_ input119/X _06696_/A input96/X _05101_/A VGND VGND VPWR VPWR _06921_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06852_ _10403_/Q VGND VGND VPWR VPWR _06852_/Y sky130_fd_sc_hd__inv_2
X_09640_ _10427_/Q _06835_/X _09680_/S VGND VGND VPWR VPWR _09640_/X sky130_fd_sc_hd__mux2_1
X_06783_ _09826_/Q VGND VGND VPWR VPWR _06783_/Y sky130_fd_sc_hd__clkinv_4
X_09571_ input84/X input67/X _10298_/Q VGND VGND VPWR VPWR _09571_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05803_ _10221_/Q _05796_/A _09660_/A1 _05797_/A VGND VGND VPWR VPWR _10221_/D sky130_fd_sc_hd__a22o_1
X_05734_ _10263_/Q _05729_/X _09579_/X _05731_/X VGND VGND VPWR VPWR _10263_/D sky130_fd_sc_hd__a22o_1
X_08522_ _09155_/A _08957_/A VGND VGND VPWR VPWR _08523_/A sky130_fd_sc_hd__or2_1
X_08453_ _08530_/D VGND VGND VPWR VPWR _08483_/D sky130_fd_sc_hd__buf_2
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05665_ _05665_/A VGND VGND VPWR VPWR _05665_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07404_ _07402_/Y _05874_/B _07403_/Y _05314_/A VGND VGND VPWR VPWR _07404_/X sky130_fd_sc_hd__o22a_1
X_08384_ _09102_/D VGND VGND VPWR VPWR _08491_/A sky130_fd_sc_hd__inv_2
X_05596_ _05597_/A VGND VGND VPWR VPWR _05596_/X sky130_fd_sc_hd__clkbuf_2
X_07335_ _07333_/Y _06329_/B _07907_/A _06280_/B VGND VGND VPWR VPWR _07335_/X sky130_fd_sc_hd__o22a_1
X_07266_ _10234_/Q VGND VGND VPWR VPWR _07266_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09005_ _09005_/A VGND VGND VPWR VPWR _09204_/A sky130_fd_sc_hd__buf_2
X_06217_ _09994_/Q _06208_/A _09659_/A1 _06209_/A VGND VGND VPWR VPWR _09994_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07197_ _09870_/Q VGND VGND VPWR VPWR _07197_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06148_ _06137_/A _06150_/A _06260_/C VGND VGND VPWR VPWR _06148_/Y sky130_fd_sc_hd__o21ai_1
X_06079_ _06087_/A _06079_/B VGND VGND VPWR VPWR _06081_/A sky130_fd_sc_hd__or2_1
X_09907_ _10023_/CLK _09907_/D repeater409/X VGND VGND VPWR VPWR _09907_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _10191_/CLK _09838_/D repeater410/X VGND VGND VPWR VPWR _09838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09769_ _10127_/CLK _09769_/D VGND VGND VPWR VPWR _09769_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10475_ _10478_/CLK _10475_/D _05034_/A VGND VGND VPWR VPWR _10475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05450_ _05450_/A VGND VGND VPWR VPWR _05493_/D sky130_fd_sc_hd__inv_2
XANTENNA_28 _07237_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05381_ _09770_/Q VGND VGND VPWR VPWR _06579_/D sky130_fd_sc_hd__inv_2
XANTENNA_17 _06931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _07590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07120_ _09963_/Q VGND VGND VPWR VPWR _09479_/A sky130_fd_sc_hd__clkinv_4
XFILLER_173_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07051_ _07049_/Y _05603_/B _07050_/Y _06024_/B VGND VGND VPWR VPWR _07051_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06002_ _06087_/A _06002_/B VGND VGND VPWR VPWR _06004_/A sky130_fd_sc_hd__or2_1
XFILLER_141_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07953_ _07141_/Y _07532_/A _07146_/Y _07811_/A _07952_/X VGND VGND VPWR VPWR _07961_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06904_ _06881_/Y _06481_/B _06884_/X _06890_/X _06903_/X VGND VGND VPWR VPWR _06904_/X
+ sky130_fd_sc_hd__o2111a_2
X_07884_ _05254_/Y _07825_/X _05175_/Y _07827_/X _07883_/X VGND VGND VPWR VPWR _07885_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09623_ _09622_/X _09885_/Q _09776_/Q VGND VGND VPWR VPWR _09623_/X sky130_fd_sc_hd__mux2_1
X_06835_ _06835_/A VGND VGND VPWR VPWR _06835_/X sky130_fd_sc_hd__buf_4
XFILLER_102_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06766_ _10465_/Q _06853_/B _10457_/Q _05089_/A VGND VGND VPWR VPWR _06766_/X sky130_fd_sc_hd__a22o_1
X_09554_ _09982_/Q _10483_/Q _09791_/Q VGND VGND VPWR VPWR _09554_/X sky130_fd_sc_hd__mux2_8
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ _09485_/A VGND VGND VPWR VPWR _09486_/A sky130_fd_sc_hd__clkbuf_1
X_08505_ _08505_/A VGND VGND VPWR VPWR _09102_/A sky130_fd_sc_hd__clkbuf_2
X_05717_ _05717_/A VGND VGND VPWR VPWR _05717_/X sky130_fd_sc_hd__clkbuf_2
X_06697_ _06697_/A VGND VGND VPWR VPWR _06697_/X sky130_fd_sc_hd__buf_2
X_08436_ _08774_/A _08775_/A VGND VGND VPWR VPWR _08771_/A sky130_fd_sc_hd__or2_2
X_05648_ _10310_/Q _05641_/A _09660_/A1 _05642_/A VGND VGND VPWR VPWR _10310_/D sky130_fd_sc_hd__a22o_1
X_08367_ _09788_/Q _08367_/B VGND VGND VPWR VPWR _08367_/X sky130_fd_sc_hd__and2_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07318_ _10008_/Q VGND VGND VPWR VPWR _07318_/Y sky130_fd_sc_hd__clkinv_2
X_05579_ _05579_/A VGND VGND VPWR VPWR _05579_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08298_ _07073_/Y _08188_/A _07074_/Y _08189_/A VGND VGND VPWR VPWR _08298_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07249_ _07244_/Y _04871_/B _07245_/Y _05807_/A _07248_/X VGND VGND VPWR VPWR _07262_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_191_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10260_ _10289_/CLK _10260_/D repeater402/X VGND VGND VPWR VPWR _10260_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10191_ _10191_/CLK _10191_/D repeater410/X VGND VGND VPWR VPWR _10191_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_6
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_8
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10458_ _10486_/CLK _10458_/D repeater409/X VGND VGND VPWR VPWR _10458_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_184_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10389_ _10500_/CLK _10389_/D repeater407/X VGND VGND VPWR VPWR _10389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04950_ _09678_/X _04947_/Y _06684_/B1 _10470_/Q _04948_/X VGND VGND VPWR VPWR _10470_/D
+ sky130_fd_sc_hd__a32o_1
X_04881_ _05318_/B VGND VGND VPWR VPWR _05305_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06620_ _09802_/Q _06604_/X _09647_/X _06606_/X VGND VGND VPWR VPWR _09802_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06551_ _06635_/A _06551_/B VGND VGND VPWR VPWR _06553_/A sky130_fd_sc_hd__or2_1
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05502_ _05518_/A VGND VGND VPWR VPWR _05503_/A sky130_fd_sc_hd__clkbuf_1
X_06482_ _06483_/A VGND VGND VPWR VPWR _06482_/X sky130_fd_sc_hd__clkbuf_2
X_09270_ _09270_/A _09421_/A _09343_/B _09400_/B VGND VGND VPWR VPWR _09274_/A sky130_fd_sc_hd__or4_1
XFILLER_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ _06751_/Y _08173_/X _06708_/A _08174_/X VGND VGND VPWR VPWR _08221_/X sky130_fd_sc_hd__o22a_1
X_05433_ _05433_/A VGND VGND VPWR VPWR _05434_/B sky130_fd_sc_hd__buf_4
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08152_ _08152_/A _08152_/B _08152_/C _08152_/D VGND VGND VPWR VPWR _08153_/D sky130_fd_sc_hd__and4_2
X_05364_ _05364_/A _05364_/B _05364_/C _05364_/D VGND VGND VPWR VPWR _05365_/D sky130_fd_sc_hd__and4_1
XFILLER_173_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05295_ _05329_/A _05311_/B VGND VGND VPWR VPWR _05838_/A sky130_fd_sc_hd__or2_4
X_08083_ _08202_/A VGND VGND VPWR VPWR _08083_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07103_ _10360_/Q VGND VGND VPWR VPWR _09457_/A sky130_fd_sc_hd__inv_4
X_07034_ _10048_/Q _05084_/Y _10440_/Q _05091_/X VGND VGND VPWR VPWR _07034_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _08997_/A _08985_/B VGND VGND VPWR VPWR _08985_/X sky130_fd_sc_hd__or2_1
XFILLER_114_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07936_ _07936_/A _07936_/B _07936_/C _07936_/D VGND VGND VPWR VPWR _07937_/C sky130_fd_sc_hd__and4_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07867_ _05267_/Y _07794_/X _05260_/Y _07795_/X VGND VGND VPWR VPWR _07867_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06818_ _10217_/Q VGND VGND VPWR VPWR _06818_/Y sky130_fd_sc_hd__clkinv_2
X_09606_ _08274_/Y _10325_/Q _09700_/S VGND VGND VPWR VPWR _09606_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07798_ _10035_/Q VGND VGND VPWR VPWR _07798_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06749_ _06747_/Y _06439_/B _06748_/Y _06313_/B VGND VGND VPWR VPWR _06749_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09468_ _09468_/A VGND VGND VPWR VPWR _09468_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08419_ _08640_/A VGND VGND VPWR VPWR _08695_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09399_ _09432_/A _09399_/B _09399_/C VGND VGND VPWR VPWR _09425_/C sky130_fd_sc_hd__or3_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10312_ _10313_/CLK _10312_/D repeater404/X VGND VGND VPWR VPWR _10312_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10243_ _10244_/CLK _10243_/D repeater402/X VGND VGND VPWR VPWR _10243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10174_ _10313_/CLK _10174_/D repeater403/X VGND VGND VPWR VPWR _10174_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05080_ _05080_/A VGND VGND VPWR VPWR _05080_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater402 repeater403/X VGND VGND VPWR VPWR repeater402/X sky130_fd_sc_hd__buf_12
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08853_/B VGND VGND VPWR VPWR _09352_/B sky130_fd_sc_hd__clkbuf_4
X_05982_ _05982_/A VGND VGND VPWR VPWR _05983_/A sky130_fd_sc_hd__inv_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07721_ _06943_/Y _07618_/X _06987_/Y _07619_/X _07720_/X VGND VGND VPWR VPWR _07744_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04933_ _05118_/A _05261_/B VGND VGND VPWR VPWR _05081_/A sky130_fd_sc_hd__or2_1
X_04864_ _05318_/B VGND VGND VPWR VPWR _05313_/A sky130_fd_sc_hd__clkbuf_2
X_07652_ _07812_/A VGND VGND VPWR VPWR _07652_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07583_ _07583_/A VGND VGND VPWR VPWR _07793_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_51_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _10487_/CLK sky130_fd_sc_hd__clkbuf_16
X_06603_ _09773_/Q _06602_/X _06585_/A VGND VGND VPWR VPWR _06605_/A sky130_fd_sc_hd__o21ai_4
X_06534_ _09830_/Q _06530_/X _09660_/A1 _06531_/Y VGND VGND VPWR VPWR _09830_/D sky130_fd_sc_hd__a22o_1
X_09322_ _08483_/D _08552_/X _08548_/A VGND VGND VPWR VPWR _09322_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06465_ _08492_/C _06465_/B _06465_/C _06464_/X VGND VGND VPWR VPWR _06466_/D sky130_fd_sc_hd__or4b_1
X_09253_ _09253_/A _09253_/B _09253_/C VGND VGND VPWR VPWR _09337_/B sky130_fd_sc_hd__or3_2
X_06396_ _09906_/Q _06394_/X _09578_/X _06395_/Y VGND VGND VPWR VPWR _09906_/D sky130_fd_sc_hd__a22o_1
X_05416_ _05588_/A VGND VGND VPWR VPWR _05417_/A sky130_fd_sc_hd__clkbuf_1
X_09184_ _09184_/A _09184_/B VGND VGND VPWR VPWR _09433_/C sky130_fd_sc_hd__or2_2
X_08204_ _06790_/Y _08199_/X _06823_/Y _08200_/X _08203_/X VGND VGND VPWR VPWR _08217_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05347_ _05347_/A VGND VGND VPWR VPWR _05419_/B sky130_fd_sc_hd__buf_4
X_08135_ _08135_/A _08135_/B _08135_/C _08135_/D VGND VGND VPWR VPWR _08135_/Y sky130_fd_sc_hd__nand4_4
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05278_ _05349_/A _05359_/B VGND VGND VPWR VPWR _06550_/A sky130_fd_sc_hd__or2_1
X_08066_ _07377_/Y _08065_/X _07375_/Y _06188_/X VGND VGND VPWR VPWR _08066_/X sky130_fd_sc_hd__o22a_1
X_07017_ _09924_/Q VGND VGND VPWR VPWR _07017_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08968_ _09046_/A _08968_/B VGND VGND VPWR VPWR _09214_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08899_ _09057_/A VGND VGND VPWR VPWR _09277_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07919_ _07231_/Y _07794_/X _07215_/Y _07795_/X VGND VGND VPWR VPWR _07919_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10244_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10226_ _10349_/CLK _10226_/D repeater405/X VGND VGND VPWR VPWR _10226_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10157_ _10157_/CLK _10157_/D repeater406/X VGND VGND VPWR VPWR _10157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10088_ _10374_/CLK _10088_/D hold41/X VGND VGND VPWR VPWR _10088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xnet399_2 net399_2/A VGND VGND VPWR VPWR _07505_/A sky130_fd_sc_hd__inv_2
XFILLER_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06250_ _06250_/A VGND VGND VPWR VPWR _06251_/B sky130_fd_sc_hd__buf_4
XFILLER_175_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05201_ _05213_/A _05213_/B _05201_/C VGND VGND VPWR VPWR _05338_/B sky130_fd_sc_hd__or3_2
X_06181_ _08038_/A VGND VGND VPWR VPWR _07989_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05132_ _09946_/Q _06633_/A _10337_/Q _05126_/Y _05131_/X VGND VGND VPWR VPWR _05141_/C
+ sky130_fd_sc_hd__a221o_1
X_09940_ _10310_/CLK _09940_/D repeater403/X VGND VGND VPWR VPWR _09940_/Q sky130_fd_sc_hd__dfrtp_1
X_05063_ _10423_/Q _05041_/A _09641_/X _05042_/A VGND VGND VPWR VPWR _10423_/D sky130_fd_sc_hd__a22o_1
X_09871_ _10490_/CLK _09871_/D repeater404/X VGND VGND VPWR VPWR _09871_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08822_ _08823_/A _08822_/B VGND VGND VPWR VPWR _09388_/A sky130_fd_sc_hd__nor2_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08753_ _09226_/A _08753_/B _08753_/C VGND VGND VPWR VPWR _09415_/C sky130_fd_sc_hd__and3_1
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05965_ _10125_/Q _05961_/X _06683_/B1 _05962_/Y VGND VGND VPWR VPWR _10125_/D sky130_fd_sc_hd__a22o_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04916_ _10482_/Q _04915_/Y _09536_/A3 _04915_/A _09678_/X VGND VGND VPWR VPWR _10482_/D
+ sky130_fd_sc_hd__o221a_1
X_07704_ _07503_/Y _07639_/X _09517_/A _07641_/X _07703_/X VGND VGND VPWR VPWR _07707_/C
+ sky130_fd_sc_hd__o221a_1
X_05896_ _05896_/A _05896_/B VGND VGND VPWR VPWR _05898_/A sky130_fd_sc_hd__or2_2
X_08684_ _08684_/A _09048_/A VGND VGND VPWR VPWR _09324_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _07795_/A VGND VGND VPWR VPWR _07635_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04847_ _04847_/A VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__buf_6
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07566_ _07579_/A _07653_/A _07572_/A _07573_/A VGND VGND VPWR VPWR _07567_/D sky130_fd_sc_hd__and4_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09305_ _08491_/B _09303_/Y _09353_/A _09209_/C VGND VGND VPWR VPWR _09407_/D sky130_fd_sc_hd__a211o_1
X_06517_ _06518_/A VGND VGND VPWR VPWR _06517_/X sky130_fd_sc_hd__clkbuf_2
X_09236_ _09236_/A _09236_/B VGND VGND VPWR VPWR _09236_/Y sky130_fd_sc_hd__nor2_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07497_ _07497_/A VGND VGND VPWR VPWR _07498_/A sky130_fd_sc_hd__buf_2
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06448_ _09870_/Q _06441_/A _09660_/A1 _06442_/A VGND VGND VPWR VPWR _09870_/D sky130_fd_sc_hd__a22o_1
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06379_ _06374_/X _09605_/X _09650_/X _09915_/Q VGND VGND VPWR VPWR _09915_/D sky130_fd_sc_hd__o22a_1
X_09167_ _09167_/A _09446_/C _09167_/C _09326_/C VGND VGND VPWR VPWR _09172_/A sky130_fd_sc_hd__or4_1
XFILLER_134_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09098_ _09098_/A VGND VGND VPWR VPWR _09109_/B sky130_fd_sc_hd__clkbuf_2
X_08118_ _09487_/A _08219_/A _09477_/A _08220_/A VGND VGND VPWR VPWR _08118_/X sky130_fd_sc_hd__o22a_1
XFILLER_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08049_ _08049_/A _08049_/B _08049_/C _08049_/D VGND VGND VPWR VPWR _08050_/D sky130_fd_sc_hd__and4_1
XFILLER_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10011_ _10500_/CLK _10011_/D repeater407/X VGND VGND VPWR VPWR _10011_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10209_ _10355_/CLK _10209_/D repeater406/X VGND VGND VPWR VPWR _10209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05750_ _05751_/A VGND VGND VPWR VPWR _05750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05681_ _10296_/Q _05678_/X _09581_/X _05680_/X VGND VGND VPWR VPWR _10296_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07420_ _07420_/A _07420_/B _07419_/X VGND VGND VPWR VPWR _07421_/A sky130_fd_sc_hd__or3b_2
X_07351_ _09877_/Q VGND VGND VPWR VPWR _07351_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06302_ _09960_/Q _06293_/A _09659_/A1 _06294_/A VGND VGND VPWR VPWR _09960_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07282_ _09843_/Q VGND VGND VPWR VPWR _07282_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_31_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06233_ _07473_/A _06177_/Y _06227_/Y _06184_/A _06232_/X VGND VGND VPWR VPWR _06234_/A
+ sky130_fd_sc_hd__o32a_1
X_09021_ _09021_/A _09021_/B VGND VGND VPWR VPWR _09309_/C sky130_fd_sc_hd__or2_1
XFILLER_191_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06164_ _10013_/Q _06156_/A _09661_/A1 _06157_/A VGND VGND VPWR VPWR _10013_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05115_ _05163_/B _05284_/B VGND VGND VPWR VPWR _06838_/A sky130_fd_sc_hd__nor2_2
XFILLER_144_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06095_ _06095_/A VGND VGND VPWR VPWR _06096_/B sky130_fd_sc_hd__clkbuf_4
X_09923_ _10000_/CLK _09923_/D repeater405/X VGND VGND VPWR VPWR _09923_/Q sky130_fd_sc_hd__dfrtp_1
X_05046_ _10428_/Q _05040_/X _09640_/X _05042_/X VGND VGND VPWR VPWR _10428_/D sky130_fd_sc_hd__a22o_1
X_09854_ _10490_/CLK _09854_/D repeater404/X VGND VGND VPWR VPWR _09854_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08805_ _08819_/B _08823_/B VGND VGND VPWR VPWR _09060_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _10382_/CLK _09785_/D _06656_/X VGND VGND VPWR VPWR _09785_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06997_ _10374_/Q VGND VGND VPWR VPWR _06997_/Y sky130_fd_sc_hd__clkinv_4
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _08736_/A VGND VGND VPWR VPWR _09229_/A sky130_fd_sc_hd__buf_2
X_05948_ _10136_/Q _05941_/X _09658_/A1 _05943_/X VGND VGND VPWR VPWR _10136_/D sky130_fd_sc_hd__a22o_1
XANTENNA_107 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ _08667_/A _08781_/B VGND VGND VPWR VPWR _09092_/B sky130_fd_sc_hd__or2b_1
X_05879_ _10177_/Q _05875_/X _09576_/X _05876_/Y VGND VGND VPWR VPWR _10177_/D sky130_fd_sc_hd__a22o_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07777_/A VGND VGND VPWR VPWR _07618_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08598_ _08598_/A _08598_/B VGND VGND VPWR VPWR _08598_/X sky130_fd_sc_hd__and2_1
XFILLER_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07549_ _07582_/B _07549_/B VGND VGND VPWR VPWR _07789_/A sky130_fd_sc_hd__or2_1
XFILLER_167_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09219_ _08385_/B _09278_/B _09299_/A _09385_/A VGND VGND VPWR VPWR _09220_/D sky130_fd_sc_hd__a211o_1
X_10491_ _10491_/CLK _10491_/D repeater403/X VGND VGND VPWR VPWR _10491_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput306 _10439_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_2
Xoutput317 _10462_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_2
XFILLER_141_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput328 _10448_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_2
Xoutput339 _09554_/X VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_2
XFILLER_141_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06920_ _09572_/A1 _06693_/A input65/X _06844_/X _06919_/X VGND VGND VPWR VPWR _06925_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06851_ _10138_/Q VGND VGND VPWR VPWR _06851_/Y sky130_fd_sc_hd__inv_2
X_09570_ _07503_/Y input92/X input76/X VGND VGND VPWR VPWR _09570_/X sky130_fd_sc_hd__mux2_2
XFILLER_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06782_ input98/X _05101_/X input116/X _05112_/X _06781_/Y VGND VGND VPWR VPWR _06789_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05802_ _10222_/Q _05795_/X _09550_/A0 _05797_/X VGND VGND VPWR VPWR _10222_/D sky130_fd_sc_hd__a22o_1
X_05733_ _10264_/Q _05729_/X _09580_/X _05731_/X VGND VGND VPWR VPWR _10264_/D sky130_fd_sc_hd__a22o_1
X_08521_ _09233_/A _08561_/B _08537_/C _09236_/A VGND VGND VPWR VPWR _08957_/A sky130_fd_sc_hd__or4_4
X_08452_ _09372_/C _08812_/A VGND VGND VPWR VPWR _09299_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05664_ _06644_/A VGND VGND VPWR VPWR _05665_/A sky130_fd_sc_hd__clkbuf_1
X_07403_ _10254_/Q VGND VGND VPWR VPWR _07403_/Y sky130_fd_sc_hd__clkinv_2
X_08383_ _08687_/A VGND VGND VPWR VPWR _09102_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05595_ _05775_/A _05595_/B VGND VGND VPWR VPWR _05597_/A sky130_fd_sc_hd__or2_1
X_07334_ _09970_/Q VGND VGND VPWR VPWR _07907_/A sky130_fd_sc_hd__clkinv_4
XFILLER_176_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07265_ _10229_/Q VGND VGND VPWR VPWR _07265_/Y sky130_fd_sc_hd__inv_2
X_09004_ _09159_/A _09354_/B VGND VGND VPWR VPWR _09004_/Y sky130_fd_sc_hd__nor2_2
X_06216_ _09995_/Q _06208_/A _09661_/A1 _06209_/A VGND VGND VPWR VPWR _09995_/D sky130_fd_sc_hd__a22o_1
X_07196_ _10388_/Q VGND VGND VPWR VPWR _07196_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06147_ _06227_/B VGND VGND VPWR VPWR _06147_/X sky130_fd_sc_hd__buf_2
X_06078_ _06078_/A VGND VGND VPWR VPWR _06079_/B sky130_fd_sc_hd__clkbuf_4
X_09906_ _10119_/CLK _09906_/D repeater403/X VGND VGND VPWR VPWR _09906_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05029_ _06780_/A _05355_/A VGND VGND VPWR VPWR _05031_/B sky130_fd_sc_hd__or2_1
XFILLER_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _10191_/CLK _09837_/D repeater410/X VGND VGND VPWR VPWR _09837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09768_ _10127_/CLK _09768_/D VGND VGND VPWR VPWR _09768_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08719_ _08719_/A _09326_/B VGND VGND VPWR VPWR _08721_/A sky130_fd_sc_hd__nor2_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09699_ _05677_/B hold1/A _09699_/S VGND VGND VPWR VPWR _09699_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10474_ _10478_/CLK _10474_/D _05034_/A VGND VGND VPWR VPWR _10474_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_29 _07932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05380_ _09809_/Q _09808_/Q _06579_/B VGND VGND VPWR VPWR _05671_/B sky130_fd_sc_hd__and3_1
XANTENNA_18 _06932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07050_ _10084_/Q VGND VGND VPWR VPWR _07050_/Y sky130_fd_sc_hd__inv_6
XFILLER_146_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06001_ _06327_/A VGND VGND VPWR VPWR _06087_/A sky130_fd_sc_hd__buf_4
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07952_ _07086_/Y _07812_/A _07048_/Y _07653_/A VGND VGND VPWR VPWR _07952_/X sky130_fd_sc_hd__o22a_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07883_ _05208_/Y _07828_/X _05298_/Y _07829_/X VGND VGND VPWR VPWR _07883_/X sky130_fd_sc_hd__o22a_1
X_06903_ _06891_/Y _06096_/B _06893_/X _06896_/X _06902_/X VGND VGND VPWR VPWR _06903_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09622_ _07776_/Y _10334_/Q _09682_/S VGND VGND VPWR VPWR _09622_/X sky130_fd_sc_hd__mux2_1
X_06834_ _06834_/A _06834_/B _06814_/X _06833_/X VGND VGND VPWR VPWR _06835_/A sky130_fd_sc_hd__or4bb_4
X_09553_ _09579_/X _10305_/Q _09677_/S VGND VGND VPWR VPWR _09553_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08504_ _08620_/A _08504_/B VGND VGND VPWR VPWR _08598_/A sky130_fd_sc_hd__or2_2
XFILLER_102_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06765_ _06759_/X _06762_/X _09765_/Q _06764_/X VGND VGND VPWR VPWR _09765_/D sky130_fd_sc_hd__o22a_1
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09484_ _09484_/A VGND VGND VPWR VPWR _09484_/X sky130_fd_sc_hd__clkbuf_1
X_05716_ _05718_/A VGND VGND VPWR VPWR _05717_/A sky130_fd_sc_hd__inv_2
XFILLER_102_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06696_ _06696_/A VGND VGND VPWR VPWR _06696_/X sky130_fd_sc_hd__buf_2
X_08435_ _09247_/C _09224_/B VGND VGND VPWR VPWR _08775_/A sky130_fd_sc_hd__or2_4
X_05647_ _10311_/Q _05640_/X _09550_/A0 _05642_/X VGND VGND VPWR VPWR _10311_/D sky130_fd_sc_hd__a22o_1
X_08366_ _09790_/Q input185/X _09789_/Q input168/X _08365_/X VGND VGND VPWR VPWR _08366_/X
+ sky130_fd_sc_hd__a221o_1
X_05578_ _05578_/A VGND VGND VPWR VPWR _05579_/A sky130_fd_sc_hd__inv_2
X_07317_ _07317_/A _07317_/B _07317_/C _07317_/D VGND VGND VPWR VPWR _07324_/C sky130_fd_sc_hd__or4_1
X_08297_ _07097_/Y _08184_/A _07086_/Y _08158_/A VGND VGND VPWR VPWR _08297_/X sky130_fd_sc_hd__o22a_1
XFILLER_191_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07248_ _07246_/Y _06251_/B _07247_/Y _05575_/A VGND VGND VPWR VPWR _07248_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ input22/X _06704_/A _07178_/Y _05177_/A VGND VGND VPWR VPWR _07179_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10190_ _10224_/CLK _10190_/D repeater410/X VGND VGND VPWR VPWR _10190_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_2
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_6
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_4
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10457_ _10486_/CLK _10457_/D repeater409/X VGND VGND VPWR VPWR _10457_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_184_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10388_ _10500_/CLK _10388_/D repeater407/X VGND VGND VPWR VPWR _10388_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04880_ _05806_/A VGND VGND VPWR VPWR _04993_/A sky130_fd_sc_hd__buf_4
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06550_ _06550_/A VGND VGND VPWR VPWR _06551_/B sky130_fd_sc_hd__clkbuf_4
X_05501_ _06646_/A VGND VGND VPWR VPWR _05518_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06481_ _06481_/A _06481_/B VGND VGND VPWR VPWR _06483_/A sky130_fd_sc_hd__or2_2
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08220_ _08220_/A VGND VGND VPWR VPWR _08220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05432_ _05806_/A VGND VGND VPWR VPWR _05603_/A sky130_fd_sc_hd__buf_4
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08151_ _07010_/Y _08092_/X _07738_/A _08093_/X _08150_/X VGND VGND VPWR VPWR _08152_/D
+ sky130_fd_sc_hd__o221a_1
X_05363_ _05354_/Y _06312_/A _05356_/Y _05527_/A _05362_/X VGND VGND VPWR VPWR _05364_/D
+ sky130_fd_sc_hd__o221a_1
X_05294_ _10193_/Q VGND VGND VPWR VPWR _05294_/Y sky130_fd_sc_hd__clkinv_4
X_08082_ _08201_/A VGND VGND VPWR VPWR _08082_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07102_ _10188_/Q VGND VGND VPWR VPWR _09513_/A sky130_fd_sc_hd__inv_6
XFILLER_161_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07033_ _10126_/Q _05073_/Y _10475_/Q _06776_/A _07032_/X VGND VGND VPWR VPWR _07040_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08984_ _09297_/B _09433_/A _08984_/C VGND VGND VPWR VPWR _08985_/B sky130_fd_sc_hd__or3_1
XFILLER_142_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07935_ _07228_/Y _07825_/X _07178_/Y _07827_/X _07934_/X VGND VGND VPWR VPWR _07936_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07866_ _05360_/Y _07787_/X _05276_/Y _07788_/X _07865_/X VGND VGND VPWR VPWR _07875_/A
+ sky130_fd_sc_hd__o221a_1
X_09605_ _09604_/X _09914_/Q _09776_/Q VGND VGND VPWR VPWR _09605_/X sky130_fd_sc_hd__mux2_1
X_06817_ _10095_/Q VGND VGND VPWR VPWR _06817_/Y sky130_fd_sc_hd__inv_2
X_07797_ _06821_/Y _07792_/X _06799_/Y _07793_/X _07796_/X VGND VGND VPWR VPWR _07810_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06748_ _09954_/Q VGND VGND VPWR VPWR _06748_/Y sky130_fd_sc_hd__inv_2
X_09536_ _09678_/X _04822_/Y _09536_/A3 _10513_/Q _04827_/X VGND VGND VPWR VPWR _10513_/D
+ sky130_fd_sc_hd__a32o_1
X_09467_ _09467_/A VGND VGND VPWR VPWR _09468_/A sky130_fd_sc_hd__clkbuf_1
X_08418_ _08634_/B VGND VGND VPWR VPWR _08640_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06679_ _06679_/A _06679_/B _06679_/C VGND VGND VPWR VPWR _06680_/A sky130_fd_sc_hd__or3_1
X_09398_ _09398_/A _09398_/B _09398_/C _09398_/D VGND VGND VPWR VPWR _09421_/D sky130_fd_sc_hd__or4_2
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08349_ _09813_/Q VGND VGND VPWR VPWR _08349_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10311_ _10504_/CLK _10311_/D repeater404/X VGND VGND VPWR VPWR _10311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10242_ _10244_/CLK _10242_/D repeater402/X VGND VGND VPWR VPWR _10242_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10173_ _10491_/CLK _10173_/D repeater403/X VGND VGND VPWR VPWR _10173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10509_ _10512_/CLK _10509_/D _07492_/B VGND VGND VPWR VPWR _10509_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater403 repeater404/X VGND VGND VPWR VPWR repeater403/X sky130_fd_sc_hd__buf_12
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07720_ _06980_/Y _07620_/X _07718_/Y _07621_/X _07719_/X VGND VGND VPWR VPWR _07720_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05981_ _05982_/A VGND VGND VPWR VPWR _05981_/X sky130_fd_sc_hd__clkbuf_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04932_ _05340_/A VGND VGND VPWR VPWR _05261_/B sky130_fd_sc_hd__clkbuf_8
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_07651_ _07811_/A VGND VGND VPWR VPWR _07651_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04863_ _09663_/X _05201_/C _05135_/C VGND VGND VPWR VPWR _05318_/B sky130_fd_sc_hd__or3_4
X_07582_ _07608_/A _07582_/B VGND VGND VPWR VPWR _07792_/A sky130_fd_sc_hd__or2_4
X_06602_ _09772_/Q _06602_/B _07489_/B VGND VGND VPWR VPWR _06602_/X sky130_fd_sc_hd__and3_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06533_ _09831_/Q _06530_/X _09577_/X _06531_/Y VGND VGND VPWR VPWR _09831_/D sky130_fd_sc_hd__a22o_1
X_09321_ _09321_/A VGND VGND VPWR VPWR _09378_/C sky130_fd_sc_hd__inv_2
XFILLER_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06464_ _08492_/A _08378_/A VGND VGND VPWR VPWR _06464_/X sky130_fd_sc_hd__or2_1
X_09252_ _09252_/A VGND VGND VPWR VPWR _09252_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06395_ _06395_/A VGND VGND VPWR VPWR _06395_/Y sky130_fd_sc_hd__inv_2
X_05415_ hold44/A _05397_/A hold48/A _05398_/A VGND VGND VPWR VPWR _10413_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09183_ _09415_/C _09329_/A _09183_/C VGND VGND VPWR VPWR _09185_/A sky130_fd_sc_hd__or3_1
X_08203_ _06816_/Y _08201_/X _06798_/Y _08202_/X VGND VGND VPWR VPWR _08203_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08134_ _08134_/A _08134_/B _08134_/C _08134_/D VGND VGND VPWR VPWR _08135_/D sky130_fd_sc_hd__and4_2
X_05346_ _05346_/A _05361_/B VGND VGND VPWR VPWR _05347_/A sky130_fd_sc_hd__or2_1
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05277_ _05277_/A VGND VGND VPWR VPWR _05359_/B sky130_fd_sc_hd__clkbuf_2
X_08065_ _08184_/A VGND VGND VPWR VPWR _08065_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07016_ _10402_/Q VGND VGND VPWR VPWR _07016_/Y sky130_fd_sc_hd__clkinv_4
X_08967_ _08967_/A _09291_/B VGND VGND VPWR VPWR _08969_/A sky130_fd_sc_hd__or2_1
XFILLER_76_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08898_ _08898_/A VGND VGND VPWR VPWR _09184_/B sky130_fd_sc_hd__inv_2
X_07918_ _07185_/Y _07787_/X _07222_/Y _07788_/X _07917_/X VGND VGND VPWR VPWR _07926_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07849_ _06724_/Y _07812_/X _06742_/Y _07813_/X VGND VGND VPWR VPWR _07849_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09519_ _09519_/A VGND VGND VPWR VPWR _09520_/A sky130_fd_sc_hd__clkbuf_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10225_ _10349_/CLK _10225_/D repeater405/X VGND VGND VPWR VPWR _10225_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10156_ _10354_/CLK _10156_/D repeater406/X VGND VGND VPWR VPWR _10156_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_94_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10087_ _10374_/CLK _10087_/D hold41/X VGND VGND VPWR VPWR _10087_/Q sky130_fd_sc_hd__dfrtp_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05200_ _09894_/Q VGND VGND VPWR VPWR _05200_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06180_ _08027_/A VGND VGND VPWR VPWR _08038_/A sky130_fd_sc_hd__clkbuf_2
X_05131_ input4/X _05129_/X _10443_/Q _06688_/A VGND VGND VPWR VPWR _05131_/X sky130_fd_sc_hd__a22o_2
X_05062_ _05062_/A VGND VGND VPWR VPWR _05062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09870_ _10350_/CLK _09870_/D repeater404/X VGND VGND VPWR VPWR _09870_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _09060_/A _08821_/B _09283_/A _09395_/B VGND VGND VPWR VPWR _08825_/A sky130_fd_sc_hd__or4_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08752_ _08752_/A VGND VGND VPWR VPWR _09226_/A sky130_fd_sc_hd__clkinv_4
X_05964_ _10126_/Q _05961_/X _09658_/A1 _05962_/Y VGND VGND VPWR VPWR _10126_/D sky130_fd_sc_hd__a22o_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ _08683_/A VGND VGND VPWR VPWR _09048_/A sky130_fd_sc_hd__buf_2
X_07703_ _09515_/A _07568_/B _09479_/A _07642_/X VGND VGND VPWR VPWR _07703_/X sky130_fd_sc_hd__o22a_4
X_04915_ _04915_/A VGND VGND VPWR VPWR _04915_/Y sky130_fd_sc_hd__inv_2
X_05895_ _05895_/A VGND VGND VPWR VPWR _05896_/B sky130_fd_sc_hd__buf_2
X_07634_ _07794_/A VGND VGND VPWR VPWR _07634_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04846_ _10373_/Q _09798_/Q input67/X VGND VGND VPWR VPWR _04847_/A sky130_fd_sc_hd__or3_4
XFILLER_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07565_ _07565_/A _07608_/B VGND VGND VPWR VPWR _07573_/A sky130_fd_sc_hd__or2_1
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09304_ _09304_/A VGND VGND VPWR VPWR _09353_/A sky130_fd_sc_hd__inv_2
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07496_ _10297_/Q input88/X VGND VGND VPWR VPWR _07497_/A sky130_fd_sc_hd__or2_1
X_06516_ _06538_/A _06516_/B VGND VGND VPWR VPWR _06518_/A sky130_fd_sc_hd__or2_2
X_09235_ _09324_/B _09235_/B _09235_/C _09378_/A VGND VGND VPWR VPWR _09240_/B sky130_fd_sc_hd__or4_2
X_06447_ _09871_/Q _06440_/X _09550_/A0 _06442_/X VGND VGND VPWR VPWR _09871_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06378_ _06374_/X _09607_/X _09650_/X _09916_/Q VGND VGND VPWR VPWR _09916_/D sky130_fd_sc_hd__o22a_1
X_09166_ _09010_/X _09024_/A _08466_/A _09260_/A VGND VGND VPWR VPWR _09326_/C sky130_fd_sc_hd__o22ai_2
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09097_ _09253_/C VGND VGND VPWR VPWR _09098_/A sky130_fd_sc_hd__inv_2
X_05329_ _05329_/A _05361_/B VGND VGND VPWR VPWR _06480_/A sky130_fd_sc_hd__or2_4
X_08117_ _08117_/A _08117_/B _08117_/C _08117_/D VGND VGND VPWR VPWR _08117_/Y sky130_fd_sc_hd__nand4_4
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08048_ _05335_/Y _08211_/A _07606_/A _08212_/A _08047_/X VGND VGND VPWR VPWR _08049_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ _10500_/CLK _10010_/D repeater407/X VGND VGND VPWR VPWR _10010_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09999_ _10364_/CLK _09999_/D repeater410/X VGND VGND VPWR VPWR _09999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _10486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10208_ _10354_/CLK _10208_/D repeater406/X VGND VGND VPWR VPWR _10208_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10139_ _10371_/CLK _10139_/D repeater410/X VGND VGND VPWR VPWR _10139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05680_ _05680_/A VGND VGND VPWR VPWR _05680_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07350_ _09869_/Q VGND VGND VPWR VPWR _07350_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06301_ _09961_/Q _06293_/A _09661_/A1 _06294_/A VGND VGND VPWR VPWR _09961_/D sky130_fd_sc_hd__a22o_1
XFILLER_176_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07281_ _09976_/Q VGND VGND VPWR VPWR _07690_/A sky130_fd_sc_hd__inv_2
X_09020_ _09020_/A _09023_/A VGND VGND VPWR VPWR _09198_/C sky130_fd_sc_hd__nor2_1
XFILLER_148_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06232_ _06232_/A VGND VGND VPWR VPWR _06232_/X sky130_fd_sc_hd__buf_2
X_06163_ _10014_/Q _06156_/A _09660_/A1 _06157_/A VGND VGND VPWR VPWR _10014_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_18_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10289_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05114_ _05114_/A VGND VGND VPWR VPWR _05114_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_144_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06094_ _10045_/Q _06088_/X _09536_/A3 _06089_/Y VGND VGND VPWR VPWR _10045_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09922_ _10000_/CLK _09922_/D repeater405/X VGND VGND VPWR VPWR _09922_/Q sky130_fd_sc_hd__dfrtp_1
X_05045_ _05045_/A VGND VGND VPWR VPWR _05045_/X sky130_fd_sc_hd__clkbuf_1
X_09853_ _10288_/CLK _09853_/D repeater406/X VGND VGND VPWR VPWR _09853_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _10382_/CLK _09784_/D _06658_/X VGND VGND VPWR VPWR _09784_/Q sky130_fd_sc_hd__dfrtp_1
X_08804_ _08804_/A VGND VGND VPWR VPWR _09096_/B sky130_fd_sc_hd__buf_4
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _10106_/Q VGND VGND VPWR VPWR _06996_/Y sky130_fd_sc_hd__clkinv_4
X_08735_ _08787_/B _09265_/A _08734_/Y VGND VGND VPWR VPWR _08739_/A sky130_fd_sc_hd__o21ba_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05947_ _10137_/Q _05941_/X _09545_/A1 _05943_/X VGND VGND VPWR VPWR _10137_/D sky130_fd_sc_hd__a22o_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05878_ _10178_/Q _05875_/X _09577_/X _05876_/Y VGND VGND VPWR VPWR _10178_/D sky130_fd_sc_hd__a22o_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08841_/B VGND VGND VPWR VPWR _09262_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_119 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _08504_/B _08883_/A _08596_/Y VGND VGND VPWR VPWR _08598_/B sky130_fd_sc_hd__o21ba_1
X_07617_ _07617_/A VGND VGND VPWR VPWR _07617_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04829_ _05155_/A VGND VGND VPWR VPWR _05149_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07548_ _07799_/A VGND VGND VPWR VPWR _07639_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07479_ _07479_/A VGND VGND VPWR VPWR _07479_/Y sky130_fd_sc_hd__inv_2
X_09218_ _09218_/A _09372_/B _09372_/C VGND VGND VPWR VPWR _09315_/C sky130_fd_sc_hd__nor3_1
X_10490_ _10490_/CLK _10490_/D repeater404/X VGND VGND VPWR VPWR _10490_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09149_ _09149_/A _09149_/B VGND VGND VPWR VPWR _09157_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput307 _10443_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_2
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 _10449_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_2
Xoutput318 _10444_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_2
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06850_ _10060_/Q _05162_/X _10112_/Q _05094_/Y _06849_/X VGND VGND VPWR VPWR _06855_/C
+ sky130_fd_sc_hd__a221o_1
X_05801_ _10223_/Q _05795_/X _09547_/A1 _05797_/X VGND VGND VPWR VPWR _10223_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06781_ _06779_/Y _05980_/B _06780_/X VGND VGND VPWR VPWR _06781_/Y sky130_fd_sc_hd__o21ai_2
X_05732_ _10265_/Q _05729_/X _09581_/X _05731_/X VGND VGND VPWR VPWR _10265_/D sky130_fd_sc_hd__a22o_1
X_08520_ _08752_/A _08520_/B VGND VGND VPWR VPWR _09311_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05663_ _10300_/Q _05654_/A _09574_/X _05655_/A VGND VGND VPWR VPWR _10300_/D sky130_fd_sc_hd__a22o_1
X_08451_ _08687_/A _08701_/A VGND VGND VPWR VPWR _08812_/A sky130_fd_sc_hd__or2_2
XFILLER_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07402_ _10176_/Q VGND VGND VPWR VPWR _07402_/Y sky130_fd_sc_hd__inv_2
X_08382_ _09233_/A _08561_/B _08571_/C _09236_/A VGND VGND VPWR VPWR _08687_/A sky130_fd_sc_hd__or4_2
XFILLER_149_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05594_ _09771_/Q _05590_/Y _06593_/B _10342_/Q VGND VGND VPWR VPWR _10342_/D sky130_fd_sc_hd__a31o_1
X_07333_ _09942_/Q VGND VGND VPWR VPWR _07333_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07264_ _10039_/Q VGND VGND VPWR VPWR _07264_/Y sky130_fd_sc_hd__clkinv_4
X_09003_ _09003_/A VGND VGND VPWR VPWR _09159_/A sky130_fd_sc_hd__inv_2
X_06215_ _09996_/Q _06208_/A _09660_/A1 _06209_/A VGND VGND VPWR VPWR _09996_/D sky130_fd_sc_hd__a22o_1
X_07195_ _10359_/Q VGND VGND VPWR VPWR _07195_/Y sky130_fd_sc_hd__clkinv_4
X_06146_ _06140_/B _06137_/X _06150_/A _06145_/X VGND VGND VPWR VPWR _10022_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06077_ _10055_/Q _06068_/A _09536_/A3 _06069_/A VGND VGND VPWR VPWR _10055_/D sky130_fd_sc_hd__a22o_1
X_09905_ _10119_/CLK _09905_/D repeater403/X VGND VGND VPWR VPWR _09905_/Q sky130_fd_sc_hd__dfrtp_1
X_05028_ _05100_/B VGND VGND VPWR VPWR _05355_/A sky130_fd_sc_hd__buf_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _10364_/CLK _09836_/D repeater410/X VGND VGND VPWR VPWR _09836_/Q sky130_fd_sc_hd__dfrtp_2
X_06979_ _09872_/Q VGND VGND VPWR VPWR _06979_/Y sky130_fd_sc_hd__inv_2
X_09767_ _10471_/CLK _09767_/D VGND VGND VPWR VPWR _09767_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09454_/X _09440_/X _09698_/S VGND VGND VPWR VPWR _09698_/X sky130_fd_sc_hd__mux2_1
X_08718_ _08736_/A _09262_/A VGND VGND VPWR VPWR _09326_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _09085_/B _08783_/A VGND VGND VPWR VPWR _08650_/A sky130_fd_sc_hd__or2_2
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10473_ _10478_/CLK _10473_/D _05034_/A VGND VGND VPWR VPWR _10473_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_19 _06967_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06000_ _10102_/Q _05994_/X _09574_/X _05995_/Y VGND VGND VPWR VPWR _10102_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07951_ _07951_/A _07951_/B _07951_/C _07951_/D VGND VGND VPWR VPWR _07962_/B sky130_fd_sc_hd__and4_1
X_06902_ _06897_/Y _05762_/B _06898_/Y _05839_/B _06901_/X VGND VGND VPWR VPWR _06902_/X
+ sky130_fd_sc_hd__o221a_2
X_07882_ _05317_/Y _07768_/X _05244_/Y _07769_/X _07881_/X VGND VGND VPWR VPWR _07885_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06833_ _06833_/A _06833_/B _06833_/C VGND VGND VPWR VPWR _06833_/X sky130_fd_sc_hd__and3_2
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09621_ _09620_/X _09884_/Q _09776_/Q VGND VGND VPWR VPWR _09621_/X sky130_fd_sc_hd__mux2_1
X_09552_ _09578_/X _10304_/Q _09677_/S VGND VGND VPWR VPWR _09552_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06764_ _06764_/A VGND VGND VPWR VPWR _06764_/X sky130_fd_sc_hd__clkbuf_2
X_08503_ _08512_/A VGND VGND VPWR VPWR _08504_/B sky130_fd_sc_hd__buf_2
XFILLER_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05715_ _09699_/X _05715_/B VGND VGND VPWR VPWR _05718_/A sky130_fd_sc_hd__or2_4
X_09483_ _09483_/A VGND VGND VPWR VPWR _09484_/A sky130_fd_sc_hd__clkbuf_1
X_06695_ _10088_/Q _06692_/Y input70/X _09679_/S _06694_/X VGND VGND VPWR VPWR _06701_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08434_ _08476_/A _08476_/B _09247_/B VGND VGND VPWR VPWR _09224_/B sky130_fd_sc_hd__o21ai_2
X_05646_ _10312_/Q _05640_/X _09547_/A1 _05642_/X VGND VGND VPWR VPWR _10312_/D sky130_fd_sc_hd__a22o_1
X_08365_ _09788_/Q _08365_/B VGND VGND VPWR VPWR _08365_/X sky130_fd_sc_hd__and2_1
X_05577_ _05578_/A VGND VGND VPWR VPWR _05577_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07316_ input44/X _06697_/X _10444_/Q _06688_/A _07315_/X VGND VGND VPWR VPWR _07317_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08296_ _07121_/Y _08177_/A _07126_/Y _08178_/A _08295_/X VGND VGND VPWR VPWR _08310_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ _10345_/Q VGND VGND VPWR VPWR _07247_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07178_ _10073_/Q VGND VGND VPWR VPWR _07178_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_132_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06129_ _10024_/Q _06123_/X _09536_/A3 _06124_/Y VGND VGND VPWR VPWR _10024_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09819_ _10354_/CLK _09819_/D repeater406/X VGND VGND VPWR VPWR _09819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_2
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_2
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__buf_6
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10456_ _10486_/CLK _10456_/D repeater409/X VGND VGND VPWR VPWR _10456_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10387_ _10500_/CLK _10387_/D repeater407/X VGND VGND VPWR VPWR _10387_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05500_ _05500_/A VGND VGND VPWR VPWR _10384_/D sky130_fd_sc_hd__clkbuf_1
X_06480_ _06480_/A VGND VGND VPWR VPWR _06481_/B sky130_fd_sc_hd__buf_2
X_05431_ _10420_/Q _05430_/Y _10406_/Q _05430_/A VGND VGND VPWR VPWR _10406_/D sky130_fd_sc_hd__a22o_1
X_08150_ _06981_/Y _08094_/X _06932_/Y _08095_/X VGND VGND VPWR VPWR _08150_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07101_ _09511_/A _05807_/A _07097_/Y _05830_/B _07100_/X VGND VGND VPWR VPWR _07114_/B
+ sky130_fd_sc_hd__o221a_1
X_05362_ _05358_/Y _06528_/A _05360_/Y _06471_/A VGND VGND VPWR VPWR _05362_/X sky130_fd_sc_hd__o22a_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05293_ _05293_/A VGND VGND VPWR VPWR _05952_/B sky130_fd_sc_hd__buf_2
X_08081_ _08200_/A VGND VGND VPWR VPWR _08081_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07032_ _10327_/Q _05156_/Y _10340_/Q _05126_/Y VGND VGND VPWR VPWR _07032_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _10023_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08983_ _09184_/B _08983_/B VGND VGND VPWR VPWR _08984_/C sky130_fd_sc_hd__or2_1
X_07934_ _07266_/Y _07828_/X _07213_/Y _07829_/X VGND VGND VPWR VPWR _07934_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07865_ _05332_/Y _07749_/X _05358_/Y _07789_/X VGND VGND VPWR VPWR _07865_/X sky130_fd_sc_hd__o22a_1
X_09604_ _08256_/Y _10324_/Q _09700_/S VGND VGND VPWR VPWR _09604_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07796_ _06805_/Y _07794_/X _06803_/Y _07795_/X VGND VGND VPWR VPWR _07796_/X sky130_fd_sc_hd__o22a_1
X_06816_ _10018_/Q VGND VGND VPWR VPWR _06816_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09535_ _09535_/A _09535_/B VGND VGND VPWR VPWR _09782_/D sky130_fd_sc_hd__nor2_1
X_06747_ _09875_/Q VGND VGND VPWR VPWR _06747_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09466_ _09466_/A VGND VGND VPWR VPWR _09466_/X sky130_fd_sc_hd__clkbuf_1
X_06678_ _06678_/A VGND VGND VPWR VPWR _06678_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08417_ _08417_/A VGND VGND VPWR VPWR _08634_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05629_ _05629_/A VGND VGND VPWR VPWR _05629_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09397_ _09397_/A _09397_/B VGND VGND VPWR VPWR _09398_/B sky130_fd_sc_hd__or2_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08348_ _09812_/Q VGND VGND VPWR VPWR _08348_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08279_ _07271_/Y _08184_/X _07246_/Y _08158_/A VGND VGND VPWR VPWR _08279_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10310_ _10310_/CLK _10310_/D repeater404/X VGND VGND VPWR VPWR _10310_/Q sky130_fd_sc_hd__dfrtp_1
X_10241_ _10244_/CLK _10241_/D repeater402/X VGND VGND VPWR VPWR _10241_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10172_ _10491_/CLK _10172_/D repeater403/X VGND VGND VPWR VPWR _10172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10508_ _10508_/CLK _10508_/D repeater402/X VGND VGND VPWR VPWR _10508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10439_ _10478_/CLK _10439_/D repeater409/X VGND VGND VPWR VPWR _10439_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05980_ _06011_/A _05980_/B VGND VGND VPWR VPWR _05982_/A sky130_fd_sc_hd__or2_2
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater404 repeater405/X VGND VGND VPWR VPWR repeater404/X sky130_fd_sc_hd__buf_12
XFILLER_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04931_ _09670_/X _05109_/D _05082_/A _09676_/X VGND VGND VPWR VPWR _05340_/A sky130_fd_sc_hd__or4_4
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07650_ _07650_/A _07650_/B _07650_/C _07650_/D VGND VGND VPWR VPWR _07672_/B sky130_fd_sc_hd__and4_1
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04862_ _06630_/C VGND VGND VPWR VPWR _05541_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07581_ _05225_/Y _07627_/A _05248_/Y _07788_/A _07580_/X VGND VGND VPWR VPWR _07595_/A
+ sky130_fd_sc_hd__o221a_1
X_06601_ _09812_/Q _06601_/B VGND VGND VPWR VPWR _07489_/B sky130_fd_sc_hd__nand2_1
X_06532_ _09832_/Q _06530_/X _09547_/A1 _06531_/Y VGND VGND VPWR VPWR _09832_/D sky130_fd_sc_hd__a22o_1
X_09320_ _09204_/A _08620_/A _09006_/B _08704_/C _09155_/X VGND VGND VPWR VPWR _09321_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09251_ _09415_/B _09317_/A _09417_/A _09250_/Y VGND VGND VPWR VPWR _09252_/A sky130_fd_sc_hd__or4b_1
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06463_ _08492_/B VGND VGND VPWR VPWR _08378_/A sky130_fd_sc_hd__inv_2
X_08202_ _08202_/A VGND VGND VPWR VPWR _08202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06394_ _06395_/A VGND VGND VPWR VPWR _06394_/X sky130_fd_sc_hd__clkbuf_2
X_05414_ _05414_/A VGND VGND VPWR VPWR _05414_/X sky130_fd_sc_hd__clkbuf_1
X_09182_ _09182_/A _09182_/B VGND VGND VPWR VPWR _09183_/C sky130_fd_sc_hd__or2_1
XFILLER_146_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05345_ _10407_/Q VGND VGND VPWR VPWR _05345_/Y sky130_fd_sc_hd__inv_2
X_08133_ _09465_/A _08092_/X _09481_/A _08093_/X _08132_/X VGND VGND VPWR VPWR _08134_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08064_ _08183_/A VGND VGND VPWR VPWR _08064_/X sky130_fd_sc_hd__clkbuf_2
X_07015_ _09906_/Q VGND VGND VPWR VPWR _07015_/Y sky130_fd_sc_hd__clkinv_4
X_05276_ _09815_/Q VGND VGND VPWR VPWR _05276_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08966_ _09372_/A _08968_/B VGND VGND VPWR VPWR _09291_/B sky130_fd_sc_hd__nor2_1
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08897_ _08897_/A _08897_/B VGND VGND VPWR VPWR _09433_/A sky130_fd_sc_hd__nor2_2
X_07917_ _07239_/Y _07527_/A _07234_/Y _07789_/X VGND VGND VPWR VPWR _07917_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07848_ _07848_/A _07848_/B _07848_/C _07848_/D VGND VGND VPWR VPWR _07860_/B sky130_fd_sc_hd__and4_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09518_ _09518_/A VGND VGND VPWR VPWR _09518_/X sky130_fd_sc_hd__clkbuf_1
X_07779_ _07779_/A VGND VGND VPWR VPWR _07779_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _08674_/X _09265_/B _09448_/X _09340_/X VGND VGND VPWR VPWR _09449_/Y sky130_fd_sc_hd__o211ai_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10224_ _10224_/CLK _10224_/D repeater405/X VGND VGND VPWR VPWR _10224_/Q sky130_fd_sc_hd__dfrtp_1
X_10155_ _10157_/CLK _10155_/D repeater406/X VGND VGND VPWR VPWR _10155_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10086_ _10374_/CLK _10086_/D repeater410/X VGND VGND VPWR VPWR _10086_/Q sky130_fd_sc_hd__dfrtp_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05130_ _05130_/A VGND VGND VPWR VPWR _06688_/A sky130_fd_sc_hd__inv_2
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05061_ _05378_/A VGND VGND VPWR VPWR _05062_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08837_/A _08823_/A VGND VGND VPWR VPWR _09395_/B sky130_fd_sc_hd__nor2_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08751_ _08751_/A _08751_/B VGND VGND VPWR VPWR _08754_/A sky130_fd_sc_hd__or2_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05963_ _10127_/Q _05961_/X _09545_/A1 _05962_/Y VGND VGND VPWR VPWR _10127_/D sky130_fd_sc_hd__a22o_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05894_ _10167_/Q _05885_/A _09659_/A1 _05886_/A VGND VGND VPWR VPWR _10167_/D sky130_fd_sc_hd__a22o_1
X_08682_ _08809_/B _08737_/B VGND VGND VPWR VPWR _08683_/A sky130_fd_sc_hd__or2_1
X_07702_ _09495_/A _07632_/X _09475_/A _07633_/X _07701_/X VGND VGND VPWR VPWR _07707_/B
+ sky130_fd_sc_hd__o221a_2
X_04914_ _05286_/A _06780_/A VGND VGND VPWR VPWR _04915_/A sky130_fd_sc_hd__or2_1
X_07633_ _07793_/A VGND VGND VPWR VPWR _07633_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04845_ _04845_/A VGND VGND VPWR VPWR _05677_/B sky130_fd_sc_hd__buf_8
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07564_ _07585_/C _07612_/A _07564_/C VGND VGND VPWR VPWR _07572_/A sky130_fd_sc_hd__or3_1
XFILLER_34_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09303_ _09218_/A _09206_/A _08546_/B _09105_/A VGND VGND VPWR VPWR _09303_/Y sky130_fd_sc_hd__o211ai_1
X_06515_ _06515_/A VGND VGND VPWR VPWR _06516_/B sky130_fd_sc_hd__buf_4
X_07495_ _07495_/A VGND VGND VPWR VPWR _07495_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09234_ _09233_/Y _09225_/Y _09237_/A _09157_/A VGND VGND VPWR VPWR _09378_/A sky130_fd_sc_hd__a31o_1
X_06446_ _09872_/Q _06440_/X _09547_/A1 _06442_/X VGND VGND VPWR VPWR _09872_/D sky130_fd_sc_hd__a22o_1
X_09165_ _08746_/A _08581_/B _08714_/X VGND VGND VPWR VPWR _09167_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08116_ _08116_/A _08116_/B _08116_/C _08116_/D VGND VGND VPWR VPWR _08117_/D sky130_fd_sc_hd__and4_2
X_06377_ _06374_/X _09609_/X _09650_/X _09917_/Q VGND VGND VPWR VPWR _09917_/D sky130_fd_sc_hd__o22a_1
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05328_ _09854_/Q VGND VGND VPWR VPWR _05328_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09096_ _09226_/B _09096_/B VGND VGND VPWR VPWR _09253_/C sky130_fd_sc_hd__or2_1
X_05259_ _05248_/Y _06537_/A _05251_/Y _05918_/B _05258_/X VGND VGND VPWR VPWR _05281_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08047_ _05197_/Y _08213_/A _05274_/Y _08214_/A VGND VGND VPWR VPWR _08047_/X sky130_fd_sc_hd__o22a_1
XFILLER_122_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09998_ _10000_/CLK _09998_/D repeater410/X VGND VGND VPWR VPWR _09998_/Q sky130_fd_sc_hd__dfrtp_1
X_08949_ _09024_/A _08957_/B VGND VGND VPWR VPWR _09289_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10207_ _10409_/CLK _10207_/D repeater406/X VGND VGND VPWR VPWR _10207_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10138_ _10374_/CLK _10138_/D _07492_/B VGND VGND VPWR VPWR _10138_/Q sky130_fd_sc_hd__dfrtp_1
X_10069_ _10350_/CLK _10069_/D repeater405/X VGND VGND VPWR VPWR _10069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06300_ _09962_/Q _06293_/A _09660_/A1 _06294_/A VGND VGND VPWR VPWR _09962_/D sky130_fd_sc_hd__a22o_1
X_07280_ _07275_/Y _05918_/B _07276_/Y _05896_/B _07279_/X VGND VGND VPWR VPWR _07287_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06231_ _07768_/A VGND VGND VPWR VPWR _06232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06162_ _10015_/Q _06155_/X _09550_/A0 _06157_/X VGND VGND VPWR VPWR _10015_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_144_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06093_ _10046_/Q _06088_/X _06684_/B1 _06089_/Y VGND VGND VPWR VPWR _10046_/D sky130_fd_sc_hd__a22o_1
X_05113_ _05677_/B VGND VGND VPWR VPWR _05114_/A sky130_fd_sc_hd__inv_2
X_09921_ _10224_/CLK _09921_/D repeater405/X VGND VGND VPWR VPWR _09921_/Q sky130_fd_sc_hd__dfstp_1
X_05044_ _05053_/A VGND VGND VPWR VPWR _05045_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_171_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09852_ _10355_/CLK _09852_/D repeater406/X VGND VGND VPWR VPWR _09852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10382_/CLK _09783_/D _06660_/X VGND VGND VPWR VPWR _09783_/Q sky130_fd_sc_hd__dfrtp_1
X_08803_ _08822_/B VGND VGND VPWR VPWR _08804_/A sky130_fd_sc_hd__inv_2
XFILLER_98_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _06990_/Y _05567_/B _06991_/Y _05576_/B _06994_/X VGND VGND VPWR VPWR _06995_/X
+ sky130_fd_sc_hd__o221a_1
X_08734_ _09265_/A _08743_/A _08733_/X VGND VGND VPWR VPWR _08734_/Y sky130_fd_sc_hd__o21ai_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05946_ _10138_/Q _05941_/X _09579_/X _05943_/X VGND VGND VPWR VPWR _10138_/D sky130_fd_sc_hd__a22o_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05877_ _10179_/Q _05875_/X _09578_/X _05876_/Y VGND VGND VPWR VPWR _10179_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08665_ _08841_/B VGND VGND VPWR VPWR _08665_/Y sky130_fd_sc_hd__inv_2
XANTENNA_109 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08596_/A _08596_/B VGND VGND VPWR VPWR _08596_/Y sky130_fd_sc_hd__nand2_1
X_07616_ _07616_/A _07616_/B _07616_/C VGND VGND VPWR VPWR _07617_/A sky130_fd_sc_hd__and3_1
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04828_ _09678_/X _04822_/Y _06683_/B1 _10512_/Q _04827_/X VGND VGND VPWR VPWR _10512_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07547_ _07565_/A _07574_/B VGND VGND VPWR VPWR _07799_/A sky130_fd_sc_hd__or2_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07478_ _07470_/Y _06176_/A _07476_/Y _07479_/A VGND VGND VPWR VPWR _09777_/D sky130_fd_sc_hd__o22ai_1
X_09217_ _09217_/A _09405_/A _09312_/B _09374_/B VGND VGND VPWR VPWR _09220_/B sky130_fd_sc_hd__or4_1
X_06429_ _06429_/A VGND VGND VPWR VPWR _06430_/B sky130_fd_sc_hd__clkbuf_4
X_09148_ _09010_/X _08925_/A _08662_/A _08808_/X VGND VGND VPWR VPWR _09377_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09079_ _09079_/A _09405_/B VGND VGND VPWR VPWR _09294_/A sky130_fd_sc_hd__or2_2
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput308 _10453_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_2
XFILLER_99_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput319 _10463_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_2
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05800_ _10224_/Q _05795_/X _09579_/X _05797_/X VGND VGND VPWR VPWR _10224_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06780_ _06780_/A _06780_/B VGND VGND VPWR VPWR _06780_/X sky130_fd_sc_hd__or2_2
XFILLER_55_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05731_ _05731_/A VGND VGND VPWR VPWR _05731_/X sky130_fd_sc_hd__clkbuf_2
X_05662_ _10301_/Q _05654_/A hold46/X _05655_/A VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__a22o_1
X_08450_ _08494_/A _09344_/A VGND VGND VPWR VPWR _08701_/A sky130_fd_sc_hd__or2_1
X_07401_ _09816_/Q VGND VGND VPWR VPWR _07401_/Y sky130_fd_sc_hd__clkinv_2
X_08381_ _08980_/C VGND VGND VPWR VPWR _08385_/B sky130_fd_sc_hd__clkbuf_2
X_07332_ _10202_/Q VGND VGND VPWR VPWR _07332_/Y sky130_fd_sc_hd__inv_2
X_05593_ _06589_/B VGND VGND VPWR VPWR _06593_/B sky130_fd_sc_hd__clkinv_2
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07263_ _09856_/Q VGND VGND VPWR VPWR _07263_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07194_ _09878_/Q VGND VGND VPWR VPWR _07194_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09002_ _09023_/A VGND VGND VPWR VPWR _09002_/Y sky130_fd_sc_hd__inv_2
X_06214_ _09997_/Q _06207_/X _09550_/A0 _06209_/X VGND VGND VPWR VPWR _09997_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06145_ _06140_/B _06260_/C _06137_/A _06142_/B VGND VGND VPWR VPWR _06145_/X sky130_fd_sc_hd__o31a_1
X_06076_ _10056_/Q _06068_/A _06684_/B1 _06069_/A VGND VGND VPWR VPWR _10056_/D sky130_fd_sc_hd__a22o_1
X_09904_ _10119_/CLK _09904_/D repeater403/X VGND VGND VPWR VPWR _09904_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05027_ _05027_/A _09668_/X _09674_/X _09676_/X VGND VGND VPWR VPWR _05100_/B sky130_fd_sc_hd__or4_2
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09835_ _10191_/CLK _09835_/D repeater410/X VGND VGND VPWR VPWR _09835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06978_ _06973_/Y _06480_/A _06974_/Y _06472_/B _06977_/X VGND VGND VPWR VPWR _06985_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09766_ _10471_/CLK _09766_/D VGND VGND VPWR VPWR _09766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05929_ _05930_/A VGND VGND VPWR VPWR _05929_/X sky130_fd_sc_hd__clkbuf_2
X_09697_ _09437_/Y _09409_/X _09698_/S VGND VGND VPWR VPWR _09697_/X sky130_fd_sc_hd__mux2_1
X_08717_ _08717_/A VGND VGND VPWR VPWR _08736_/A sky130_fd_sc_hd__buf_2
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _08855_/A VGND VGND VPWR VPWR _09265_/A sky130_fd_sc_hd__clkbuf_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _08934_/A _09010_/A _08576_/X _08577_/X _09162_/A VGND VGND VPWR VPWR _08579_/X
+ sky130_fd_sc_hd__o2111a_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10472_ _10478_/CLK _10472_/D _05034_/A VGND VGND VPWR VPWR _10472_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07950_ _07151_/Y _07645_/A _07948_/Y _07523_/A _07949_/X VGND VGND VPWR VPWR _07951_/D
+ sky130_fd_sc_hd__o221a_1
X_06901_ _06899_/Y _05727_/A _06900_/Y _05895_/A VGND VGND VPWR VPWR _06901_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07881_ _07881_/A _07932_/B VGND VGND VPWR VPWR _07881_/X sky130_fd_sc_hd__or2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06832_ _06827_/Y _05749_/B _06828_/Y _05839_/B _06831_/X VGND VGND VPWR VPWR _06833_/C
+ sky130_fd_sc_hd__o221a_1
X_09620_ _07744_/Y _10333_/Q _09682_/S VGND VGND VPWR VPWR _09620_/X sky130_fd_sc_hd__mux2_1
X_09551_ _09576_/X _10302_/Q _09677_/S VGND VGND VPWR VPWR _09551_/X sky130_fd_sc_hd__mux2_1
X_06763_ _06763_/A VGND VGND VPWR VPWR _06764_/A sky130_fd_sc_hd__inv_2
X_08502_ _09372_/B _09005_/A VGND VGND VPWR VPWR _08512_/A sky130_fd_sc_hd__or2_1
X_05714_ _05376_/X _05592_/B _10274_/Q _05713_/Y _05390_/X VGND VGND VPWR VPWR _10274_/D
+ sky130_fd_sc_hd__o221a_1
X_09482_ _09482_/A VGND VGND VPWR VPWR _09482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06694_ input33/X _05129_/X _10479_/Q _06776_/A VGND VGND VPWR VPWR _06694_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08433_ _08695_/B VGND VGND VPWR VPWR _09247_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05645_ _10313_/Q _05640_/X _09579_/X _05642_/X VGND VGND VPWR VPWR _10313_/D sky130_fd_sc_hd__a22o_1
X_08364_ _09790_/Q input184/X _09789_/Q input167/X _08363_/X VGND VGND VPWR VPWR _08364_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05576_ _05603_/A _05576_/B VGND VGND VPWR VPWR _05578_/A sky130_fd_sc_hd__or2_2
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07315_ input15/X _05129_/A _10030_/Q _05080_/A VGND VGND VPWR VPWR _07315_/X sky130_fd_sc_hd__a22o_1
X_08295_ _07128_/Y _08179_/A _07110_/Y _08180_/A VGND VGND VPWR VPWR _08295_/X sky130_fd_sc_hd__o22a_1
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07246_ _09985_/Q VGND VGND VPWR VPWR _07246_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07177_ _10083_/Q VGND VGND VPWR VPWR _07177_/Y sky130_fd_sc_hd__clkinv_4
X_06128_ _10025_/Q _06123_/X _06684_/B1 _06124_/Y VGND VGND VPWR VPWR _10025_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06059_ _10069_/Q _06055_/X _09580_/X _06057_/X VGND VGND VPWR VPWR _10069_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09818_ _10353_/CLK _09818_/D repeater403/X VGND VGND VPWR VPWR _09818_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09749_ _09752_/CLK _09749_/D VGND VGND VPWR VPWR _09749_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10455_ _10486_/CLK _10455_/D repeater409/X VGND VGND VPWR VPWR _10455_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10386_ _10500_/CLK _10386_/D repeater407/X VGND VGND VPWR VPWR _10386_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05430_ _05430_/A VGND VGND VPWR VPWR _05430_/Y sky130_fd_sc_hd__inv_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05361_ _06630_/B _05361_/B VGND VGND VPWR VPWR _06471_/A sky130_fd_sc_hd__or2_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07100_ _07098_/Y _05993_/B _09465_/A _06502_/A VGND VGND VPWR VPWR _07100_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05292_ _05292_/A _05316_/B VGND VGND VPWR VPWR _05293_/A sky130_fd_sc_hd__or2_1
X_08080_ _08199_/A VGND VGND VPWR VPWR _08080_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07031_ _06762_/X _07030_/X _09762_/Q _06764_/X VGND VGND VPWR VPWR _09762_/D sky130_fd_sc_hd__o22a_2
XFILLER_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08982_ _09248_/A _08982_/B VGND VGND VPWR VPWR _08983_/B sky130_fd_sc_hd__or2_1
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07933_ _07271_/Y _06232_/A _07284_/Y _07519_/A _07932_/X VGND VGND VPWR VPWR _07936_/C
+ sky130_fd_sc_hd__o221a_1
X_07864_ _05312_/Y _07777_/X _05186_/Y _07778_/X _07863_/X VGND VGND VPWR VPWR _07886_/A
+ sky130_fd_sc_hd__o221a_1
X_06815_ _10494_/Q VGND VGND VPWR VPWR _06815_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09603_ _09602_/X _09913_/Q _09776_/Q VGND VGND VPWR VPWR _09603_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07795_ _07795_/A VGND VGND VPWR VPWR _07795_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09534_ _09534_/A _09535_/B VGND VGND VPWR VPWR _09783_/D sky130_fd_sc_hd__nor2_1
X_06746_ _10070_/Q VGND VGND VPWR VPWR _06746_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09465_ _09465_/A VGND VGND VPWR VPWR _09466_/A sky130_fd_sc_hd__clkbuf_1
X_06677_ _06677_/A VGND VGND VPWR VPWR _06678_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08416_ _08564_/A _08565_/B VGND VGND VPWR VPWR _08774_/A sky130_fd_sc_hd__or2_1
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05628_ _05628_/A VGND VGND VPWR VPWR _05629_/A sky130_fd_sc_hd__inv_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09396_ _08808_/X _09337_/B _09113_/A _09395_/X _09341_/B VGND VGND VPWR VPWR _09401_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_165_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05559_ _10359_/Q _05552_/A _09660_/A1 _05553_/A VGND VGND VPWR VPWR _10359_/D sky130_fd_sc_hd__a22o_1
X_08347_ _09805_/Q _08344_/B _08346_/Y _09806_/Q _08344_/Y VGND VGND VPWR VPWR _08347_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08278_ _07253_/Y _08177_/X _07222_/Y _08178_/X _08277_/X VGND VGND VPWR VPWR _08292_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_180_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07229_ _07227_/Y _05927_/A _07228_/Y _06079_/B VGND VGND VPWR VPWR _07229_/X sky130_fd_sc_hd__o22a_1
X_10240_ _10290_/CLK _10240_/D repeater402/X VGND VGND VPWR VPWR _10240_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10171_ _10313_/CLK _10171_/D repeater403/X VGND VGND VPWR VPWR _10171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10507_ _10508_/CLK _10507_/D repeater402/X VGND VGND VPWR VPWR _10507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10438_ _10478_/CLK _10438_/D _05034_/A VGND VGND VPWR VPWR _10438_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_124_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10369_ _10369_/CLK _10369_/D repeater407/X VGND VGND VPWR VPWR _10369_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater405 _07492_/B VGND VGND VPWR VPWR repeater405/X sky130_fd_sc_hd__buf_12
X_04930_ _05149_/A VGND VGND VPWR VPWR _05118_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_04861_ _06679_/A VGND VGND VPWR VPWR _06630_/C sky130_fd_sc_hd__clkbuf_2
X_07580_ _05343_/Y _07527_/A _05212_/Y _07629_/A VGND VGND VPWR VPWR _07580_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06600_ _06600_/A VGND VGND VPWR VPWR _06600_/X sky130_fd_sc_hd__clkbuf_1
X_06531_ _06531_/A VGND VGND VPWR VPWR _06531_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09250_ _09250_/A _09329_/B _09417_/D _09331_/D VGND VGND VPWR VPWR _09250_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06462_ _08485_/A VGND VGND VPWR VPWR _08492_/A sky130_fd_sc_hd__inv_2
X_08201_ _08201_/A VGND VGND VPWR VPWR _08201_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05413_ _05588_/A VGND VGND VPWR VPWR _05414_/A sky130_fd_sc_hd__clkbuf_1
X_06393_ _06472_/A _06393_/B VGND VGND VPWR VPWR _06395_/A sky130_fd_sc_hd__or2_1
X_09181_ _09179_/Y _09180_/Y _08750_/A _09420_/C VGND VGND VPWR VPWR _09182_/B sky130_fd_sc_hd__a31o_1
XFILLER_186_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08132_ _09503_/A _08094_/X _09479_/A _08095_/X VGND VGND VPWR VPWR _08132_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05344_ _06780_/B _05357_/B VGND VGND VPWR VPWR _05549_/A sky130_fd_sc_hd__or2_4
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05275_ _05286_/A _05275_/B VGND VGND VPWR VPWR _06290_/A sky130_fd_sc_hd__or2_2
X_08063_ _07407_/Y _08058_/X _07327_/Y _08059_/X _08062_/X VGND VGND VPWR VPWR _08099_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07014_ _07009_/Y _05793_/A _07010_/Y _06502_/A _07013_/X VGND VGND VPWR VPWR _07027_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08965_ _08965_/A VGND VGND VPWR VPWR _09372_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07916_ _07209_/Y _07777_/X _07265_/Y _07778_/X _07915_/X VGND VGND VPWR VPWR _07937_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08896_ _09083_/C VGND VGND VPWR VPWR _09045_/C sky130_fd_sc_hd__inv_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07847_ _06722_/Y _07805_/X _06725_/Y _07758_/X _07846_/X VGND VGND VPWR VPWR _07848_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07778_ _07778_/A VGND VGND VPWR VPWR _07778_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09517_ _09517_/A VGND VGND VPWR VPWR _09518_/A sky130_fd_sc_hd__clkbuf_1
X_06729_ _10252_/Q VGND VGND VPWR VPWR _06729_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _08858_/A _09260_/A _08714_/X _09119_/Y VGND VGND VPWR VPWR _09448_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _09379_/A _09379_/B VGND VGND VPWR VPWR _09380_/B sky130_fd_sc_hd__or2_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10223_ _10349_/CLK _10223_/D repeater405/X VGND VGND VPWR VPWR _10223_/Q sky130_fd_sc_hd__dfrtp_1
X_10154_ _10157_/CLK _10154_/D repeater406/X VGND VGND VPWR VPWR _10154_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10085_ _10374_/CLK _10085_/D repeater410/X VGND VGND VPWR VPWR _10085_/Q sky130_fd_sc_hd__dfrtp_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05060_ _10424_/Q _05041_/A _09642_/X _05042_/A VGND VGND VPWR VPWR _10424_/D sky130_fd_sc_hd__a22o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08753_/B _08750_/C VGND VGND VPWR VPWR _08751_/B sky130_fd_sc_hd__and3_1
X_05962_ _05962_/A VGND VGND VPWR VPWR _05962_/Y sky130_fd_sc_hd__inv_2
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05893_ _10168_/Q _05885_/A _09661_/A1 _05886_/A VGND VGND VPWR VPWR _10168_/D sky130_fd_sc_hd__a22o_1
X_07701_ _09497_/A _07634_/X _09507_/A _07635_/X VGND VGND VPWR VPWR _07701_/X sky130_fd_sc_hd__o22a_1
X_08681_ _08819_/B VGND VGND VPWR VPWR _09109_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_04913_ _05163_/B VGND VGND VPWR VPWR _06780_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07632_ _07792_/A VGND VGND VPWR VPWR _07632_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04844_ _05118_/B _05164_/B VGND VGND VPWR VPWR _04845_/A sky130_fd_sc_hd__or2_1
XFILLER_179_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09302_ _09317_/B _09252_/Y _09275_/X _09301_/X VGND VGND VPWR VPWR _09302_/Y sky130_fd_sc_hd__o211ai_1
X_07563_ _07813_/A VGND VGND VPWR VPWR _07653_/A sky130_fd_sc_hd__buf_2
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06514_ _09841_/Q _06505_/A _09659_/A1 _06506_/A VGND VGND VPWR VPWR _09841_/D sky130_fd_sc_hd__a22o_1
X_07494_ _07494_/A VGND VGND VPWR VPWR _07495_/A sky130_fd_sc_hd__buf_2
XFILLER_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09233_ _09233_/A _09247_/B _09233_/C VGND VGND VPWR VPWR _09233_/Y sky130_fd_sc_hd__nor3_4
XFILLER_166_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06445_ _09873_/Q _06440_/X _09579_/X _06442_/X VGND VGND VPWR VPWR _09873_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09164_ _09010_/X _09020_/A _08661_/A _08674_/X VGND VGND VPWR VPWR _09446_/C sky130_fd_sc_hd__o22ai_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08115_ _07282_/Y _08092_/X _07690_/A _08093_/X _08114_/X VGND VGND VPWR VPWR _08116_/D
+ sky130_fd_sc_hd__o221a_1
X_06376_ _06374_/X _09611_/X _09650_/X _09918_/Q VGND VGND VPWR VPWR _09918_/D sky130_fd_sc_hd__o22a_1
XFILLER_162_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09095_ _09095_/A VGND VGND VPWR VPWR _09226_/B sky130_fd_sc_hd__inv_2
X_05327_ _05327_/A _05349_/B VGND VGND VPWR VPWR _06392_/A sky130_fd_sc_hd__or2_1
X_05258_ _05254_/Y _06078_/A _05256_/Y _06121_/A VGND VGND VPWR VPWR _05258_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08046_ _08046_/A _10002_/Q _08046_/C _10006_/Q VGND VGND VPWR VPWR _08214_/A sky130_fd_sc_hd__or4_4
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05189_ _10185_/Q VGND VGND VPWR VPWR _05189_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_135_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09997_ _10000_/CLK _09997_/D repeater410/X VGND VGND VPWR VPWR _09997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08948_ _08948_/A _09309_/B VGND VGND VPWR VPWR _08950_/A sky130_fd_sc_hd__or2_1
X_08879_ _08879_/A VGND VGND VPWR VPWR _09222_/A sky130_fd_sc_hd__inv_2
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10206_ _10354_/CLK _10206_/D repeater406/X VGND VGND VPWR VPWR _10206_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10137_ _10374_/CLK _10137_/D _07492_/B VGND VGND VPWR VPWR _10137_/Q sky130_fd_sc_hd__dfrtp_1
X_10068_ _10349_/CLK _10068_/D repeater405/X VGND VGND VPWR VPWR _10068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06230_ _07534_/A _07612_/C VGND VGND VPWR VPWR _07768_/A sky130_fd_sc_hd__or2_1
XFILLER_129_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06161_ _10016_/Q _06155_/X _09547_/A1 _06157_/X VGND VGND VPWR VPWR _10016_/D sky130_fd_sc_hd__a22o_1
X_06092_ _10047_/Q _06088_/X _06683_/B1 _06089_/Y VGND VGND VPWR VPWR _10047_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05112_ _05112_/A VGND VGND VPWR VPWR _05112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05043_ _10429_/Q _05040_/X _09656_/X _05042_/X VGND VGND VPWR VPWR _10429_/D sky130_fd_sc_hd__a22o_1
X_09920_ _10224_/CLK _09920_/D repeater405/X VGND VGND VPWR VPWR _09920_/Q sky130_fd_sc_hd__dfstp_1
X_09851_ _10157_/CLK _09851_/D repeater406/X VGND VGND VPWR VPWR _09851_/Q sky130_fd_sc_hd__dfstp_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _10382_/CLK _09782_/D _06662_/X VGND VGND VPWR VPWR _09787_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06994_ _06992_/Y _06167_/B _06993_/Y _06430_/B VGND VGND VPWR VPWR _06994_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08802_ _08847_/B VGND VGND VPWR VPWR _09253_/B sky130_fd_sc_hd__clkinv_4
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08733_/A _09175_/A VGND VGND VPWR VPWR _08733_/X sky130_fd_sc_hd__and2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05945_ _10139_/Q _05941_/X _09580_/X _05943_/X VGND VGND VPWR VPWR _10139_/D sky130_fd_sc_hd__a22o_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05876_ _05876_/A VGND VGND VPWR VPWR _05876_/Y sky130_fd_sc_hd__inv_2
X_08664_ _08679_/B _08672_/B VGND VGND VPWR VPWR _08841_/B sky130_fd_sc_hd__or2_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _09030_/A _08595_/B VGND VGND VPWR VPWR _08596_/B sky130_fd_sc_hd__and2_1
X_07615_ _07615_/A _07615_/B _07615_/C _07615_/D VGND VGND VPWR VPWR _07616_/C sky130_fd_sc_hd__and4_1
X_04827_ _05031_/A _04827_/B VGND VGND VPWR VPWR _04827_/X sky130_fd_sc_hd__or2_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07546_ _09991_/Q _07551_/B _07546_/C VGND VGND VPWR VPWR _07574_/B sky130_fd_sc_hd__or3_1
XFILLER_179_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09216_ _08385_/B _08484_/Y _09102_/A _08398_/C _09036_/B VGND VGND VPWR VPWR _09374_/B
+ sky130_fd_sc_hd__a41o_1
X_07477_ _07477_/A _09554_/X _07477_/C VGND VGND VPWR VPWR _07479_/A sky130_fd_sc_hd__or3_1
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06428_ _09650_/X _07477_/A _06427_/Y _06417_/A _09881_/Q VGND VGND VPWR VPWR _09881_/D
+ sky130_fd_sc_hd__a32o_1
X_09147_ _09226_/A _08753_/B _08750_/C _08751_/B VGND VGND VPWR VPWR _09329_/A sky130_fd_sc_hd__a31o_1
X_06359_ _06359_/A VGND VGND VPWR VPWR _06360_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_146_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09078_ _09078_/A _09357_/C _09291_/C _09427_/C VGND VGND VPWR VPWR _09081_/A sky130_fd_sc_hd__or4_4
XFILLER_146_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08029_ _05283_/Y _08195_/A _05310_/Y _08196_/A VGND VGND VPWR VPWR _08029_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 _10454_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_2
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05730_ _05730_/A VGND VGND VPWR VPWR _05731_/A sky130_fd_sc_hd__inv_2
X_05661_ _10302_/Q _05654_/A _09576_/X _05655_/A VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__a22o_1
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07400_ _10160_/Q VGND VGND VPWR VPWR _07400_/Y sky130_fd_sc_hd__inv_2
X_08380_ _08621_/C VGND VGND VPWR VPWR _08980_/C sky130_fd_sc_hd__inv_2
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07331_ _09975_/Q VGND VGND VPWR VPWR _07663_/A sky130_fd_sc_hd__inv_2
X_05592_ _06585_/A _05592_/B VGND VGND VPWR VPWR _06589_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07262_ _07262_/A _07262_/B _07262_/C VGND VGND VPWR VPWR _07288_/C sky130_fd_sc_hd__and3_1
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09001_ _09001_/A VGND VGND VPWR VPWR _09023_/A sky130_fd_sc_hd__buf_4
X_07193_ _07193_/A _07193_/B _07187_/X _07192_/X VGND VGND VPWR VPWR _07289_/B sky130_fd_sc_hd__or4bb_1
X_06213_ _09998_/Q _06207_/X _09547_/A1 _06209_/X VGND VGND VPWR VPWR _09998_/D sky130_fd_sc_hd__a22o_1
X_06144_ _06140_/B _06137_/X _06140_/A _06142_/X _06143_/Y VGND VGND VPWR VPWR _10023_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06075_ _10057_/Q _06068_/A _06683_/B1 _06069_/A VGND VGND VPWR VPWR _10057_/D sky130_fd_sc_hd__a22o_1
X_09903_ _10353_/CLK _09903_/D repeater403/X VGND VGND VPWR VPWR _09903_/Q sky130_fd_sc_hd__dfrtp_1
X_05026_ _10432_/Q _05020_/X _09536_/A3 _05021_/Y VGND VGND VPWR VPWR _10432_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09834_ _10062_/CLK _09834_/D repeater410/X VGND VGND VPWR VPWR _09834_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06977_ _06975_/Y _06304_/B _06976_/Y _06401_/A VGND VGND VPWR VPWR _06977_/X sky130_fd_sc_hd__o22a_1
X_09765_ _09919_/CLK _09765_/D VGND VGND VPWR VPWR _09765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05928_ _06011_/A _05928_/B VGND VGND VPWR VPWR _05930_/A sky130_fd_sc_hd__or2_2
X_09696_ _09404_/Y _09376_/X _09698_/S VGND VGND VPWR VPWR _09696_/X sky130_fd_sc_hd__mux2_1
X_08716_ _08661_/A _09260_/A _08715_/X VGND VGND VPWR VPWR _08719_/A sky130_fd_sc_hd__o21ai_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08647_ _08851_/B VGND VGND VPWR VPWR _08855_/A sky130_fd_sc_hd__clkbuf_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05859_ _10189_/Q _05853_/X _09547_/A1 _05855_/X VGND VGND VPWR VPWR _10189_/D sky130_fd_sc_hd__a22o_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _08586_/A _08578_/B VGND VGND VPWR VPWR _09162_/A sky130_fd_sc_hd__or2_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _07554_/C VGND VGND VPWR VPWR _07562_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10471_ _10471_/CLK _10471_/D _05034_/A VGND VGND VPWR VPWR _10471_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_6_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_csclk _09582_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06900_ _10164_/Q VGND VGND VPWR VPWR _06900_/Y sky130_fd_sc_hd__inv_2
X_07880_ _05339_/Y _07816_/X _05256_/Y _07817_/X _07879_/X VGND VGND VPWR VPWR _07885_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06831_ _06829_/Y _06360_/B _06830_/Y _05762_/B VGND VGND VPWR VPWR _06831_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09550_ _09550_/A0 _10303_/Q _09677_/S VGND VGND VPWR VPWR _09550_/X sky130_fd_sc_hd__mux2_1
X_06762_ _06763_/A VGND VGND VPWR VPWR _06762_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09481_ _09481_/A VGND VGND VPWR VPWR _09482_/A sky130_fd_sc_hd__clkbuf_1
X_08501_ _09103_/A VGND VGND VPWR VPWR _09005_/A sky130_fd_sc_hd__clkbuf_2
X_05713_ _05713_/A _06593_/B VGND VGND VPWR VPWR _05713_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08432_ _08530_/D _08430_/B _08431_/B VGND VGND VPWR VPWR _08695_/B sky130_fd_sc_hd__a21o_1
X_06693_ _06693_/A VGND VGND VPWR VPWR _09679_/S sky130_fd_sc_hd__buf_6
X_05644_ _10314_/Q _05640_/X _09580_/X _05642_/X VGND VGND VPWR VPWR _10314_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08363_ _09788_/Q _08363_/B VGND VGND VPWR VPWR _08363_/X sky130_fd_sc_hd__and2_1
XFILLER_189_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05575_ _05575_/A VGND VGND VPWR VPWR _05576_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08294_ _07092_/Y _08219_/X _07138_/Y _08220_/X _08293_/X VGND VGND VPWR VPWR _08310_/A
+ sky130_fd_sc_hd__o221a_1
X_07314_ input124/X _05101_/A _10433_/Q _05121_/Y _07313_/X VGND VGND VPWR VPWR _07317_/C
+ sky130_fd_sc_hd__a221o_1
X_07245_ _10213_/Q VGND VGND VPWR VPWR _07245_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07176_ _10047_/Q VGND VGND VPWR VPWR _07176_/Y sky130_fd_sc_hd__inv_4
XFILLER_191_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06127_ _10026_/Q _06123_/X _06683_/B1 _06124_/Y VGND VGND VPWR VPWR _10026_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06058_ _10070_/Q _06055_/X _09581_/X _06057_/X VGND VGND VPWR VPWR _10070_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05009_ _05009_/A VGND VGND VPWR VPWR _05010_/A sky130_fd_sc_hd__inv_2
X_09817_ _10238_/CLK _09817_/D repeater406/X VGND VGND VPWR VPWR _09817_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _09752_/CLK _09748_/D VGND VGND VPWR VPWR _09748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _05677_/B split1/X _09679_/S VGND VGND VPWR VPWR _09679_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_2
XFILLER_168_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10454_ _10486_/CLK _10454_/D _05034_/A VGND VGND VPWR VPWR _10454_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_182_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10385_ _04811_/A1 _10385_/D _05483_/X VGND VGND VPWR VPWR _10385_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05360_ _09862_/Q VGND VGND VPWR VPWR _05360_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05291_ _10128_/Q VGND VGND VPWR VPWR _05291_/Y sky130_fd_sc_hd__inv_2
X_07030_ _07030_/A VGND VGND VPWR VPWR _07030_/X sky130_fd_sc_hd__buf_1
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08981_ _08981_/A _09035_/B VGND VGND VPWR VPWR _08982_/B sky130_fd_sc_hd__or2_1
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07932_ _07932_/A _07932_/B VGND VGND VPWR VPWR _07932_/X sky130_fd_sc_hd__or2_1
X_07863_ _05348_/Y _07779_/X _07861_/Y _07781_/X _07862_/X VGND VGND VPWR VPWR _07863_/X
+ sky130_fd_sc_hd__o221a_1
X_06814_ _06814_/A _06814_/B _06814_/C _06814_/D VGND VGND VPWR VPWR _06814_/X sky130_fd_sc_hd__and4_2
X_09602_ _08238_/Y _10336_/Q _09700_/S VGND VGND VPWR VPWR _09602_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09533_ _09533_/A _09535_/B VGND VGND VPWR VPWR _09784_/D sky130_fd_sc_hd__nor2_1
X_07794_ _07794_/A VGND VGND VPWR VPWR _07794_/X sky130_fd_sc_hd__clkbuf_2
X_06745_ _10218_/Q VGND VGND VPWR VPWR _06745_/Y sky130_fd_sc_hd__clkinv_2
X_09464_ _09464_/A VGND VGND VPWR VPWR _09464_/X sky130_fd_sc_hd__clkbuf_1
X_06676_ _06676_/A VGND VGND VPWR VPWR _06676_/X sky130_fd_sc_hd__clkbuf_1
X_08415_ _08644_/A _08408_/Y _08485_/A _08408_/A _08895_/A VGND VGND VPWR VPWR _08565_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09395_ _09395_/A _09395_/B VGND VGND VPWR VPWR _09395_/X sky130_fd_sc_hd__or2_1
X_05627_ _05628_/A VGND VGND VPWR VPWR _05627_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08346_ _09806_/Q VGND VGND VPWR VPWR _08346_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05558_ _10360_/Q _05551_/X _09658_/A1 _05553_/X VGND VGND VPWR VPWR _10360_/D sky130_fd_sc_hd__a22o_1
X_05489_ _08354_/A _05489_/B VGND VGND VPWR VPWR _05489_/X sky130_fd_sc_hd__and2_1
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08277_ _07239_/Y _08179_/X _07213_/Y _08180_/X VGND VGND VPWR VPWR _08277_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07228_ _10052_/Q VGND VGND VPWR VPWR _07228_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07159_ _07159_/A VGND VGND VPWR VPWR _07159_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_16_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10353_/CLK sky130_fd_sc_hd__clkbuf_16
X_10170_ _10313_/CLK _10170_/D repeater403/X VGND VGND VPWR VPWR _10170_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10506_ _10508_/CLK _10506_/D repeater402/X VGND VGND VPWR VPWR _10506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10437_ _10478_/CLK _10437_/D _05034_/A VGND VGND VPWR VPWR _10437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10368_ _10500_/CLK _10368_/D repeater407/X VGND VGND VPWR VPWR _10368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10382_/CLK _10299_/D _05665_/X VGND VGND VPWR VPWR _10299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater406 repeater407/X VGND VGND VPWR VPWR repeater406/X sky130_fd_sc_hd__buf_12
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04860_ _10501_/Q _04851_/A _09589_/X _04852_/A VGND VGND VPWR VPWR _10501_/D sky130_fd_sc_hd__o22a_1
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06530_ _06531_/A VGND VGND VPWR VPWR _06530_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06461_ _06461_/A _06461_/B input164/X VGND VGND VPWR VPWR _06465_/C sky130_fd_sc_hd__or3b_1
XFILLER_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05412_ hold50/A _05396_/X hold44/A _05398_/X VGND VGND VPWR VPWR _10414_/D sky130_fd_sc_hd__a22o_1
X_08200_ _08200_/A VGND VGND VPWR VPWR _08200_/X sky130_fd_sc_hd__buf_2
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09180_ _09180_/A VGND VGND VPWR VPWR _09180_/Y sky130_fd_sc_hd__clkinv_2
X_06392_ _06392_/A VGND VGND VPWR VPWR _06393_/B sky130_fd_sc_hd__clkbuf_4
X_08131_ _09467_/A _08086_/X _09507_/A _08087_/X _08130_/X VGND VGND VPWR VPWR _08134_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05343_ _10357_/Q VGND VGND VPWR VPWR _05343_/Y sky130_fd_sc_hd__clkinv_4
X_05274_ _09960_/Q VGND VGND VPWR VPWR _05274_/Y sky130_fd_sc_hd__clkinv_4
X_08062_ _07394_/Y _08060_/X _07356_/Y _08061_/X VGND VGND VPWR VPWR _08062_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07013_ _07011_/Y _05830_/B _07012_/Y _06329_/B VGND VGND VPWR VPWR _07013_/X sky130_fd_sc_hd__o22a_1
XFILLER_161_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08964_ _08964_/A _09311_/B VGND VGND VPWR VPWR _08967_/A sky130_fd_sc_hd__or2_1
X_07915_ _07203_/Y _07779_/X _07913_/Y _07781_/X _07914_/X VGND VGND VPWR VPWR _07915_/X
+ sky130_fd_sc_hd__o221a_1
X_08895_ _08895_/A _08895_/B _08895_/C VGND VGND VPWR VPWR _09083_/C sky130_fd_sc_hd__or3_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07846_ _06735_/Y _07806_/X _06728_/Y _07807_/X VGND VGND VPWR VPWR _07846_/X sky130_fd_sc_hd__o22a_1
X_07777_ _07777_/A VGND VGND VPWR VPWR _07777_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04989_ _10452_/Q _04981_/A _06684_/B1 _04982_/A VGND VGND VPWR VPWR _10452_/D sky130_fd_sc_hd__a22o_1
X_09516_ _09516_/A VGND VGND VPWR VPWR _09516_/X sky130_fd_sc_hd__clkbuf_1
X_06728_ _10495_/Q VGND VGND VPWR VPWR _06728_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _09447_/A _09447_/B _09447_/C _09447_/D VGND VGND VPWR VPWR _09447_/X sky130_fd_sc_hd__or4_1
XFILLER_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06659_ _06663_/A VGND VGND VPWR VPWR _06660_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09378_ _09378_/A _09378_/B _09378_/C _09378_/D VGND VGND VPWR VPWR _09447_/D sky130_fd_sc_hd__or4_2
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08329_ _09771_/Q _09774_/Q VGND VGND VPWR VPWR _08329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10222_ _10224_/CLK _10222_/D repeater405/X VGND VGND VPWR VPWR _10222_/Q sky130_fd_sc_hd__dfrtp_1
X_10153_ _10411_/CLK _10153_/D repeater407/X VGND VGND VPWR VPWR _10153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10084_ _10374_/CLK _10084_/D hold41/X VGND VGND VPWR VPWR _10084_/Q sky130_fd_sc_hd__dfrtp_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07700_ _09469_/A _07627_/X _09461_/A _07628_/X _07699_/X VGND VGND VPWR VPWR _07707_/A
+ sky130_fd_sc_hd__o221a_1
X_05961_ _05962_/A VGND VGND VPWR VPWR _05961_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05892_ _10169_/Q _05885_/A _09660_/A1 _05886_/A VGND VGND VPWR VPWR _10169_/D sky130_fd_sc_hd__a22o_1
X_08680_ _08807_/A VGND VGND VPWR VPWR _08819_/B sky130_fd_sc_hd__clkbuf_2
X_04912_ _04992_/A VGND VGND VPWR VPWR _05163_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07631_ _07350_/Y _07627_/X _07327_/Y _07628_/X _07630_/X VGND VGND VPWR VPWR _07650_/A
+ sky130_fd_sc_hd__o221a_1
X_04843_ _05213_/A _09672_/X _05135_/C VGND VGND VPWR VPWR _05164_/B sky130_fd_sc_hd__or3_4
X_07562_ _07584_/B _07562_/B VGND VGND VPWR VPWR _07813_/A sky130_fd_sc_hd__or2_1
X_09301_ _09362_/B _09362_/C _09363_/B _09300_/X VGND VGND VPWR VPWR _09301_/X sky130_fd_sc_hd__or4b_2
X_06513_ _09842_/Q _06505_/A _09661_/A1 _06506_/A VGND VGND VPWR VPWR _09842_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07493_ _10298_/Q input86/X VGND VGND VPWR VPWR _07494_/A sky130_fd_sc_hd__or2b_1
XFILLER_34_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09232_ _09231_/Y _09225_/Y _09237_/A _09152_/A VGND VGND VPWR VPWR _09235_/C sky130_fd_sc_hd__a31o_1
X_06444_ _09874_/Q _06440_/X _09580_/X _06442_/X VGND VGND VPWR VPWR _09874_/D sky130_fd_sc_hd__a22o_1
X_09163_ _09163_/A _09163_/B VGND VGND VPWR VPWR _09167_/A sky130_fd_sc_hd__or2_1
X_06375_ _09919_/Q _09650_/X _09613_/X _06374_/X VGND VGND VPWR VPWR _09919_/D sky130_fd_sc_hd__o22a_1
X_05326_ _09902_/Q VGND VGND VPWR VPWR _05326_/Y sky130_fd_sc_hd__inv_2
X_08114_ _07220_/Y _08094_/X _07270_/Y _08095_/X VGND VGND VPWR VPWR _08114_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09094_ _08788_/B _09105_/B _08865_/X VGND VGND VPWR VPWR _09343_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05257_ _05333_/A _05316_/B VGND VGND VPWR VPWR _06121_/A sky130_fd_sc_hd__or2_1
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08045_ _08046_/A _10002_/Q _08045_/C _08045_/D VGND VGND VPWR VPWR _08213_/A sky130_fd_sc_hd__or4_4
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05188_ _05188_/A VGND VGND VPWR VPWR _05785_/B sky130_fd_sc_hd__buf_2
XFILLER_103_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09996_ _10364_/CLK _09996_/D repeater410/X VGND VGND VPWR VPWR _09996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08947_ _08947_/A VGND VGND VPWR VPWR _09309_/B sky130_fd_sc_hd__inv_2
X_08878_ _08878_/A _09348_/B VGND VGND VPWR VPWR _08993_/A sky130_fd_sc_hd__or2_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07829_ _07829_/A VGND VGND VPWR VPWR _07829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10205_ _10513_/CLK _10205_/D _07492_/B VGND VGND VPWR VPWR _10205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10136_ _10374_/CLK _10136_/D _07492_/B VGND VGND VPWR VPWR _10136_/Q sky130_fd_sc_hd__dfrtp_4
X_10067_ _10350_/CLK _10067_/D repeater405/X VGND VGND VPWR VPWR _10067_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06160_ _10017_/Q _06155_/X _09579_/X _06157_/X VGND VGND VPWR VPWR _10017_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06091_ _10048_/Q _06088_/X _09658_/A1 _06089_/Y VGND VGND VPWR VPWR _10048_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05111_ _05157_/A _05284_/B VGND VGND VPWR VPWR _05112_/A sky130_fd_sc_hd__nor2_2
X_05042_ _05042_/A VGND VGND VPWR VPWR _05042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09850_ _10354_/CLK _09850_/D repeater406/X VGND VGND VPWR VPWR _09850_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09781_/CLK _09781_/D _06664_/X VGND VGND VPWR VPWR _09781_/Q sky130_fd_sc_hd__dfstp_1
X_08801_ _09337_/A _08980_/B _08801_/C VGND VGND VPWR VPWR _09420_/B sky130_fd_sc_hd__and3_2
X_06993_ _09880_/Q VGND VGND VPWR VPWR _06993_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_112_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08732_/A _08855_/A VGND VGND VPWR VPWR _09175_/A sky130_fd_sc_hd__or2_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05944_ _10140_/Q _05941_/X _09581_/X _05943_/X VGND VGND VPWR VPWR _10140_/D sky130_fd_sc_hd__a22o_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _09233_/A _08781_/B _08668_/A VGND VGND VPWR VPWR _08679_/B sky130_fd_sc_hd__or3_4
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05875_ _05876_/A VGND VGND VPWR VPWR _05875_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _09327_/A _08594_/B VGND VGND VPWR VPWR _08595_/B sky130_fd_sc_hd__nor2_1
X_07614_ _05310_/Y _07825_/A _07609_/Y _07827_/A _07613_/X VGND VGND VPWR VPWR _07615_/D
+ sky130_fd_sc_hd__o221a_1
X_04826_ _06635_/A VGND VGND VPWR VPWR _05031_/A sky130_fd_sc_hd__clkbuf_2
X_07545_ _07802_/A VGND VGND VPWR VPWR _07642_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_179_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07476_ _07565_/A _07582_/B VGND VGND VPWR VPWR _07476_/Y sky130_fd_sc_hd__nor2_2
X_09215_ _08546_/A _08548_/A _08504_/B _09000_/B _08598_/A VGND VGND VPWR VPWR _09312_/B
+ sky130_fd_sc_hd__o221ai_1
X_06427_ _09682_/X VGND VGND VPWR VPWR _06427_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06358_ _09928_/Q _06352_/X _09574_/X _06353_/Y VGND VGND VPWR VPWR _09928_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09146_ _09223_/A _09229_/B VGND VGND VPWR VPWR _09415_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05309_ _05302_/Y _05761_/A _05304_/Y _05793_/A _05308_/X VGND VGND VPWR VPWR _05321_/C
+ sky130_fd_sc_hd__o221a_1
X_09077_ _09420_/D _09214_/B VGND VGND VPWR VPWR _09427_/C sky130_fd_sc_hd__or2_1
X_06289_ _10020_/Q _09778_/Q _06288_/Y _09968_/Q _06264_/A VGND VGND VPWR VPWR _09968_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08028_ _08034_/A _08044_/A _08040_/C VGND VGND VPWR VPWR _08196_/A sky130_fd_sc_hd__or3_4
XFILLER_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09979_ _10350_/CLK _09979_/D repeater405/X VGND VGND VPWR VPWR _09979_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10119_ _10119_/CLK _10119_/D repeater402/X VGND VGND VPWR VPWR _10119_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05660_ _10303_/Q _05653_/X _09550_/A0 _05655_/X VGND VGND VPWR VPWR _10303_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05591_ _09772_/Q _09773_/Q VGND VGND VPWR VPWR _05592_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07330_ _07325_/Y _06339_/B _07326_/Y _06053_/A _07329_/X VGND VGND VPWR VPWR _07349_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_188_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07261_ _07256_/Y _06010_/A _07257_/Y _06339_/B _07260_/X VGND VGND VPWR VPWR _07262_/C
+ sky130_fd_sc_hd__o221a_1
X_09000_ _09103_/A _09000_/B VGND VGND VPWR VPWR _09001_/A sky130_fd_sc_hd__or2_1
XFILLER_176_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07192_ _07188_/Y _06066_/B _07189_/Y _06108_/B _07191_/X VGND VGND VPWR VPWR _07192_/X
+ sky130_fd_sc_hd__o221a_1
X_06212_ _09999_/Q _06207_/X _09579_/X _06209_/X VGND VGND VPWR VPWR _09999_/D sky130_fd_sc_hd__a22o_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06143_ _06140_/B _06137_/X _06140_/A VGND VGND VPWR VPWR _06143_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06074_ _10058_/Q _06067_/X _09658_/A1 _06069_/X VGND VGND VPWR VPWR _10058_/D sky130_fd_sc_hd__a22o_1
X_09902_ _10353_/CLK _09902_/D repeater406/X VGND VGND VPWR VPWR _09902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05025_ _10433_/Q _05020_/X _06684_/B1 _05021_/Y VGND VGND VPWR VPWR _10433_/D sky130_fd_sc_hd__a22o_1
X_09833_ _10062_/CLK _09833_/D repeater410/X VGND VGND VPWR VPWR _09833_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06976_ _09898_/Q VGND VGND VPWR VPWR _06976_/Y sky130_fd_sc_hd__inv_2
X_09764_ _09919_/CLK _09764_/D VGND VGND VPWR VPWR _09764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05927_ _05927_/A VGND VGND VPWR VPWR _05928_/B sky130_fd_sc_hd__buf_2
X_09695_ _09367_/Y _09316_/X _09698_/S VGND VGND VPWR VPWR _09695_/X sky130_fd_sc_hd__mux2_1
X_08715_ _08743_/A _08836_/B _08712_/X _09118_/A _08714_/X VGND VGND VPWR VPWR _08715_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08786_/B _08809_/A VGND VGND VPWR VPWR _08851_/B sky130_fd_sc_hd__or2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05858_ _10190_/Q _05853_/X _09579_/X _05855_/X VGND VGND VPWR VPWR _10190_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04809_ _10281_/Q input77/X _09521_/B VGND VGND VPWR VPWR _09705_/A sky130_fd_sc_hd__mux2_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05789_ _10230_/Q _05786_/X _09577_/X _05787_/Y VGND VGND VPWR VPWR _10230_/D sky130_fd_sc_hd__a22o_1
X_08577_ _08585_/A _08578_/B VGND VGND VPWR VPWR _08577_/X sky130_fd_sc_hd__or2_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _07528_/A _09990_/Q VGND VGND VPWR VPWR _07602_/C sky130_fd_sc_hd__or2_1
X_07459_ _07290_/X _07452_/A _09736_/Q _07453_/A VGND VGND VPWR VPWR _09736_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10470_ _10471_/CLK _10470_/D _05034_/A VGND VGND VPWR VPWR _10470_/Q sky130_fd_sc_hd__dfrtp_4
X_09129_ _09342_/C VGND VGND VPWR VPWR _09129_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06830_ _10243_/Q VGND VGND VPWR VPWR _06830_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06761_ _07450_/A _06761_/B VGND VGND VPWR VPWR _06763_/A sky130_fd_sc_hd__or2_2
X_09480_ _09480_/A VGND VGND VPWR VPWR _09480_/X sky130_fd_sc_hd__clkbuf_1
X_08500_ _09155_/A VGND VGND VPWR VPWR _09103_/A sky130_fd_sc_hd__clkbuf_2
X_05712_ _05712_/A VGND VGND VPWR VPWR _05712_/X sky130_fd_sc_hd__clkbuf_1
X_06692_ _06692_/A VGND VGND VPWR VPWR _06692_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08431_ _09233_/A _08431_/B VGND VGND VPWR VPWR _08476_/B sky130_fd_sc_hd__nor2_1
X_05643_ _10315_/Q _05640_/X _09581_/X _05642_/X VGND VGND VPWR VPWR _10315_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08362_ _09790_/Q input183/X _09789_/Q input166/X _08361_/X VGND VGND VPWR VPWR _08362_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05574_ _10351_/Q _05568_/X _09659_/A1 _05569_/Y VGND VGND VPWR VPWR _10351_/D sky130_fd_sc_hd__a22o_1
X_08293_ _07071_/Y _08173_/A _07152_/Y _08174_/A VGND VGND VPWR VPWR _08293_/X sky130_fd_sc_hd__o22a_1
X_07313_ _09767_/Q _05146_/Y _10046_/Q _05084_/Y VGND VGND VPWR VPWR _07313_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07244_ _10498_/Q VGND VGND VPWR VPWR _07244_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07175_ input58/X _06693_/A input13/X _06698_/A _07174_/X VGND VGND VPWR VPWR _07181_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06126_ _10027_/Q _06123_/X _09577_/X _06124_/Y VGND VGND VPWR VPWR _10027_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06057_ _06057_/A VGND VGND VPWR VPWR _06057_/X sky130_fd_sc_hd__clkbuf_2
X_05008_ _05009_/A VGND VGND VPWR VPWR _05008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09816_ _10353_/CLK _09816_/D repeater403/X VGND VGND VPWR VPWR _09816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09747_ _09752_/CLK _09747_/D VGND VGND VPWR VPWR _09747_/Q sky130_fd_sc_hd__dfxtp_1
X_06959_ _06954_/Y _05549_/A _06955_/Y _06551_/B _06958_/X VGND VGND VPWR VPWR _06960_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _10421_/Q _10481_/Q _10299_/Q VGND VGND VPWR VPWR _09678_/X sky130_fd_sc_hd__mux2_8
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08629_ _08757_/A VGND VGND VPWR VPWR _09223_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10453_ _10486_/CLK _10453_/D repeater409/X VGND VGND VPWR VPWR _10453_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10384_ _04811_/A1 _10384_/D _05498_/X VGND VGND VPWR VPWR _10384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05290_ _05282_/Y _04871_/B _05283_/Y _06010_/A _05289_/X VGND VGND VPWR VPWR _05321_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _09337_/A _08980_/B _08980_/C VGND VGND VPWR VPWR _09035_/B sky130_fd_sc_hd__and3_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07931_ _07196_/Y _07816_/X _07238_/Y _07817_/X _07930_/X VGND VGND VPWR VPWR _07936_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07862_ _05296_/Y _07782_/X _05192_/Y _07783_/X VGND VGND VPWR VPWR _07862_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06813_ _06808_/Y _06708_/B _06809_/Y _05550_/B _06812_/X VGND VGND VPWR VPWR _06814_/D
+ sky130_fd_sc_hd__o221a_1
X_09601_ _09600_/X _09912_/Q _09776_/Q VGND VGND VPWR VPWR _09601_/X sky130_fd_sc_hd__mux2_1
X_09532_ _09532_/A _09535_/B VGND VGND VPWR VPWR _09785_/D sky130_fd_sc_hd__nor2_1
X_07793_ _07793_/A VGND VGND VPWR VPWR _07793_/X sky130_fd_sc_hd__clkbuf_2
X_06744_ _06742_/Y _06503_/B _07854_/A _06267_/B VGND VGND VPWR VPWR _06744_/X sky130_fd_sc_hd__o22a_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ _09463_/A VGND VGND VPWR VPWR _09464_/A sky130_fd_sc_hd__clkbuf_1
X_06675_ _06677_/A VGND VGND VPWR VPWR _06676_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08414_ _08913_/A VGND VGND VPWR VPWR _08895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09394_ _09432_/B _09434_/A _09434_/B _09435_/A VGND VGND VPWR VPWR _09394_/X sky130_fd_sc_hd__or4_2
X_05626_ _05626_/A VGND VGND VPWR VPWR _05628_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05557_ _10361_/Q _05551_/X _09547_/A1 _05553_/X VGND VGND VPWR VPWR _10361_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08345_ _09805_/Q _08344_/B _08344_/Y VGND VGND VPWR VPWR _08345_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05488_ _09789_/Q VGND VGND VPWR VPWR _09534_/A sky130_fd_sc_hd__inv_2
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08276_ _07238_/Y _08219_/X _07203_/Y _08220_/X _08275_/X VGND VGND VPWR VPWR _08292_/A
+ sky130_fd_sc_hd__o221a_1
X_07227_ _10143_/Q VGND VGND VPWR VPWR _07227_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07158_ _07158_/A _07158_/B _07064_/X _07157_/X VGND VGND VPWR VPWR _07159_/A sky130_fd_sc_hd__or4bb_4
XFILLER_118_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06109_ _06110_/A VGND VGND VPWR VPWR _06109_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07089_ _07089_/A _07089_/B _07089_/C _07089_/D VGND VGND VPWR VPWR _07157_/A sky130_fd_sc_hd__and4_1
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10505_ _10508_/CLK _10505_/D repeater402/X VGND VGND VPWR VPWR _10505_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10436_ _10483_/CLK _10436_/D _05034_/A VGND VGND VPWR VPWR _10436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10367_ _10369_/CLK _10367_/D repeater407/X VGND VGND VPWR VPWR _10367_/Q sky130_fd_sc_hd__dfstp_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10298_ _10406_/CLK _10298_/D _05670_/X VGND VGND VPWR VPWR _10298_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater407 repeater409/X VGND VGND VPWR VPWR repeater407/X sky130_fd_sc_hd__buf_12
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06460_ _06460_/A _06460_/B input150/X input153/X VGND VGND VPWR VPWR _06465_/B sky130_fd_sc_hd__or4bb_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05411_ _05411_/A VGND VGND VPWR VPWR _05411_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08130_ _09471_/A _08088_/X _09509_/A _08089_/X VGND VGND VPWR VPWR _08130_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06391_ _09650_/X _07477_/A _06389_/Y _06390_/X _09907_/Q VGND VGND VPWR VPWR _09907_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05342_ _05332_/Y _05567_/B _05335_/Y _06502_/A _05341_/X VGND VGND VPWR VPWR _05364_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05273_ _10488_/Q VGND VGND VPWR VPWR _05273_/Y sky130_fd_sc_hd__clkinv_4
X_08061_ _08180_/A VGND VGND VPWR VPWR _08061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07012_ _09945_/Q VGND VGND VPWR VPWR _07012_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ _08972_/A _08968_/B VGND VGND VPWR VPWR _09311_/B sky130_fd_sc_hd__nor2_1
X_07914_ _07214_/Y _07782_/X _07277_/Y _07783_/X VGND VGND VPWR VPWR _07914_/X sky130_fd_sc_hd__o22a_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _08908_/B VGND VGND VPWR VPWR _09045_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_110_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07845_ _07842_/Y _07799_/X _07843_/Y _07801_/X _07844_/X VGND VGND VPWR VPWR _07848_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07776_ _07776_/A _07776_/B _07776_/C VGND VGND VPWR VPWR _07776_/Y sky130_fd_sc_hd__nand3_2
X_04988_ _10453_/Q _04981_/A _06683_/B1 _04982_/A VGND VGND VPWR VPWR _10453_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09515_ _09515_/A VGND VGND VPWR VPWR _09516_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06727_ _06722_/Y _06402_/B _06723_/Y _05550_/B _06726_/X VGND VGND VPWR VPWR _06740_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _09446_/A _09446_/B _09446_/C _09446_/D VGND VGND VPWR VPWR _09447_/B sky130_fd_sc_hd__or4_1
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06658_ _06658_/A VGND VGND VPWR VPWR _06658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09377_ _09377_/A _09377_/B _08543_/X VGND VGND VPWR VPWR _09378_/B sky130_fd_sc_hd__or3b_1
X_06589_ _09807_/Q _06589_/B _09808_/Q VGND VGND VPWR VPWR _06589_/X sky130_fd_sc_hd__and3_1
X_05609_ _10334_/Q _05604_/X _09579_/X _05606_/X VGND VGND VPWR VPWR _10334_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08328_ _08328_/A _08328_/B _08328_/C _08328_/D VGND VGND VPWR VPWR _08328_/Y sky130_fd_sc_hd__nand4_2
X_08259_ _07370_/Y _08179_/X _07364_/Y _08180_/X VGND VGND VPWR VPWR _08259_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10221_ _10224_/CLK _10221_/D repeater405/X VGND VGND VPWR VPWR _10221_/Q sky130_fd_sc_hd__dfrtp_1
X_10152_ _10257_/CLK _10152_/D repeater407/X VGND VGND VPWR VPWR _10152_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 _09538_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_2
X_10083_ _10135_/CLK _10083_/D hold41/X VGND VGND VPWR VPWR _10083_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10419_ _09572_/A1 _10419_/D _05387_/X VGND VGND VPWR VPWR _10419_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05960_ _05993_/A _05960_/B VGND VGND VPWR VPWR _05962_/A sky130_fd_sc_hd__or2_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05891_ _10170_/Q _05884_/X _09550_/A0 _05886_/X VGND VGND VPWR VPWR _10170_/D sky130_fd_sc_hd__a22o_1
X_04911_ _09663_/X _09672_/X _05213_/B VGND VGND VPWR VPWR _04992_/A sky130_fd_sc_hd__or3_2
X_07630_ _07394_/Y _07533_/C _07387_/Y _07629_/X VGND VGND VPWR VPWR _07630_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04842_ _04818_/Y _09666_/X _09665_/X VGND VGND VPWR VPWR _05135_/C sky130_fd_sc_hd__a21bo_1
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07561_ _07564_/C _07574_/B VGND VGND VPWR VPWR _07579_/A sky130_fd_sc_hd__or2_1
XFILLER_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ _09432_/B _09300_/B _09417_/A _09393_/A VGND VGND VPWR VPWR _09300_/X sky130_fd_sc_hd__or4_1
X_06512_ _09843_/Q _06505_/A _09660_/A1 _06506_/A VGND VGND VPWR VPWR _09843_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10238_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07492_ _10297_/Q _07492_/B VGND VGND VPWR VPWR _07492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09231_ _09231_/A VGND VGND VPWR VPWR _09231_/Y sky130_fd_sc_hd__clkinv_2
X_06443_ _09875_/Q _06440_/X _09581_/X _06442_/X VGND VGND VPWR VPWR _09875_/D sky130_fd_sc_hd__a22o_1
X_09162_ _09162_/A _09162_/B VGND VGND VPWR VPWR _09163_/B sky130_fd_sc_hd__nand2_1
X_06374_ _06417_/A VGND VGND VPWR VPWR _06374_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08113_ _07263_/Y _08086_/X _07184_/Y _08087_/X _08112_/X VGND VGND VPWR VPWR _08116_/C
+ sky130_fd_sc_hd__o221a_1
X_05325_ _05325_/A _05361_/B VGND VGND VPWR VPWR _05433_/A sky130_fd_sc_hd__or2_4
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09093_ _09093_/A _09344_/B VGND VGND VPWR VPWR _09399_/B sky130_fd_sc_hd__nor2_1
X_05256_ _10024_/Q VGND VGND VPWR VPWR _05256_/Y sky130_fd_sc_hd__inv_2
X_08044_ _08044_/A _08044_/B _10006_/Q VGND VGND VPWR VPWR _08212_/A sky130_fd_sc_hd__or3_4
X_05187_ _05313_/A _05292_/A VGND VGND VPWR VPWR _05188_/A sky130_fd_sc_hd__or2_1
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09995_ _10000_/CLK _09995_/D repeater410/X VGND VGND VPWR VPWR _09995_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08946_ _08972_/A _08951_/B VGND VGND VPWR VPWR _08947_/A sky130_fd_sc_hd__or2_1
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08877_ _08786_/A _09092_/A _08787_/B _09788_/Q VGND VGND VPWR VPWR _09348_/B sky130_fd_sc_hd__o31ai_4
XFILLER_57_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07828_ _07828_/A VGND VGND VPWR VPWR _07828_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07759_ _06888_/Y _07646_/X _06856_/Y _07647_/X VGND VGND VPWR VPWR _07759_/X sky130_fd_sc_hd__o22a_1
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09429_ _09352_/A _08858_/A _09352_/A _09352_/B VGND VGND VPWR VPWR _09429_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10204_ _10513_/CLK _10204_/D _07492_/B VGND VGND VPWR VPWR _10204_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10135_ _10135_/CLK _10135_/D _07492_/B VGND VGND VPWR VPWR _10135_/Q sky130_fd_sc_hd__dfrtp_1
X_10066_ _10350_/CLK _10066_/D repeater405/X VGND VGND VPWR VPWR _10066_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05110_ _05325_/A VGND VGND VPWR VPWR _05284_/B sky130_fd_sc_hd__buf_4
X_06090_ _10049_/Q _06088_/X _09545_/A1 _06089_/Y VGND VGND VPWR VPWR _10049_/D sky130_fd_sc_hd__a22o_1
X_05041_ _05041_/A VGND VGND VPWR VPWR _05042_/A sky130_fd_sc_hd__inv_2
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _09057_/A VGND VGND VPWR VPWR _08801_/C sky130_fd_sc_hd__inv_2
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06992_ _10011_/Q VGND VGND VPWR VPWR _06992_/Y sky130_fd_sc_hd__inv_2
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09780_/CLK _09780_/D _06667_/X VGND VGND VPWR VPWR _09780_/Q sky130_fd_sc_hd__dfstp_1
X_08731_ _08731_/A _09327_/B VGND VGND VPWR VPWR _08733_/A sky130_fd_sc_hd__nor2_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05943_ _05943_/A VGND VGND VPWR VPWR _05943_/X sky130_fd_sc_hd__clkbuf_2
X_08662_ _08662_/A VGND VGND VPWR VPWR _09253_/A sky130_fd_sc_hd__buf_4
X_05874_ _05874_/A _05874_/B VGND VGND VPWR VPWR _05876_/A sky130_fd_sc_hd__or2_1
X_07613_ _05197_/Y _07828_/A _05304_/Y _07829_/A VGND VGND VPWR VPWR _07613_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08593_ _09006_/A _08520_/B _08592_/Y VGND VGND VPWR VPWR _08594_/B sky130_fd_sc_hd__o21ai_1
X_04825_ _06679_/A VGND VGND VPWR VPWR _06635_/A sky130_fd_sc_hd__buf_4
XFILLER_179_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07544_ _07558_/A _07611_/A _07549_/B VGND VGND VPWR VPWR _07802_/A sky130_fd_sc_hd__or3_4
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07475_ _09991_/Q _07551_/B _07524_/A VGND VGND VPWR VPWR _07582_/B sky130_fd_sc_hd__or3_2
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09214_ _09327_/A _09214_/B _09214_/C VGND VGND VPWR VPWR _09405_/A sky130_fd_sc_hd__or3_2
X_06426_ _06390_/X _09615_/X _09650_/X _09882_/Q VGND VGND VPWR VPWR _09882_/D sky130_fd_sc_hd__o22a_1
XFILLER_167_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06357_ _09929_/Q _06352_/X hold46/X _06353_/Y VGND VGND VPWR VPWR _09929_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09145_ _09344_/A _09145_/B VGND VGND VPWR VPWR _09416_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05308_ _05308_/A _05882_/A VGND VGND VPWR VPWR _05308_/X sky130_fd_sc_hd__or2_1
X_09076_ _09076_/A _09311_/B VGND VGND VPWR VPWR _09291_/C sky130_fd_sc_hd__or2_1
X_06288_ _06288_/A VGND VGND VPWR VPWR _06288_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05239_ _10343_/Q VGND VGND VPWR VPWR _05239_/Y sky130_fd_sc_hd__clkinv_2
X_08027_ _08027_/A _08043_/B _08040_/C VGND VGND VPWR VPWR _08195_/A sky130_fd_sc_hd__or3_4
XFILLER_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09978_ _10000_/CLK _09978_/D repeater405/X VGND VGND VPWR VPWR _09978_/Q sky130_fd_sc_hd__dfrtp_1
X_08929_ _08929_/A _08943_/A VGND VGND VPWR VPWR _09354_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10118_ _10289_/CLK _10118_/D repeater402/X VGND VGND VPWR VPWR _10118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsplit1 hold1/A VGND VGND VPWR VPWR split1/X sky130_fd_sc_hd__buf_4
XFILLER_152_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10049_ _10127_/CLK _10049_/D repeater409/X VGND VGND VPWR VPWR _10049_/Q sky130_fd_sc_hd__dfstp_1
X_05590_ _09774_/Q VGND VGND VPWR VPWR _05590_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07260_ _07258_/Y _05229_/A _07259_/Y _06537_/A VGND VGND VPWR VPWR _07260_/X sky130_fd_sc_hd__o22a_1
X_07191_ _05139_/B _05333_/A _07190_/Y _06705_/A _06780_/X VGND VGND VPWR VPWR _07191_/X
+ sky130_fd_sc_hd__o221a_1
X_06211_ _10000_/Q _06207_/X _09580_/X _06209_/X VGND VGND VPWR VPWR _10000_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06142_ _06150_/A _06142_/B VGND VGND VPWR VPWR _06142_/X sky130_fd_sc_hd__or2_1
XFILLER_144_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06073_ _10059_/Q _06067_/X _09545_/A1 _06069_/X VGND VGND VPWR VPWR _10059_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09901_ _10310_/CLK _09901_/D repeater404/X VGND VGND VPWR VPWR _09901_/Q sky130_fd_sc_hd__dfrtp_1
X_05024_ _10434_/Q _05020_/X _06683_/B1 _05021_/Y VGND VGND VPWR VPWR _10434_/D sky130_fd_sc_hd__a22o_1
X_09832_ _10355_/CLK _09832_/D repeater406/X VGND VGND VPWR VPWR _09832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09763_ _09919_/CLK _09763_/D VGND VGND VPWR VPWR _09763_/Q sky130_fd_sc_hd__dfxtp_1
X_06975_ _09959_/Q VGND VGND VPWR VPWR _06975_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08714_ _08732_/A _08836_/B VGND VGND VPWR VPWR _08714_/X sky130_fd_sc_hd__or2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _09302_/Y _09221_/X _09698_/S VGND VGND VPWR VPWR _09694_/X sky130_fd_sc_hd__mux2_1
X_05926_ _06337_/A VGND VGND VPWR VPWR _06011_/A sky130_fd_sc_hd__buf_6
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _08645_/A _08668_/A VGND VGND VPWR VPWR _08809_/A sky130_fd_sc_hd__or2_2
X_05857_ _10191_/Q _05853_/X _09580_/X _05855_/X VGND VGND VPWR VPWR _10191_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08583_/A _08578_/B _08543_/X _08574_/X _09003_/A VGND VGND VPWR VPWR _08576_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_81_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04808_ _10266_/Q input67/X _10406_/Q VGND VGND VPWR VPWR _09707_/A sky130_fd_sc_hd__mux2_2
X_05788_ _10231_/Q _05786_/X _09578_/X _05787_/Y VGND VGND VPWR VPWR _10231_/D sky130_fd_sc_hd__a22o_1
X_07527_ _07527_/A VGND VGND VPWR VPWR _07533_/C sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07458_ _07159_/X _07451_/X _09737_/Q _07453_/X VGND VGND VPWR VPWR _09737_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ _10259_/Q VGND VGND VPWR VPWR _07389_/Y sky130_fd_sc_hd__inv_2
X_06409_ _09898_/Q _06403_/X _09547_/A1 _06405_/X VGND VGND VPWR VPWR _09898_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09128_ _09327_/B _09290_/A VGND VGND VPWR VPWR _09342_/C sky130_fd_sc_hd__or2_1
XFILLER_108_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09059_ _08851_/A _09048_/X _09049_/Y _08918_/X _09058_/X VGND VGND VPWR VPWR _09062_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput190 wb_dat_i[3] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__clkbuf_1
X_06760_ _09784_/Q VGND VGND VPWR VPWR _06761_/B sky130_fd_sc_hd__clkinv_4
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05711_ _06568_/A VGND VGND VPWR VPWR _05712_/A sky130_fd_sc_hd__clkbuf_1
X_06691_ _10114_/Q _05094_/Y _10450_/Q _06688_/X _06690_/X VGND VGND VPWR VPWR _06701_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08430_ _08530_/D _08430_/B VGND VGND VPWR VPWR _08431_/B sky130_fd_sc_hd__nor2_1
X_05642_ _05642_/A VGND VGND VPWR VPWR _05642_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08361_ _09788_/Q _08361_/B VGND VGND VPWR VPWR _08361_/X sky130_fd_sc_hd__and2_1
X_05573_ _10352_/Q _05568_/X _09661_/A1 _05569_/Y VGND VGND VPWR VPWR _10352_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08292_ _08292_/A _08292_/B _08292_/C _08292_/D VGND VGND VPWR VPWR _08292_/Y sky130_fd_sc_hd__nand4_2
X_07312_ _10338_/Q _05126_/Y input110/X _05112_/A _07311_/X VGND VGND VPWR VPWR _07317_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07243_ _07243_/A _07243_/B _07243_/C _07243_/D VGND VGND VPWR VPWR _07288_/B sky130_fd_sc_hd__and4_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07174_ _10125_/Q _05073_/Y input26/X _05129_/A VGND VGND VPWR VPWR _07174_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06125_ _10028_/Q _06123_/X _09545_/A1 _06124_/Y VGND VGND VPWR VPWR _10028_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06056_ _06056_/A VGND VGND VPWR VPWR _06057_/A sky130_fd_sc_hd__inv_2
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05007_ _06538_/A _05090_/A VGND VGND VPWR VPWR _05009_/A sky130_fd_sc_hd__or2_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09815_ _10353_/CLK _09815_/D repeater403/X VGND VGND VPWR VPWR _09815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09746_ _09752_/CLK _09746_/D VGND VGND VPWR VPWR _09746_/Q sky130_fd_sc_hd__dfxtp_1
X_06958_ _06956_/Y _05865_/B _06957_/Y _04871_/B VGND VGND VPWR VPWR _06958_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05909_ _05909_/A VGND VGND VPWR VPWR _05910_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09677_ split1/X _05677_/B _09677_/S VGND VGND VPWR VPWR _09677_/X sky130_fd_sc_hd__mux2_1
X_08628_ _08766_/B _08858_/A VGND VGND VPWR VPWR _09297_/B sky130_fd_sc_hd__nor2_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _06887_/Y _06339_/B _06888_/Y _06360_/B VGND VGND VPWR VPWR _06889_/X sky130_fd_sc_hd__o22a_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08552_/A _09006_/A _09155_/A _09006_/B VGND VGND VPWR VPWR _08559_/X sky130_fd_sc_hd__a211o_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10452_ _10486_/CLK _10452_/D _05034_/A VGND VGND VPWR VPWR _10452_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10383_ _04811_/A1 _10383_/D _05503_/X VGND VGND VPWR VPWR _10383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07930_ _07212_/Y _07818_/X _07929_/Y _07819_/X VGND VGND VPWR VPWR _07930_/X sky130_fd_sc_hd__o22a_1
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07861_ _10097_/Q VGND VGND VPWR VPWR _07861_/Y sky130_fd_sc_hd__inv_2
X_07792_ _07792_/A VGND VGND VPWR VPWR _07792_/X sky130_fd_sc_hd__clkbuf_2
X_06812_ _07823_/A _06267_/B _06811_/Y _05852_/B VGND VGND VPWR VPWR _06812_/X sky130_fd_sc_hd__o22a_1
X_09600_ _08218_/Y _10335_/Q _09700_/S VGND VGND VPWR VPWR _09600_/X sky130_fd_sc_hd__mux2_1
X_09531_ _09531_/A VGND VGND VPWR VPWR _09535_/B sky130_fd_sc_hd__inv_2
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06743_ _09981_/Q VGND VGND VPWR VPWR _07854_/A sky130_fd_sc_hd__inv_2
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06674_ _06674_/A VGND VGND VPWR VPWR _06674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09462_ _09462_/A VGND VGND VPWR VPWR _09462_/X sky130_fd_sc_hd__clkbuf_1
X_08413_ _08485_/A _08492_/B _08412_/Y _08492_/C _06464_/X VGND VGND VPWR VPWR _08913_/A
+ sky130_fd_sc_hd__a32o_1
X_09393_ _09393_/A _09393_/B _09393_/C VGND VGND VPWR VPWR _09435_/A sky130_fd_sc_hd__or3_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05625_ _06337_/A _05651_/B _05625_/C VGND VGND VPWR VPWR _05626_/A sky130_fd_sc_hd__or3_2
XFILLER_149_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05556_ _10362_/Q _05551_/X _09579_/X _05553_/X VGND VGND VPWR VPWR _10362_/D sky130_fd_sc_hd__a22o_1
X_08344_ _09805_/Q _08344_/B VGND VGND VPWR VPWR _08344_/Y sky130_fd_sc_hd__nand2_1
X_05487_ _08354_/A _08354_/B _09535_/A VGND VGND VPWR VPWR _05493_/B sky130_fd_sc_hd__a21oi_1
XFILLER_137_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08275_ _07206_/Y _08173_/X _07284_/Y _08174_/X VGND VGND VPWR VPWR _08275_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07226_ _10169_/Q VGND VGND VPWR VPWR _07226_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07157_ _07157_/A _07157_/B _07157_/C _07157_/D VGND VGND VPWR VPWR _07157_/X sky130_fd_sc_hd__and4_4
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06108_ _06108_/A _06108_/B VGND VGND VPWR VPWR _06110_/A sky130_fd_sc_hd__or2_2
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07088_ _07957_/A _06280_/B _09477_/A _06313_/B _07087_/X VGND VGND VPWR VPWR _07089_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06039_ _06039_/A VGND VGND VPWR VPWR _06039_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09729_ _10295_/Q _09511_/A VGND VGND VPWR VPWR _09729_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10504_ _10504_/CLK _10504_/D repeater402/X VGND VGND VPWR VPWR _10504_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10435_ _10478_/CLK _10435_/D _05034_/A VGND VGND VPWR VPWR _10435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10366_ _10366_/CLK _10366_/D repeater407/X VGND VGND VPWR VPWR _10366_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10297_ _10406_/CLK _10297_/D _05674_/X VGND VGND VPWR VPWR _10297_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater408 repeater409/X VGND VGND VPWR VPWR _05034_/A sky130_fd_sc_hd__buf_12
XFILLER_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ _05588_/A VGND VGND VPWR VPWR _05411_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ _06390_/A VGND VGND VPWR VPWR _06390_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05341_ _05337_/Y _06166_/A _05339_/Y _05473_/A VGND VGND VPWR VPWR _05341_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05272_ _05286_/B _05329_/A VGND VGND VPWR VPWR _05895_/A sky130_fd_sc_hd__or2_4
X_08060_ _08179_/A VGND VGND VPWR VPWR _08060_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07011_ _10205_/Q VGND VGND VPWR VPWR _07011_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08962_ _08962_/A _09357_/B VGND VGND VPWR VPWR _08964_/A sky130_fd_sc_hd__or2_1
X_08893_ _09233_/A _09295_/B _09295_/C VGND VGND VPWR VPWR _08908_/B sky130_fd_sc_hd__or3_1
XFILLER_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07913_ _10099_/Q VGND VGND VPWR VPWR _07913_/Y sky130_fd_sc_hd__inv_2
X_07844_ _06730_/Y _07755_/X _06709_/Y _07802_/X VGND VGND VPWR VPWR _07844_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07775_ _07775_/A _07775_/B _07775_/C _07775_/D VGND VGND VPWR VPWR _07776_/C sky130_fd_sc_hd__and4_1
X_04987_ _10454_/Q _04980_/X _09658_/A1 _04982_/X VGND VGND VPWR VPWR _10454_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09514_ _09514_/A VGND VGND VPWR VPWR _09514_/X sky130_fd_sc_hd__clkbuf_1
X_06726_ _06724_/Y _06206_/B _06725_/Y _05576_/B VGND VGND VPWR VPWR _06726_/X sky130_fd_sc_hd__o22a_1
X_06657_ _06663_/A VGND VGND VPWR VPWR _06658_/A sky130_fd_sc_hd__clkbuf_1
X_09445_ _09445_/A VGND VGND VPWR VPWR _09445_/Y sky130_fd_sc_hd__inv_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05608_ _10335_/Q _05604_/X _09580_/X _05606_/X VGND VGND VPWR VPWR _10335_/D sky130_fd_sc_hd__a22o_1
X_09376_ _09376_/A VGND VGND VPWR VPWR _09376_/X sky130_fd_sc_hd__clkbuf_1
X_06588_ _06588_/A VGND VGND VPWR VPWR _06588_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08327_ _08327_/A _08327_/B _08327_/C _08327_/D VGND VGND VPWR VPWR _08328_/D sky130_fd_sc_hd__and4_1
X_05539_ _10370_/Q _05530_/A _09659_/A1 _05531_/A VGND VGND VPWR VPWR _10370_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08258_ _07337_/Y _08219_/X _07333_/Y _08220_/X _08257_/X VGND VGND VPWR VPWR _08274_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07209_ _10255_/Q VGND VGND VPWR VPWR _07209_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08189_ _08189_/A VGND VGND VPWR VPWR _08189_/X sky130_fd_sc_hd__clkbuf_2
X_10220_ _10224_/CLK _10220_/D repeater405/X VGND VGND VPWR VPWR _10220_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10151_ _10257_/CLK _10151_/D repeater407/X VGND VGND VPWR VPWR _10151_/Q sky130_fd_sc_hd__dfstp_1
Xoutput280 _09706_/Z VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput291 _07498_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_2
X_10082_ _10374_/CLK _10082_/D hold41/A VGND VGND VPWR VPWR _10082_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10418_ _04807_/A1 _10418_/D _05394_/X VGND VGND VPWR VPWR _10418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10349_ _10349_/CLK _10349_/D repeater404/X VGND VGND VPWR VPWR _10349_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04910_ _05118_/B VGND VGND VPWR VPWR _05286_/A sky130_fd_sc_hd__clkbuf_4
X_05890_ _10171_/Q _05884_/X _09547_/A1 _05886_/X VGND VGND VPWR VPWR _10171_/D sky130_fd_sc_hd__a22o_1
X_04841_ _09663_/X VGND VGND VPWR VPWR _05213_/A sky130_fd_sc_hd__inv_2
X_07560_ _07646_/A _07610_/A _07589_/A _07583_/A VGND VGND VPWR VPWR _07567_/C sky130_fd_sc_hd__and4_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06511_ _09844_/Q _06504_/X _09550_/A0 _06506_/X VGND VGND VPWR VPWR _09844_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09230_ _08753_/C _08753_/B _09229_/Y _08700_/B VGND VGND VPWR VPWR _09235_/B sky130_fd_sc_hd__a31o_1
X_07491_ _10298_/Q _07492_/B VGND VGND VPWR VPWR _07491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_7_0_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_7_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
X_06442_ _06442_/A VGND VGND VPWR VPWR _06442_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09161_ _09377_/A _09161_/B _09161_/C _09319_/C VGND VGND VPWR VPWR _09163_/A sky130_fd_sc_hd__or4_1
X_06373_ _06390_/A VGND VGND VPWR VPWR _06417_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09092_ _09092_/A _09092_/B VGND VGND VPWR VPWR _09344_/B sky130_fd_sc_hd__or2_2
X_08112_ _07252_/Y _08088_/X _07200_/Y _08089_/X VGND VGND VPWR VPWR _08112_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05324_ _10398_/Q VGND VGND VPWR VPWR _05324_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08043_ _08044_/A _08043_/B _10006_/Q VGND VGND VPWR VPWR _08211_/A sky130_fd_sc_hd__or3_4
XFILLER_174_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05255_ _05327_/A _05307_/B VGND VGND VPWR VPWR _06078_/A sky130_fd_sc_hd__or2_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05186_ _10227_/Q VGND VGND VPWR VPWR _05186_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _10364_/CLK _09994_/D repeater410/X VGND VGND VPWR VPWR _09994_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08945_ _08945_/A _09198_/B _09021_/B VGND VGND VPWR VPWR _08948_/A sky130_fd_sc_hd__or3_1
X_08876_ _09141_/B _08876_/B VGND VGND VPWR VPWR _08878_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07827_ _07827_/A VGND VGND VPWR VPWR _07827_/X sky130_fd_sc_hd__clkbuf_2
X_07758_ _07758_/A VGND VGND VPWR VPWR _07758_/X sky130_fd_sc_hd__buf_4
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06709_ _09967_/Q VGND VGND VPWR VPWR _06709_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07689_ _07221_/Y _07656_/X _07264_/Y _07657_/X _07688_/X VGND VGND VPWR VPWR _07694_/B
+ sky130_fd_sc_hd__o221a_1
X_09428_ _09428_/A _09428_/B _09428_/C _09428_/D VGND VGND VPWR VPWR _09441_/A sky130_fd_sc_hd__or4_2
XFILLER_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09359_ _09359_/A _09428_/C _09390_/C _09433_/C VGND VGND VPWR VPWR _09359_/Y sky130_fd_sc_hd__nor4_1
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _10513_/CLK _10203_/D _07492_/B VGND VGND VPWR VPWR _10203_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10134_ _10135_/CLK _10134_/D _07492_/B VGND VGND VPWR VPWR _10134_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10065_ _10224_/CLK _10065_/D repeater405/X VGND VGND VPWR VPWR _10065_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05040_ _05041_/A VGND VGND VPWR VPWR _05040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _10347_/Q VGND VGND VPWR VPWR _06991_/Y sky130_fd_sc_hd__inv_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08730_ _08736_/A _08855_/A VGND VGND VPWR VPWR _09327_/B sky130_fd_sc_hd__nor2_2
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05942_ _05942_/A VGND VGND VPWR VPWR _05943_/A sky130_fd_sc_hd__inv_2
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05873_ _05873_/A VGND VGND VPWR VPWR _05874_/B sky130_fd_sc_hd__clkbuf_2
X_08661_ _08661_/A VGND VGND VPWR VPWR _08662_/A sky130_fd_sc_hd__inv_2
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07612_ _07612_/A _07612_/B _07612_/C VGND VGND VPWR VPWR _07829_/A sky130_fd_sc_hd__or3_4
X_04824_ _05651_/A VGND VGND VPWR VPWR _06679_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08592_ _09311_/A _08592_/B VGND VGND VPWR VPWR _08592_/Y sky130_fd_sc_hd__nor2_1
X_07543_ _07983_/B _07627_/A _07659_/A _07645_/A VGND VGND VPWR VPWR _07567_/A sky130_fd_sc_hd__and4_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07474_ _07539_/A VGND VGND VPWR VPWR _07565_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06425_ _06390_/X _09617_/X _09650_/X _09883_/Q VGND VGND VPWR VPWR _09883_/D sky130_fd_sc_hd__o22a_1
X_09213_ _09309_/D _09311_/D _09369_/C _09212_/X VGND VGND VPWR VPWR _09217_/A sky130_fd_sc_hd__or4b_4
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09144_ _09144_/A _09144_/B VGND VGND VPWR VPWR _09195_/A sky130_fd_sc_hd__nand2_1
X_06356_ _09930_/Q _06352_/X _09576_/X _06353_/Y VGND VGND VPWR VPWR _09930_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06287_ _09969_/Q _06281_/X _09574_/X _06282_/Y VGND VGND VPWR VPWR _09969_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05307_ _05336_/A _05307_/B VGND VGND VPWR VPWR _05882_/A sky130_fd_sc_hd__or2_4
X_09075_ _09342_/B _09075_/B VGND VGND VPWR VPWR _09357_/C sky130_fd_sc_hd__or2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05238_ _05284_/B _05355_/B VGND VGND VPWR VPWR _06338_/A sky130_fd_sc_hd__or2_4
X_08026_ _08026_/A _10002_/Q _08046_/C _08038_/C VGND VGND VPWR VPWR _08194_/A sky130_fd_sc_hd__or4_4
XFILLER_150_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05169_ input43/X _06697_/A input61/X _06844_/A VGND VGND VPWR VPWR _05169_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09977_ _10000_/CLK _09977_/D repeater405/X VGND VGND VPWR VPWR _09977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08928_ _08928_/A VGND VGND VPWR VPWR _09064_/B sky130_fd_sc_hd__inv_2
XFILLER_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08859_ _08859_/A _09420_/D VGND VGND VPWR VPWR _08861_/A sky130_fd_sc_hd__or2_1
XFILLER_55_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10409_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10117_ _10119_/CLK _10117_/D repeater402/X VGND VGND VPWR VPWR _10117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10048_ _10127_/CLK _10048_/D repeater409/X VGND VGND VPWR VPWR _10048_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06210_ _10001_/Q _06207_/X _09581_/X _06209_/X VGND VGND VPWR VPWR _10001_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07190_ _10135_/Q VGND VGND VPWR VPWR _07190_/Y sky130_fd_sc_hd__inv_2
X_06141_ _09776_/Q _07477_/C _09778_/Q VGND VGND VPWR VPWR _06142_/B sky130_fd_sc_hd__a21o_1
XFILLER_172_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06072_ _10060_/Q _06067_/X _09579_/X _06069_/X VGND VGND VPWR VPWR _10060_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09900_ _10268_/CLK _09900_/D repeater404/X VGND VGND VPWR VPWR _09900_/Q sky130_fd_sc_hd__dfrtp_1
X_05023_ _10435_/Q _05020_/X _09658_/A1 _05021_/Y VGND VGND VPWR VPWR _10435_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09831_ _10355_/CLK _09831_/D repeater406/X VGND VGND VPWR VPWR _09831_/Q sky130_fd_sc_hd__dfrtp_1
X_06974_ _09866_/Q VGND VGND VPWR VPWR _06974_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_86_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09762_ _09919_/CLK _09762_/D VGND VGND VPWR VPWR _09762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05925_ _10149_/Q _05919_/X _09536_/A3 _05920_/Y VGND VGND VPWR VPWR _10149_/D sky130_fd_sc_hd__a22o_1
X_08713_ _08717_/A _08836_/B VGND VGND VPWR VPWR _09118_/A sky130_fd_sc_hd__or2_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _09196_/X _09043_/X _09698_/S VGND VGND VPWR VPWR _09693_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08644_ _08644_/A _08814_/B VGND VGND VPWR VPWR _08668_/A sky130_fd_sc_hd__or2_4
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05856_ _10192_/Q _05853_/X _09581_/X _05855_/X VGND VGND VPWR VPWR _10192_/D sky130_fd_sc_hd__a22o_1
X_05787_ _05787_/A VGND VGND VPWR VPWR _05787_/Y sky130_fd_sc_hd__inv_2
X_04807_ _10267_/Q _04807_/A1 _10342_/Q VGND VGND VPWR VPWR _09708_/A sky130_fd_sc_hd__mux2_1
X_08575_ _08575_/A _08927_/B VGND VGND VPWR VPWR _09003_/A sky130_fd_sc_hd__or2_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07526_ _07749_/A VGND VGND VPWR VPWR _07527_/A sky130_fd_sc_hd__clkbuf_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07457_ _07030_/X _07451_/X _09738_/Q _07453_/X VGND VGND VPWR VPWR _09738_/D sky130_fd_sc_hd__o22a_2
X_07388_ _09903_/Q VGND VGND VPWR VPWR _07388_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06408_ _09899_/Q _06403_/X _09579_/X _06405_/X VGND VGND VPWR VPWR _09899_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06339_ _06481_/A _06339_/B VGND VGND VPWR VPWR _06341_/A sky130_fd_sc_hd__or2_2
X_09127_ _09263_/A _09099_/X _09123_/X _09126_/Y VGND VGND VPWR VPWR _09127_/X sky130_fd_sc_hd__o211a_1
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09058_ _09058_/A _09058_/B _09058_/C VGND VGND VPWR VPWR _09058_/X sky130_fd_sc_hd__and3_1
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08009_ _08032_/A _08032_/B _10006_/Q VGND VGND VPWR VPWR _08178_/A sky130_fd_sc_hd__or3_4
XFILLER_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput180 wb_dat_i[23] VGND VGND VPWR VPWR _08371_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput191 wb_dat_i[4] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05710_ _10275_/Q _05701_/A _09659_/X _05702_/A VGND VGND VPWR VPWR _10275_/D sky130_fd_sc_hd__o22a_1
X_06690_ _10466_/Q _06853_/B input42/X _06770_/A VGND VGND VPWR VPWR _06690_/X sky130_fd_sc_hd__a22o_1
X_05641_ _05641_/A VGND VGND VPWR VPWR _05642_/A sky130_fd_sc_hd__inv_2
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08360_ _09790_/Q input182/X _09789_/Q input196/X _08359_/X VGND VGND VPWR VPWR _08360_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05572_ _10353_/Q _05568_/X _09576_/X _05569_/Y VGND VGND VPWR VPWR _10353_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07311_ input129/X _05118_/Y _10438_/Q _05091_/A VGND VGND VPWR VPWR _07311_/X sky130_fd_sc_hd__a22o_1
X_08291_ _08291_/A _08291_/B _08291_/C _08291_/D VGND VGND VPWR VPWR _08292_/D sky130_fd_sc_hd__and4_2
X_07242_ _07237_/Y _06053_/A _07238_/Y _06122_/B _07241_/X VGND VGND VPWR VPWR _07243_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_176_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07173_ _10109_/Q _05094_/Y _10453_/Q _05089_/A _07172_/X VGND VGND VPWR VPWR _07181_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06124_ _06124_/A VGND VGND VPWR VPWR _06124_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06055_ _06056_/A VGND VGND VPWR VPWR _06055_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05006_ _05155_/A _05205_/A VGND VGND VPWR VPWR _05090_/A sky130_fd_sc_hd__or2_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09814_ _10406_/CLK _09814_/D _06560_/X VGND VGND VPWR VPWR _09814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09745_ _09752_/CLK _09745_/D VGND VGND VPWR VPWR _09745_/Q sky130_fd_sc_hd__dfxtp_1
X_06957_ _10500_/Q VGND VGND VPWR VPWR _06957_/Y sky130_fd_sc_hd__inv_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _09925_/Q VGND VGND VPWR VPWR _06888_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09676_ _09675_/X _10392_/Q _10299_/Q VGND VGND VPWR VPWR _09676_/X sky130_fd_sc_hd__mux2_4
X_05908_ _06327_/A VGND VGND VPWR VPWR _05993_/A sky130_fd_sc_hd__buf_4
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05839_ _05896_/A _05839_/B VGND VGND VPWR VPWR _05841_/A sky130_fd_sc_hd__or2_2
X_08627_ _08851_/A VGND VGND VPWR VPWR _08858_/A sky130_fd_sc_hd__buf_4
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08558_ _08563_/A _09006_/B VGND VGND VPWR VPWR _09149_/A sky130_fd_sc_hd__or2_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07509_ _09991_/Q _09990_/Q VGND VGND VPWR VPWR _07597_/C sky130_fd_sc_hd__or2_1
X_08489_ _09155_/A VGND VGND VPWR VPWR _08490_/A sky130_fd_sc_hd__inv_2
XFILLER_168_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10451_ _10486_/CLK _10451_/D repeater409/X VGND VGND VPWR VPWR _10451_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_182_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10382_ _10382_/CLK _10382_/D _05507_/X VGND VGND VPWR VPWR _10382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07860_ _07860_/A _07860_/B _07860_/C VGND VGND VPWR VPWR _07860_/Y sky130_fd_sc_hd__nand3_2
XFILLER_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07791_ _06790_/Y _07787_/X _06783_/Y _07788_/X _07790_/X VGND VGND VPWR VPWR _07810_/A
+ sky130_fd_sc_hd__o221a_1
X_06811_ _10191_/Q VGND VGND VPWR VPWR _06811_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06742_ _09848_/Q VGND VGND VPWR VPWR _06742_/Y sky130_fd_sc_hd__inv_2
X_09530_ _09530_/A VGND VGND VPWR VPWR _09530_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09461_ _09461_/A VGND VGND VPWR VPWR _09462_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06673_ _06677_/A VGND VGND VPWR VPWR _06674_/A sky130_fd_sc_hd__clkbuf_1
X_08412_ _08412_/A _08412_/B VGND VGND VPWR VPWR _08412_/Y sky130_fd_sc_hd__nand2_1
X_09392_ _09428_/D _09443_/D _09392_/C _09432_/A VGND VGND VPWR VPWR _09392_/Y sky130_fd_sc_hd__nor4_1
X_05624_ split1/X VGND VGND VPWR VPWR _05651_/B sky130_fd_sc_hd__clkinv_4
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05555_ _10363_/Q _05551_/X _09580_/X _05553_/X VGND VGND VPWR VPWR _10363_/D sky130_fd_sc_hd__a22o_1
X_08343_ _08343_/A VGND VGND VPWR VPWR _08344_/B sky130_fd_sc_hd__inv_2
X_08274_ _08274_/A _08274_/B _08274_/C _08274_/D VGND VGND VPWR VPWR _08274_/Y sky130_fd_sc_hd__nand4_2
X_05486_ _09790_/Q VGND VGND VPWR VPWR _09535_/A sky130_fd_sc_hd__inv_2
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07225_ _10187_/Q VGND VGND VPWR VPWR _07225_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07156_ _07156_/A _07156_/B _07156_/C _07156_/D VGND VGND VPWR VPWR _07157_/D sky130_fd_sc_hd__and4_1
X_07087_ _07085_/Y _05874_/B _07086_/Y _06251_/B VGND VGND VPWR VPWR _07087_/X sky130_fd_sc_hd__o22a_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06107_ _10037_/Q _06098_/A _09659_/A1 _06099_/A VGND VGND VPWR VPWR _10037_/D sky130_fd_sc_hd__a22o_1
XFILLER_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06038_ _06039_/A VGND VGND VPWR VPWR _06038_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09728_ _10294_/Q _09509_/A VGND VGND VPWR VPWR _09728_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07989_ _08010_/C _07989_/B _10006_/Q VGND VGND VPWR VPWR _09700_/S sky130_fd_sc_hd__nor3_4
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _10316_/Q _09659_/A1 _09679_/S VGND VGND VPWR VPWR _09659_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10503_ _10504_/CLK _10503_/D repeater404/X VGND VGND VPWR VPWR _10503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10434_ _10483_/CLK _10434_/D _05034_/A VGND VGND VPWR VPWR _10434_/Q sky130_fd_sc_hd__dfstp_2
X_10365_ _10369_/CLK _10365_/D repeater407/X VGND VGND VPWR VPWR _10365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10296_/CLK _10296_/D repeater402/X VGND VGND VPWR VPWR _10296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater409 _07492_/B VGND VGND VPWR VPWR repeater409/X sky130_fd_sc_hd__buf_12
XFILLER_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05340_ _05340_/A _05359_/B VGND VGND VPWR VPWR _05473_/A sky130_fd_sc_hd__or2_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05271_ _10159_/Q VGND VGND VPWR VPWR _05271_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07010_ _09845_/Q VGND VGND VPWR VPWR _07010_/Y sky130_fd_sc_hd__clkinv_2
X_08961_ _09029_/A _08961_/B VGND VGND VPWR VPWR _09357_/B sky130_fd_sc_hd__nor2_1
X_08892_ _09052_/A _09052_/B _08891_/X VGND VGND VPWR VPWR _09295_/C sky130_fd_sc_hd__o21ai_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07912_ _07912_/A _07912_/B _07912_/C VGND VGND VPWR VPWR _07912_/Y sky130_fd_sc_hd__nand3_2
Xclkbuf_opt_3_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07843_ _10140_/Q VGND VGND VPWR VPWR _07843_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07774_ _06893_/A _07665_/X _07772_/Y _07666_/X _07773_/X VGND VGND VPWR VPWR _07775_/D
+ sky130_fd_sc_hd__o221a_1
X_04986_ _10455_/Q _04980_/X _09545_/A1 _04982_/X VGND VGND VPWR VPWR _10455_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09513_ _09513_/A VGND VGND VPWR VPWR _09514_/A sky130_fd_sc_hd__clkbuf_1
X_06725_ _10350_/Q VGND VGND VPWR VPWR _06725_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06656_ _06656_/A VGND VGND VPWR VPWR _06656_/X sky130_fd_sc_hd__clkbuf_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09444_ _09444_/A VGND VGND VPWR VPWR _09444_/Y sky130_fd_sc_hd__inv_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05607_ _10336_/Q _05604_/X _09581_/X _05606_/X VGND VGND VPWR VPWR _10336_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09375_ _09408_/C _09439_/C _09375_/C _09433_/A VGND VGND VPWR VPWR _09376_/A sky130_fd_sc_hd__or4_1
X_06587_ _06591_/A VGND VGND VPWR VPWR _06588_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08326_ _06982_/Y _08211_/A _07983_/A _08212_/A _08325_/X VGND VGND VPWR VPWR _08327_/D
+ sky130_fd_sc_hd__o221a_1
X_05538_ _10371_/Q _05530_/A _09661_/A1 _05531_/A VGND VGND VPWR VPWR _10371_/D sky130_fd_sc_hd__a22o_1
XFILLER_165_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05469_ _09693_/X _05450_/A _10392_/Q _05493_/D VGND VGND VPWR VPWR _10392_/D sky130_fd_sc_hd__a22o_1
X_08257_ _07339_/Y _08173_/X _07382_/Y _08174_/X VGND VGND VPWR VPWR _08257_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07208_ _10490_/Q VGND VGND VPWR VPWR _07208_/Y sky130_fd_sc_hd__clkinv_4
X_08188_ _08188_/A VGND VGND VPWR VPWR _08188_/X sky130_fd_sc_hd__clkbuf_2
X_07139_ _09923_/Q VGND VGND VPWR VPWR _09473_/A sky130_fd_sc_hd__inv_4
XFILLER_133_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput270 _09731_/Z VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_2
X_10150_ _10257_/CLK _10150_/D repeater407/X VGND VGND VPWR VPWR _10150_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput281 _09707_/Z VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput292 _07498_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_2
X_10081_ _10135_/CLK _10081_/D _07492_/B VGND VGND VPWR VPWR _10081_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10417_ _04807_/A1 _10417_/D _05401_/X VGND VGND VPWR VPWR _10417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10348_ _10350_/CLK _10348_/D repeater404/X VGND VGND VPWR VPWR _10348_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10279_ _10364_/CLK _10279_/D repeater410/X VGND VGND VPWR VPWR _10279_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04840_ _04991_/A _09668_/X _09674_/X _04963_/B VGND VGND VPWR VPWR _05118_/B sky130_fd_sc_hd__or4_4
XFILLER_80_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06510_ _09845_/Q _06504_/X _09547_/A1 _06506_/X VGND VGND VPWR VPWR _09845_/D sky130_fd_sc_hd__a22o_1
X_07490_ _09773_/Q _05376_/X _09772_/Q _07489_/X VGND VGND VPWR VPWR _09772_/D sky130_fd_sc_hd__a22o_1
X_06441_ _06441_/A VGND VGND VPWR VPWR _06442_/A sky130_fd_sc_hd__inv_2
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09160_ _08934_/A _09010_/X _08661_/A _08678_/X VGND VGND VPWR VPWR _09319_/C sky130_fd_sc_hd__o22ai_1
X_06372_ _09650_/X VGND VGND VPWR VPWR _06390_/A sky130_fd_sc_hd__inv_2
X_09091_ _09362_/C _09091_/B VGND VGND VPWR VPWR _09144_/A sky130_fd_sc_hd__or2_1
X_08111_ _07197_/Y _08080_/X _07251_/Y _08081_/X _08110_/X VGND VGND VPWR VPWR _08116_/B
+ sky130_fd_sc_hd__o221a_1
X_05323_ _05357_/A _05355_/B VGND VGND VPWR VPWR _06359_/A sky130_fd_sc_hd__or2_2
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08042_ _05328_/Y _08205_/A _05263_/Y _08206_/A _08041_/X VGND VGND VPWR VPWR _08049_/C
+ sky130_fd_sc_hd__o221a_1
X_05254_ _10050_/Q VGND VGND VPWR VPWR _05254_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05185_ _05286_/A _05311_/B VGND VGND VPWR VPWR _05927_/A sky130_fd_sc_hd__or2_4
XFILLER_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09993_ _10006_/CLK _09993_/D repeater407/X VGND VGND VPWR VPWR _09993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08944_ _09024_/A _08961_/B VGND VGND VPWR VPWR _09021_/B sky130_fd_sc_hd__nor2_1
X_08875_ _09363_/A _09273_/A _09275_/A _08874_/Y VGND VGND VPWR VPWR _08876_/B sky130_fd_sc_hd__or4b_1
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07826_ _10061_/Q VGND VGND VPWR VPWR _07826_/Y sky130_fd_sc_hd__inv_2
X_04969_ _10466_/Q _04966_/X _09581_/X _04968_/X VGND VGND VPWR VPWR _10466_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07757_ _07754_/Y _07639_/X _06851_/Y _07641_/X _07756_/X VGND VGND VPWR VPWR _07761_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06708_ _06708_/A _06708_/B VGND VGND VPWR VPWR _06708_/X sky130_fd_sc_hd__or2_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07688_ _07201_/Y _07658_/X _07687_/Y _07659_/X VGND VGND VPWR VPWR _07688_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06639_ _09795_/Q _06636_/X _09550_/A0 _06637_/Y VGND VGND VPWR VPWR _09795_/D sky130_fd_sc_hd__a22o_1
X_09427_ _09427_/A _09427_/B _09427_/C VGND VGND VPWR VPWR _09428_/B sky130_fd_sc_hd__or3_1
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09358_ _09358_/A _09358_/B VGND VGND VPWR VPWR _09390_/C sky130_fd_sc_hd__or2_1
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08309_ _08309_/A _08309_/B _08309_/C _08309_/D VGND VGND VPWR VPWR _08310_/D sky130_fd_sc_hd__and4_1
X_09289_ _09289_/A _09289_/B _09289_/C VGND VGND VPWR VPWR _09387_/C sky130_fd_sc_hd__or3_1
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ _10513_/CLK _10202_/D _07492_/B VGND VGND VPWR VPWR _10202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10133_ _10135_/CLK _10133_/D _07492_/B VGND VGND VPWR VPWR _10133_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10064_ _10224_/CLK _10064_/D repeater405/X VGND VGND VPWR VPWR _10064_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _10355_/Q VGND VGND VPWR VPWR _06990_/Y sky130_fd_sc_hd__inv_2
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _05942_/A VGND VGND VPWR VPWR _05941_/X sky130_fd_sc_hd__clkbuf_2
X_05872_ _10180_/Q _05866_/X _09536_/A3 _05867_/Y VGND VGND VPWR VPWR _10180_/D sky130_fd_sc_hd__a22o_1
X_08660_ _08849_/B VGND VGND VPWR VPWR _09263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07611_ _07611_/A _07612_/B _07612_/C VGND VGND VPWR VPWR _07828_/A sky130_fd_sc_hd__or3_4
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04823_ _09678_/X VGND VGND VPWR VPWR _05651_/A sky130_fd_sc_hd__inv_2
X_08591_ _09171_/A _08591_/B VGND VGND VPWR VPWR _08592_/B sky130_fd_sc_hd__or2_1
X_07542_ _07805_/A VGND VGND VPWR VPWR _07645_/A sky130_fd_sc_hd__buf_2
X_07473_ _07473_/A _09992_/Q VGND VGND VPWR VPWR _07539_/A sky130_fd_sc_hd__or2_1
XFILLER_167_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09212_ _09209_/X _09212_/B _09212_/C VGND VGND VPWR VPWR _09212_/X sky130_fd_sc_hd__and3b_1
X_06424_ _06390_/X _09619_/X _09650_/X _09884_/Q VGND VGND VPWR VPWR _09884_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06355_ _09931_/Q _06352_/X _09550_/A0 _06353_/Y VGND VGND VPWR VPWR _09931_/D sky130_fd_sc_hd__a22o_1
X_09143_ _09348_/B _09143_/B VGND VGND VPWR VPWR _09144_/B sky130_fd_sc_hd__or2_1
X_05306_ _10167_/Q VGND VGND VPWR VPWR _05308_/A sky130_fd_sc_hd__clkinv_4
X_06286_ _09970_/Q _06281_/X hold46/X _06282_/Y VGND VGND VPWR VPWR _09970_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09074_ _09074_/A _09289_/C _09387_/A _09290_/C VGND VGND VPWR VPWR _09078_/A sky130_fd_sc_hd__or4_2
X_05237_ _09933_/Q VGND VGND VPWR VPWR _05237_/Y sky130_fd_sc_hd__inv_2
X_08025_ _08038_/A _08044_/B _10006_/Q VGND VGND VPWR VPWR _08193_/A sky130_fd_sc_hd__or3_4
X_05168_ _05689_/B VGND VGND VPWR VPWR _06844_/A sky130_fd_sc_hd__inv_2
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09976_ _10000_/CLK _09976_/D repeater405/X VGND VGND VPWR VPWR _09976_/Q sky130_fd_sc_hd__dfrtp_1
X_05099_ _05625_/C VGND VGND VPWR VPWR _06693_/A sky130_fd_sc_hd__clkinv_2
X_08927_ _08927_/A _08927_/B VGND VGND VPWR VPWR _08928_/A sky130_fd_sc_hd__or2_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08858_ _08858_/A _08862_/A VGND VGND VPWR VPWR _09420_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07809_ _06797_/Y _07805_/X _06798_/Y _07758_/X _07808_/X VGND VGND VPWR VPWR _07810_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08789_ _08794_/A _08789_/B VGND VGND VPWR VPWR _08908_/A sky130_fd_sc_hd__or2_1
XFILLER_187_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10116_ _10119_/CLK _10116_/D repeater403/X VGND VGND VPWR VPWR _10116_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10047_ _10127_/CLK _10047_/D repeater409/X VGND VGND VPWR VPWR _10047_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06140_ _06140_/A _06140_/B _10021_/Q _10020_/Q VGND VGND VPWR VPWR _07477_/C sky130_fd_sc_hd__or4_1
XANTENNA_0 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06071_ _10061_/Q _06067_/X _09580_/X _06069_/X VGND VGND VPWR VPWR _10061_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05022_ _10436_/Q _05020_/X _09545_/A1 _05021_/Y VGND VGND VPWR VPWR _10436_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09830_ _10354_/CLK _09830_/D repeater406/X VGND VGND VPWR VPWR _09830_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_112_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06973_ _09858_/Q VGND VGND VPWR VPWR _06973_/Y sky130_fd_sc_hd__clkinv_4
X_09761_ _09919_/CLK _09761_/D VGND VGND VPWR VPWR _09761_/Q sky130_fd_sc_hd__dfxtp_1
X_05924_ _10150_/Q _05919_/X _06684_/B1 _05920_/Y VGND VGND VPWR VPWR _10150_/D sky130_fd_sc_hd__a22o_1
X_08712_ _09095_/A _08674_/X _08684_/A _08831_/B _08711_/X VGND VGND VPWR VPWR _08712_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09692_ _08994_/Y _08611_/X _09698_/S VGND VGND VPWR VPWR _09692_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08643_ _08643_/A _08895_/A VGND VGND VPWR VPWR _08814_/B sky130_fd_sc_hd__or2_1
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05855_ _05855_/A VGND VGND VPWR VPWR _05855_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05786_ _05787_/A VGND VGND VPWR VPWR _05786_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08574_ _08529_/A _08925_/A _08554_/Y _08560_/X _08573_/X VGND VGND VPWR VPWR _08574_/X
+ sky130_fd_sc_hd__o2111a_1
X_04806_ _10268_/Q input58/X _10342_/Q VGND VGND VPWR VPWR _09709_/A sky130_fd_sc_hd__mux2_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _07601_/B _07549_/B VGND VGND VPWR VPWR _07749_/A sky130_fd_sc_hd__or2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07456_ _06906_/X _07451_/X _09739_/Q _07453_/X VGND VGND VPWR VPWR _09739_/D sky130_fd_sc_hd__o22a_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06407_ _09900_/Q _06403_/X _09580_/X _06405_/X VGND VGND VPWR VPWR _09900_/D sky130_fd_sc_hd__a22o_1
X_07387_ _09834_/Q VGND VGND VPWR VPWR _07387_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06338_ _06338_/A VGND VGND VPWR VPWR _06339_/B sky130_fd_sc_hd__clkbuf_4
X_09126_ _09398_/A VGND VGND VPWR VPWR _09126_/Y sky130_fd_sc_hd__inv_2
X_09057_ _09057_/A _09057_/B _09352_/C VGND VGND VPWR VPWR _09058_/C sky130_fd_sc_hd__or3_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06269_ _06269_/A VGND VGND VPWR VPWR _06270_/A sky130_fd_sc_hd__inv_2
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08008_ _08037_/B _08019_/B _10006_/Q VGND VGND VPWR VPWR _08177_/A sky130_fd_sc_hd__or3_4
XFILLER_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ _10288_/CLK _09959_/D repeater406/X VGND VGND VPWR VPWR _09959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput181 wb_dat_i[24] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__clkbuf_1
Xinput170 wb_dat_i[14] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__clkbuf_1
Xinput192 wb_dat_i[5] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05640_ _05641_/A VGND VGND VPWR VPWR _05640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05571_ _10354_/Q _05568_/X _09577_/X _05569_/Y VGND VGND VPWR VPWR _10354_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07310_ _10510_/Q _04835_/Y _10134_/Q _06705_/Y _07309_/X VGND VGND VPWR VPWR _07317_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08290_ _07182_/Y _08211_/X _07932_/A _08212_/X _08289_/X VGND VGND VPWR VPWR _08291_/D
+ sky130_fd_sc_hd__o221a_1
X_07241_ _07239_/Y _05567_/B _07240_/Y _05874_/B VGND VGND VPWR VPWR _07241_/X sky130_fd_sc_hd__o22a_1
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07172_ _10512_/Q _04822_/Y input37/X _06770_/A VGND VGND VPWR VPWR _07172_/X sky130_fd_sc_hd__a22o_1
X_06123_ _06124_/A VGND VGND VPWR VPWR _06123_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06054_ _06108_/A _06893_/B VGND VGND VPWR VPWR _06056_/A sky130_fd_sc_hd__or2_2
X_05005_ _09670_/X _09668_/X _05005_/C _09676_/X VGND VGND VPWR VPWR _05205_/A sky130_fd_sc_hd__or4_2
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09813_ _10406_/CLK _09813_/D _06569_/X VGND VGND VPWR VPWR _09813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09744_ _09752_/CLK _09744_/D VGND VGND VPWR VPWR _09744_/Q sky130_fd_sc_hd__dfxtp_1
X_06956_ _10184_/Q VGND VGND VPWR VPWR _06956_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05907_ _10159_/Q _05898_/A _09574_/X _05899_/A VGND VGND VPWR VPWR _10159_/D sky130_fd_sc_hd__a22o_1
X_06887_ _09938_/Q VGND VGND VPWR VPWR _06887_/Y sky130_fd_sc_hd__inv_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _09800_/Q _09799_/Q _09773_/Q VGND VGND VPWR VPWR _09675_/X sky130_fd_sc_hd__mux2_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05838_ _05838_/A VGND VGND VPWR VPWR _05839_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08626_ _08837_/A VGND VGND VPWR VPWR _08851_/A sky130_fd_sc_hd__buf_4
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05769_ _10241_/Q _05763_/X _09547_/A1 _05765_/X VGND VGND VPWR VPWR _10241_/D sky130_fd_sc_hd__a22o_1
X_08557_ _08921_/B VGND VGND VPWR VPWR _09006_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10355_/CLK sky130_fd_sc_hd__clkbuf_16
X_08488_ _08582_/A VGND VGND VPWR VPWR _09155_/A sky130_fd_sc_hd__clkbuf_4
X_07508_ _07608_/A VGND VGND VPWR VPWR _07601_/A sky130_fd_sc_hd__clkbuf_2
X_07439_ _07440_/A VGND VGND VPWR VPWR _07439_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10450_ _10487_/CLK _10450_/D repeater409/X VGND VGND VPWR VPWR _10450_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09109_ _09109_/A _09109_/B VGND VGND VPWR VPWR _09109_/X sky130_fd_sc_hd__or2_1
XFILLER_184_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10381_ _10382_/CLK _10381_/D _05511_/X VGND VGND VPWR VPWR _10381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_opt_9_0_csclk/X VGND VGND VPWR VPWR _10490_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07790_ _06809_/Y _07749_/X _06785_/Y _07789_/X VGND VGND VPWR VPWR _07790_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06810_ _09980_/Q VGND VGND VPWR VPWR _07823_/A sky130_fd_sc_hd__inv_2
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06741_ _10405_/Q VGND VGND VPWR VPWR _06741_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09460_ _09460_/A VGND VGND VPWR VPWR _09460_/X sky130_fd_sc_hd__clkbuf_1
X_08411_ _08913_/B VGND VGND VPWR VPWR _08644_/A sky130_fd_sc_hd__inv_2
X_06672_ _06672_/A VGND VGND VPWR VPWR _06672_/X sky130_fd_sc_hd__clkbuf_1
X_09391_ _09433_/A _09432_/C _09433_/C _09435_/C VGND VGND VPWR VPWR _09392_/C sky130_fd_sc_hd__or4_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05623_ _05651_/A VGND VGND VPWR VPWR _06337_/A sky130_fd_sc_hd__buf_2
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05554_ _10364_/Q _05551_/X _09581_/X _05553_/X VGND VGND VPWR VPWR _10364_/D sky130_fd_sc_hd__a22o_1
X_08342_ _09804_/Q _08341_/B _08343_/A VGND VGND VPWR VPWR _08342_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05485_ _08353_/A _08354_/A _09532_/A VGND VGND VPWR VPWR _05493_/A sky130_fd_sc_hd__a21oi_1
X_08273_ _08273_/A _08273_/B _08273_/C _08273_/D VGND VGND VPWR VPWR _08274_/D sky130_fd_sc_hd__and4_2
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07224_ _07219_/Y _06312_/A _07220_/Y _05749_/B _07223_/X VGND VGND VPWR VPWR _07243_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07155_ _07150_/Y _05740_/B _07151_/Y _06430_/B _07154_/X VGND VGND VPWR VPWR _07156_/D
+ sky130_fd_sc_hd__o221a_1
X_07086_ _09986_/Q VGND VGND VPWR VPWR _07086_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06106_ _10038_/Q _06098_/A _09661_/A1 _06099_/A VGND VGND VPWR VPWR _10038_/D sky130_fd_sc_hd__a22o_1
X_06037_ _06087_/A _06037_/B VGND VGND VPWR VPWR _06039_/A sky130_fd_sc_hd__or2_1
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07988_ _07988_/A _07988_/B _07988_/C VGND VGND VPWR VPWR _07988_/Y sky130_fd_sc_hd__nand3_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09727_ _10293_/Q _09507_/A VGND VGND VPWR VPWR _09727_/Z sky130_fd_sc_hd__ebufn_1
X_06939_ _10028_/Q VGND VGND VPWR VPWR _06939_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09658_ _10319_/Q _09658_/A1 _09679_/S VGND VGND VPWR VPWR _09658_/X sky130_fd_sc_hd__mux2_1
X_09589_ _09574_/X _10300_/Q _09677_/S VGND VGND VPWR VPWR _09589_/X sky130_fd_sc_hd__mux2_1
X_08609_ _09363_/A _09273_/A _08609_/C VGND VGND VPWR VPWR _08610_/B sky130_fd_sc_hd__or3_1
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10502_ _10504_/CLK _10502_/D repeater404/X VGND VGND VPWR VPWR _10502_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10433_ _10483_/CLK _10433_/D _05034_/A VGND VGND VPWR VPWR _10433_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_128_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10364_ _10364_/CLK _10364_/D repeater410/X VGND VGND VPWR VPWR _10364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10295_ _10296_/CLK _10295_/D repeater402/X VGND VGND VPWR VPWR _10295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05270_ _05260_/Y _06635_/B _05263_/Y _05727_/A _05269_/X VGND VGND VPWR VPWR _05281_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08960_ _08960_/A _09075_/B VGND VGND VPWR VPWR _08962_/A sky130_fd_sc_hd__or2_1
X_08891_ _08571_/C _08890_/Y _08494_/A _08635_/Y VGND VGND VPWR VPWR _08891_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07911_ _07911_/A _07911_/B _07911_/C _07911_/D VGND VGND VPWR VPWR _07912_/C sky130_fd_sc_hd__and4_2
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07842_ _10036_/Q VGND VGND VPWR VPWR _07842_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09512_ _09512_/A VGND VGND VPWR VPWR _09512_/X sky130_fd_sc_hd__clkbuf_1
X_07773_ _06859_/Y _07667_/X _06870_/Y _07668_/X VGND VGND VPWR VPWR _07773_/X sky130_fd_sc_hd__o22a_1
X_04985_ _10456_/Q _04980_/X _09579_/X _04982_/X VGND VGND VPWR VPWR _10456_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06724_ _10001_/Q VGND VGND VPWR VPWR _06724_/Y sky130_fd_sc_hd__inv_2
X_06655_ _06655_/A VGND VGND VPWR VPWR _06656_/A sky130_fd_sc_hd__clkbuf_1
X_09443_ _09443_/A _09443_/B _09443_/C _09443_/D VGND VGND VPWR VPWR _09443_/X sky130_fd_sc_hd__or4_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09374_ _09374_/A _09374_/B _09374_/C _09373_/X VGND VGND VPWR VPWR _09375_/C sky130_fd_sc_hd__or4b_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05606_ _05606_/A VGND VGND VPWR VPWR _05606_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08325_ _06964_/Y _08213_/A _06975_/Y _08214_/A VGND VGND VPWR VPWR _08325_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06586_ _09770_/Q _09680_/S input58/X _09810_/Q _06585_/X VGND VGND VPWR VPWR _09810_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05537_ _10372_/Q _05530_/A _09660_/A1 _05531_/A VGND VGND VPWR VPWR _10372_/D sky130_fd_sc_hd__a22o_1
X_05468_ _05468_/A VGND VGND VPWR VPWR _05468_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08256_ _08256_/A _08256_/B _08256_/C _08256_/D VGND VGND VPWR VPWR _08256_/Y sky130_fd_sc_hd__nand4_2
X_08187_ _08187_/A VGND VGND VPWR VPWR _08187_/X sky130_fd_sc_hd__clkbuf_2
X_07207_ _09922_/Q VGND VGND VPWR VPWR _07207_/Y sky130_fd_sc_hd__inv_2
X_05399_ _10418_/Q _05396_/X _10417_/Q _05398_/X VGND VGND VPWR VPWR _10418_/D sky130_fd_sc_hd__a22o_1
X_07138_ _09944_/Q VGND VGND VPWR VPWR _07138_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 _09732_/Z VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput260 _09722_/Z VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_160_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07069_ _07067_/Y _05474_/B _09503_/A _05748_/A VGND VGND VPWR VPWR _07069_/X sky130_fd_sc_hd__o22a_1
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10080_ _10411_/CLK _10080_/D repeater407/X VGND VGND VPWR VPWR _10080_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput282 _09708_/Z VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_1
Xoutput293 _10440_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_2
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10416_ _04807_/A1 _10416_/D _05404_/X VGND VGND VPWR VPWR _10416_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10347_ _10350_/CLK _10347_/D repeater404/X VGND VGND VPWR VPWR _10347_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10278_ _10405_/CLK _10278_/D hold41/X VGND VGND VPWR VPWR _10278_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06440_ _06441_/A VGND VGND VPWR VPWR _06440_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ _09920_/Q _06362_/A _09659_/A1 _06363_/A VGND VGND VPWR VPWR _09920_/D sky130_fd_sc_hd__a22o_1
X_09090_ _09090_/A _09363_/B VGND VGND VPWR VPWR _09091_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08110_ _07232_/Y _08082_/X _07247_/Y _08083_/X VGND VGND VPWR VPWR _08110_/X sky130_fd_sc_hd__o22a_1
X_05322_ _09920_/Q VGND VGND VPWR VPWR _05322_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05253_ _05253_/A VGND VGND VPWR VPWR _05918_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08041_ _05200_/Y _08207_/A _05302_/Y _08208_/A VGND VGND VPWR VPWR _08041_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05184_ _10141_/Q VGND VGND VPWR VPWR _05184_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09992_ _10006_/CLK _09992_/D repeater407/X VGND VGND VPWR VPWR _09992_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08943_ _08943_/A VGND VGND VPWR VPWR _08961_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08874_ _09253_/A _08782_/Y _08873_/X VGND VGND VPWR VPWR _08874_/Y sky130_fd_sc_hd__a21oi_1
X_07825_ _07825_/A VGND VGND VPWR VPWR _07825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07756_ _06900_/Y _07755_/X _06883_/Y _07642_/X VGND VGND VPWR VPWR _07756_/X sky130_fd_sc_hd__o22a_4
X_04968_ _04968_/A VGND VGND VPWR VPWR _04968_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06707_ _10377_/Q VGND VGND VPWR VPWR _06708_/A sky130_fd_sc_hd__inv_2
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09426_ _09426_/A _09426_/B _09426_/C _09426_/D VGND VGND VPWR VPWR _09451_/A sky130_fd_sc_hd__or4_2
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04899_ _05149_/A VGND VGND VPWR VPWR _05157_/A sky130_fd_sc_hd__clkbuf_2
X_07687_ _10109_/Q VGND VGND VPWR VPWR _07687_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06638_ _09796_/Q _06636_/X _09578_/X _06637_/Y VGND VGND VPWR VPWR _09796_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09357_ _09357_/A _09357_/B _09357_/C _09357_/D VGND VGND VPWR VPWR _09428_/C sky130_fd_sc_hd__or4_4
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06569_ _06569_/A VGND VGND VPWR VPWR _06569_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08308_ _07048_/Y _08211_/A _07957_/A _08212_/A _08307_/X VGND VGND VPWR VPWR _08309_/D
+ sky130_fd_sc_hd__o221a_1
X_09288_ _09288_/A _09354_/D _09442_/D _09288_/D VGND VGND VPWR VPWR _09292_/A sky130_fd_sc_hd__or4_1
XFILLER_60_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08239_ _05291_/Y _08173_/X _05244_/Y _08174_/X VGND VGND VPWR VPWR _08239_/X sky130_fd_sc_hd__o22a_1
XFILLER_153_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10201_ _10513_/CLK _10201_/D _07492_/B VGND VGND VPWR VPWR _10201_/Q sky130_fd_sc_hd__dfrtp_1
X_10132_ _10238_/CLK _10132_/D repeater403/X VGND VGND VPWR VPWR _10132_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10063_ _10224_/CLK _10063_/D repeater405/X VGND VGND VPWR VPWR _10063_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ _06011_/A _06705_/A VGND VGND VPWR VPWR _05942_/A sky130_fd_sc_hd__or2_2
X_05871_ _10181_/Q _05866_/X _06684_/B1 _05867_/Y VGND VGND VPWR VPWR _10181_/D sky130_fd_sc_hd__a22o_1
X_07610_ _07610_/A VGND VGND VPWR VPWR _07827_/A sky130_fd_sc_hd__clkbuf_2
X_08590_ _09379_/A _08590_/B VGND VGND VPWR VPWR _08591_/B sky130_fd_sc_hd__or2_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04822_ _04827_/B VGND VGND VPWR VPWR _04822_/Y sky130_fd_sc_hd__clkinv_2
X_07541_ _07611_/A _07612_/B _07562_/B VGND VGND VPWR VPWR _07805_/A sky130_fd_sc_hd__or3_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07472_ _09776_/Q _09554_/X _09776_/Q _07477_/C _09777_/Q VGND VGND VPWR VPWR _09776_/D
+ sky130_fd_sc_hd__a221o_1
X_09211_ _08461_/X _08578_/B _08934_/A _09206_/B _08577_/X VGND VGND VPWR VPWR _09212_/C
+ sky130_fd_sc_hd__o221a_1
X_06423_ _06390_/X _09621_/X _09650_/X _09885_/Q VGND VGND VPWR VPWR _09885_/D sky130_fd_sc_hd__o22a_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06354_ _09932_/Q _06352_/X _09578_/X _06353_/Y VGND VGND VPWR VPWR _09932_/D sky130_fd_sc_hd__a22o_1
X_09142_ _09142_/A _09348_/C VGND VGND VPWR VPWR _09143_/B sky130_fd_sc_hd__nor2_1
X_05305_ _05305_/A _05305_/B VGND VGND VPWR VPWR _05793_/A sky130_fd_sc_hd__or2_2
XFILLER_190_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06285_ _09971_/Q _06281_/X _09576_/X _06282_/Y VGND VGND VPWR VPWR _09971_/D sky130_fd_sc_hd__a22o_1
X_09073_ _09073_/A _09073_/B VGND VGND VPWR VPWR _09290_/C sky130_fd_sc_hd__or2_1
XFILLER_162_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05236_ _05236_/A _05236_/B _05236_/C _05236_/D VGND VGND VPWR VPWR _05365_/A sky130_fd_sc_hd__and4_1
X_08024_ _05324_/Y _08183_/A _08017_/X _08023_/X VGND VGND VPWR VPWR _08050_/C sky130_fd_sc_hd__o211a_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05167_ _05167_/A _05359_/A VGND VGND VPWR VPWR _05689_/B sky130_fd_sc_hd__or2_2
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09975_ _10000_/CLK _09975_/D repeater405/X VGND VGND VPWR VPWR _09975_/Q sky130_fd_sc_hd__dfstp_1
X_05098_ _05160_/A _05351_/A VGND VGND VPWR VPWR _05625_/C sky130_fd_sc_hd__or2_2
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08926_ _08926_/A _09388_/B _09370_/B _09285_/B VGND VGND VPWR VPWR _08932_/A sky130_fd_sc_hd__or4_1
X_08857_ _09420_/B _08857_/B VGND VGND VPWR VPWR _08859_/A sky130_fd_sc_hd__or2_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07808_ _06829_/Y _07806_/X _06815_/Y _07807_/X VGND VGND VPWR VPWR _07808_/X sky130_fd_sc_hd__o22a_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08788_ _08788_/A _08788_/B VGND VGND VPWR VPWR _09400_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07739_ _06950_/Y _06232_/X _06997_/Y _07533_/A _07738_/X VGND VGND VPWR VPWR _07743_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09409_ _09409_/A VGND VGND VPWR VPWR _09409_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10115_ _10119_/CLK _10115_/D repeater403/X VGND VGND VPWR VPWR _10115_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10046_ _10127_/CLK _10046_/D repeater409/X VGND VGND VPWR VPWR _10046_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _07503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06070_ _10062_/Q _06067_/X _09581_/X _06069_/X VGND VGND VPWR VPWR _10062_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05021_ _05021_/A VGND VGND VPWR VPWR _05021_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06972_ _06967_/Y _05882_/A _06968_/Y _05896_/B _06971_/X VGND VGND VPWR VPWR _06985_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09760_ _09919_/CLK _09760_/D VGND VGND VPWR VPWR _09760_/Q sky130_fd_sc_hd__dfxtp_2
X_09691_ _08372_/X input194/X _09698_/S VGND VGND VPWR VPWR _09691_/X sky130_fd_sc_hd__mux2_1
X_05923_ _10151_/Q _05919_/X _06683_/B1 _05920_/Y VGND VGND VPWR VPWR _10151_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08711_ _08684_/A _08678_/X _08708_/X _09115_/A _09162_/B VGND VGND VPWR VPWR _08711_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08642_ _08379_/B _08794_/B _08379_/B _08794_/B VGND VGND VPWR VPWR _08643_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05854_ _05854_/A VGND VGND VPWR VPWR _05855_/A sky130_fd_sc_hd__inv_2
X_04805_ _10284_/Q input78/X input79/X VGND VGND VPWR VPWR _09732_/A sky130_fd_sc_hd__mux2_2
X_05785_ _05874_/A _05785_/B VGND VGND VPWR VPWR _05787_/A sky130_fd_sc_hd__or2_1
X_08573_ _08529_/A _08552_/B _08563_/X _08570_/X _08572_/X VGND VGND VPWR VPWR _08573_/X
+ sky130_fd_sc_hd__o2111a_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ _07524_/A _07597_/C VGND VGND VPWR VPWR _07601_/B sky130_fd_sc_hd__or2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07455_ _06835_/X _07451_/X _09740_/Q _07453_/X VGND VGND VPWR VPWR _09740_/D sky130_fd_sc_hd__o22a_1
X_06406_ _09901_/Q _06403_/X _09581_/X _06405_/X VGND VGND VPWR VPWR _09901_/D sky130_fd_sc_hd__a22o_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07386_ _07381_/Y _06401_/A _07382_/Y _05541_/B _07385_/X VGND VGND VPWR VPWR _07393_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06337_ _06337_/A VGND VGND VPWR VPWR _06481_/A sky130_fd_sc_hd__clkbuf_2
X_09125_ _09379_/B _09289_/A VGND VGND VPWR VPWR _09398_/A sky130_fd_sc_hd__or2_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09056_ _09295_/A _09295_/B _09056_/C VGND VGND VPWR VPWR _09352_/C sky130_fd_sc_hd__or3_2
X_06268_ _06269_/A VGND VGND VPWR VPWR _06268_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05219_ _05338_/B VGND VGND VPWR VPWR _05349_/B sky130_fd_sc_hd__clkbuf_2
X_08007_ _08045_/C VGND VGND VPWR VPWR _08037_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06199_ _08044_/A VGND VGND VPWR VPWR _08019_/B sky130_fd_sc_hd__clkbuf_2
X_09958_ _10288_/CLK _09958_/D repeater406/X VGND VGND VPWR VPWR _09958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08909_ _09015_/B VGND VGND VPWR VPWR _08909_/Y sky130_fd_sc_hd__inv_2
X_09889_ _10397_/CLK _09889_/D repeater409/X VGND VGND VPWR VPWR _09889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 wb_dat_i[15] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__clkbuf_1
Xinput160 wb_adr_i[6] VGND VGND VPWR VPWR _08571_/C sky130_fd_sc_hd__buf_4
XFILLER_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput182 wb_dat_i[25] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__clkbuf_1
Xinput193 wb_dat_i[6] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__clkbuf_1
X_10029_ _10135_/CLK _10029_/D _07492_/B VGND VGND VPWR VPWR _10029_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05570_ _10355_/Q _05568_/X _09547_/A1 _05569_/Y VGND VGND VPWR VPWR _10355_/D sky130_fd_sc_hd__a22o_1
XFILLER_176_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07240_ _10177_/Q VGND VGND VPWR VPWR _07240_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07171_ input45/X _06697_/A _10461_/Q _06689_/A _07170_/X VGND VGND VPWR VPWR _07181_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06122_ _06304_/A _06122_/B VGND VGND VPWR VPWR _06124_/A sky130_fd_sc_hd__or2_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06053_ _06053_/A VGND VGND VPWR VPWR _06893_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_125_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05004_ _10443_/Q _04995_/A _09536_/A3 _04996_/A VGND VGND VPWR VPWR _10443_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09812_ _09572_/A1 _09812_/D _06574_/X VGND VGND VPWR VPWR _09812_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06955_ _09819_/Q VGND VGND VPWR VPWR _06955_/Y sky130_fd_sc_hd__clkinv_4
X_09743_ _09752_/CLK _09743_/D VGND VGND VPWR VPWR _09743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05906_ _10160_/Q _05898_/A hold46/X _05899_/A VGND VGND VPWR VPWR _10160_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09674_ _09673_/X _10391_/Q _10299_/Q VGND VGND VPWR VPWR _09674_/X sky130_fd_sc_hd__mux2_4
X_06886_ _10190_/Q VGND VGND VPWR VPWR _06886_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _08806_/A VGND VGND VPWR VPWR _08837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05837_ _10201_/Q _05831_/X _09536_/A3 _05832_/Y VGND VGND VPWR VPWR _10201_/D sky130_fd_sc_hd__a22o_1
X_08556_ _09233_/A _08556_/B _08571_/C _08556_/D VGND VGND VPWR VPWR _08921_/B sky130_fd_sc_hd__or4_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05768_ _10242_/Q _05763_/X _09579_/X _05765_/X VGND VGND VPWR VPWR _10242_/D sky130_fd_sc_hd__a22o_1
X_07507_ _07602_/D VGND VGND VPWR VPWR _07608_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08487_ _08921_/C VGND VGND VPWR VPWR _08582_/A sky130_fd_sc_hd__buf_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05699_ _09679_/X _05715_/B VGND VGND VPWR VPWR _05702_/A sky130_fd_sc_hd__or2_2
X_07438_ _07450_/A _07438_/B VGND VGND VPWR VPWR _07440_/A sky130_fd_sc_hd__or2_4
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07369_ _10013_/Q VGND VGND VPWR VPWR _07369_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09108_ _08736_/A _09048_/A _09101_/Y _09098_/A _09107_/X VGND VGND VPWR VPWR _09108_/X
+ sky130_fd_sc_hd__o221a_1
X_10380_ _10382_/CLK _10380_/D _05515_/X VGND VGND VPWR VPWR _10380_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09039_ _08457_/X _09218_/A _09372_/A _08457_/X VGND VGND VPWR VPWR _09039_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06740_ _06740_/A _06740_/B _06740_/C _06740_/D VGND VGND VPWR VPWR _06740_/X sky130_fd_sc_hd__and4_1
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06671_ _06677_/A VGND VGND VPWR VPWR _06672_/A sky130_fd_sc_hd__clkbuf_1
X_08410_ _08485_/A _08492_/B _06464_/X VGND VGND VPWR VPWR _08913_/B sky130_fd_sc_hd__o21ai_2
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05622_ _10324_/Q _05616_/X _09536_/A3 _05617_/Y VGND VGND VPWR VPWR _10324_/D sky130_fd_sc_hd__a22o_1
X_09390_ _09390_/A _09390_/B _09390_/C VGND VGND VPWR VPWR _09435_/C sky130_fd_sc_hd__or3_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05553_ _05553_/A VGND VGND VPWR VPWR _05553_/X sky130_fd_sc_hd__clkbuf_2
X_08341_ _09804_/Q _08341_/B VGND VGND VPWR VPWR _08343_/A sky130_fd_sc_hd__nand2_1
X_05484_ _09788_/Q VGND VGND VPWR VPWR _09532_/A sky130_fd_sc_hd__inv_2
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08272_ _07328_/Y _08211_/X _07907_/A _08212_/X _08271_/X VGND VGND VPWR VPWR _08273_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07223_ _07221_/Y _05433_/A _07222_/Y _06551_/B VGND VGND VPWR VPWR _07223_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07154_ _07152_/Y _05541_/B _07153_/Y _04871_/B VGND VGND VPWR VPWR _07154_/X sky130_fd_sc_hd__o22a_1
X_07085_ _10178_/Q VGND VGND VPWR VPWR _07085_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06105_ _10039_/Q _06098_/A _09660_/A1 _06099_/A VGND VGND VPWR VPWR _10039_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06036_ _06036_/A VGND VGND VPWR VPWR _06037_/B sky130_fd_sc_hd__buf_2
XFILLER_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07987_ _07987_/A _07987_/B _07987_/C _07987_/D VGND VGND VPWR VPWR _07988_/C sky130_fd_sc_hd__and4_1
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09726_ _10292_/Q _09505_/A VGND VGND VPWR VPWR _09726_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06938_ _10231_/Q VGND VGND VPWR VPWR _06938_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06869_ _10094_/Q VGND VGND VPWR VPWR _06869_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _08329_/Y _05713_/A _09772_/Q VGND VGND VPWR VPWR _09780_/D sky130_fd_sc_hd__mux2_1
X_09588_ _10315_/Q _09581_/X _09699_/S VGND VGND VPWR VPWR _09588_/X sky130_fd_sc_hd__mux2_1
X_08608_ _09299_/A _08608_/B VGND VGND VPWR VPWR _08609_/C sky130_fd_sc_hd__or2_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08539_ _08929_/A _08921_/C VGND VGND VPWR VPWR _08935_/B sky130_fd_sc_hd__or2_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10501_ _10504_/CLK _10501_/D repeater404/X VGND VGND VPWR VPWR _10501_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10432_ _10483_/CLK _10432_/D _05034_/A VGND VGND VPWR VPWR _10432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10363_ _10364_/CLK _10363_/D repeater410/X VGND VGND VPWR VPWR _10363_/Q sky130_fd_sc_hd__dfrtp_1
X_10294_ _10296_/CLK _10294_/D repeater402/X VGND VGND VPWR VPWR _10294_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08890_ _08890_/A _08890_/B VGND VGND VPWR VPWR _08890_/Y sky130_fd_sc_hd__nor2_1
X_07910_ _07383_/Y _07825_/X _07300_/Y _07827_/X _07909_/X VGND VGND VPWR VPWR _07911_/D
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_12_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10354_/CLK sky130_fd_sc_hd__clkbuf_16
X_07841_ _06751_/Y _07792_/X _06711_/Y _07793_/X _07840_/X VGND VGND VPWR VPWR _07848_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07772_ _10060_/Q VGND VGND VPWR VPWR _07772_/Y sky130_fd_sc_hd__inv_2
X_09511_ _09511_/A VGND VGND VPWR VPWR _09512_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04984_ _10457_/Q _04980_/X _09580_/X _04982_/X VGND VGND VPWR VPWR _10457_/D sky130_fd_sc_hd__a22o_1
X_06723_ _10364_/Q VGND VGND VPWR VPWR _06723_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10268_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06654_ _06654_/A VGND VGND VPWR VPWR _06654_/X sky130_fd_sc_hd__clkbuf_1
X_09442_ _09442_/A _09442_/B _09442_/C _09442_/D VGND VGND VPWR VPWR _09443_/B sky130_fd_sc_hd__or4_2
XFILLER_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09373_ _09372_/C _08461_/X _09372_/B _09372_/X _09267_/Y VGND VGND VPWR VPWR _09373_/X
+ sky130_fd_sc_hd__o311a_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06585_ _06585_/A _07483_/C VGND VGND VPWR VPWR _06585_/X sky130_fd_sc_hd__or2_1
X_05605_ _05605_/A VGND VGND VPWR VPWR _05606_/A sky130_fd_sc_hd__inv_2
X_08324_ _07018_/Y _08205_/A _06949_/Y _08206_/A _08323_/X VGND VGND VPWR VPWR _08327_/C
+ sky130_fd_sc_hd__o221a_1
X_05536_ _10373_/Q _05529_/X _09658_/A1 _05531_/X VGND VGND VPWR VPWR _10373_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05467_ _05497_/A VGND VGND VPWR VPWR _05468_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08255_ _08255_/A _08255_/B _08255_/C _08255_/D VGND VGND VPWR VPWR _08256_/D sky130_fd_sc_hd__and4_2
X_05398_ _05398_/A VGND VGND VPWR VPWR _05398_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07206_ _10130_/Q VGND VGND VPWR VPWR _07206_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08186_ _08186_/A VGND VGND VPWR VPWR _08186_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07137_ _09507_/A _05727_/A _09487_/A _06095_/A _07136_/X VGND VGND VPWR VPWR _07156_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_165_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput261 _09723_/Z VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_2
X_07068_ _10248_/Q VGND VGND VPWR VPWR _09503_/A sky130_fd_sc_hd__inv_6
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput250 _09713_/Z VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_1
Xoutput272 _09733_/Z VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_2
X_06019_ _10092_/Q _06012_/X _09550_/A0 _06014_/X VGND VGND VPWR VPWR _10092_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput294 _10441_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_2
Xoutput283 _09572_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09709_ _09709_/A _09471_/A VGND VGND VPWR VPWR _09709_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_74_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10415_ _04807_/A1 _10415_/D _05407_/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfrtp_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10346_ _10349_/CLK _10346_/D repeater404/X VGND VGND VPWR VPWR _10346_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10277_ _10405_/CLK _10277_/D hold41/X VGND VGND VPWR VPWR _10277_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06370_ _09921_/Q _06362_/A _09661_/A1 _06363_/A VGND VGND VPWR VPWR _09921_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05321_ _05321_/A _05321_/B _05321_/C _05321_/D VGND VGND VPWR VPWR _05365_/C sky130_fd_sc_hd__and4_1
XFILLER_174_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05252_ _05286_/B _06630_/B VGND VGND VPWR VPWR _05253_/A sky130_fd_sc_hd__or2_2
X_08040_ _08040_/A _08046_/C _08040_/C VGND VGND VPWR VPWR _08208_/A sky130_fd_sc_hd__or3_4
XFILLER_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05183_ _05183_/A _05183_/B _05183_/C _05182_/X VGND VGND VPWR VPWR _05366_/C sky130_fd_sc_hd__or4b_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09991_ _10006_/CLK _09991_/D repeater407/X VGND VGND VPWR VPWR _09991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08942_ _08951_/A _08942_/B VGND VGND VPWR VPWR _09198_/B sky130_fd_sc_hd__nor2_1
X_08873_ _09085_/B _09139_/A _08872_/X VGND VGND VPWR VPWR _08873_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07824_ _06811_/Y _07768_/X _06808_/Y _07769_/X _07823_/X VGND VGND VPWR VPWR _07832_/C
+ sky130_fd_sc_hd__o221a_1
X_07755_ _07755_/A VGND VGND VPWR VPWR _07755_/X sky130_fd_sc_hd__buf_2
X_04967_ _04967_/A VGND VGND VPWR VPWR _04968_/A sky130_fd_sc_hd__inv_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07686_ _07263_/Y _07533_/D _07232_/Y _07651_/X _07685_/X VGND VGND VPWR VPWR _07694_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06706_ input28/X _06704_/X _10140_/Q _06705_/Y VGND VGND VPWR VPWR _06715_/B sky130_fd_sc_hd__a22o_1
X_06637_ _06637_/A VGND VGND VPWR VPWR _06637_/Y sky130_fd_sc_hd__inv_2
X_09425_ _09425_/A _09425_/B _09425_/C _09425_/D VGND VGND VPWR VPWR _09426_/B sky130_fd_sc_hd__or4_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04898_ _05806_/A VGND VGND VPWR VPWR _06538_/A sky130_fd_sc_hd__buf_4
X_09356_ _09389_/D _09431_/C _09443_/A _09387_/D VGND VGND VPWR VPWR _09359_/A sky130_fd_sc_hd__or4_4
X_06568_ _06568_/A VGND VGND VPWR VPWR _06569_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05519_ _05519_/A VGND VGND VPWR VPWR _05519_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06499_ _09851_/Q _06495_/X _09576_/X _06496_/Y VGND VGND VPWR VPWR _09851_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08307_ _07093_/Y _08213_/A _07119_/Y _08214_/A VGND VGND VPWR VPWR _08307_/X sky130_fd_sc_hd__o22a_1
X_09287_ _09287_/A _09287_/B _09287_/C VGND VGND VPWR VPWR _09288_/D sky130_fd_sc_hd__or3_1
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08238_ _08238_/A _08238_/B _08238_/C _08238_/D VGND VGND VPWR VPWR _08238_/Y sky130_fd_sc_hd__nand4_4
XFILLER_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10200_ _10244_/CLK _10200_/D repeater402/X VGND VGND VPWR VPWR _10200_/Q sky130_fd_sc_hd__dfrtp_1
X_08169_ _06859_/Y _08094_/X _06883_/Y _08095_/X VGND VGND VPWR VPWR _08169_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10131_ _10238_/CLK hold49/X repeater403/X VGND VGND VPWR VPWR _10131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10062_ _10062_/CLK _10062_/D repeater405/X VGND VGND VPWR VPWR _10062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10336_/CLK _10329_/D repeater409/X VGND VGND VPWR VPWR _10329_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_112_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05870_ _10182_/Q _05866_/X _06683_/B1 _05867_/Y VGND VGND VPWR VPWR _10182_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04821_ _05318_/A _05155_/A VGND VGND VPWR VPWR _04827_/B sky130_fd_sc_hd__or2_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07540_ _07819_/A VGND VGND VPWR VPWR _07659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07471_ _06133_/Y _06262_/B _07470_/Y _09775_/Q VGND VGND VPWR VPWR _09775_/D sky130_fd_sc_hd__a2bb2o_1
X_09210_ _08925_/A _09206_/B _08543_/X _08928_/A VGND VGND VPWR VPWR _09212_/B sky130_fd_sc_hd__o211a_1
X_06422_ _06417_/X _09623_/X _09650_/X _09886_/Q VGND VGND VPWR VPWR _09886_/D sky130_fd_sc_hd__o22a_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06353_ _06353_/A VGND VGND VPWR VPWR _06353_/Y sky130_fd_sc_hd__inv_2
X_09141_ _09222_/A _09141_/B VGND VGND VPWR VPWR _09348_/C sky130_fd_sc_hd__or2_1
XFILLER_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09072_ _09397_/B _09201_/B VGND VGND VPWR VPWR _09387_/A sky130_fd_sc_hd__or2_1
X_05304_ _10219_/Q VGND VGND VPWR VPWR _05304_/Y sky130_fd_sc_hd__clkinv_2
X_06284_ _09972_/Q _06281_/X _09550_/A0 _06282_/Y VGND VGND VPWR VPWR _09972_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08023_ _05212_/Y _08186_/A _05273_/Y _08187_/A _08022_/X VGND VGND VPWR VPWR _08023_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05235_ _05225_/Y _06438_/A _05227_/Y _06351_/B _05234_/X VGND VGND VPWR VPWR _05236_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05166_ _09677_/S VGND VGND VPWR VPWR _06697_/A sky130_fd_sc_hd__clkinv_2
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09974_ _10000_/CLK _09974_/D repeater405/X VGND VGND VPWR VPWR _09974_/Q sky130_fd_sc_hd__dfstp_1
X_05097_ _05155_/B VGND VGND VPWR VPWR _05351_/A sky130_fd_sc_hd__clkbuf_4
X_08925_ _08925_/A _08933_/A VGND VGND VPWR VPWR _09285_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08856_ _08856_/A _09076_/A VGND VGND VPWR VPWR _08857_/B sky130_fd_sc_hd__or2_1
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07807_ _07807_/A VGND VGND VPWR VPWR _07807_/X sky130_fd_sc_hd__buf_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05999_ _10103_/Q _05994_/X hold46/X _05995_/Y VGND VGND VPWR VPWR _10103_/D sky130_fd_sc_hd__a22o_1
X_08787_ _08864_/A _08787_/B VGND VGND VPWR VPWR _08788_/B sky130_fd_sc_hd__or2_1
X_07738_ _07738_/A _07770_/B VGND VGND VPWR VPWR _07738_/X sky130_fd_sc_hd__or2_1
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07669_ _07346_/Y _07667_/X _07356_/Y _07668_/X VGND VGND VPWR VPWR _07669_/X sky130_fd_sc_hd__o22a_1
X_09408_ _09408_/A _09408_/B _09408_/C _09439_/D VGND VGND VPWR VPWR _09409_/A sky130_fd_sc_hd__or4_1
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09339_ _09339_/A _09339_/B _09339_/C _09339_/D VGND VGND VPWR VPWR _09398_/D sky130_fd_sc_hd__or4_2
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10114_ _10371_/CLK _10114_/D repeater405/X VGND VGND VPWR VPWR _10114_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10045_ _10127_/CLK _10045_/D repeater409/X VGND VGND VPWR VPWR _10045_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 _07504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05020_ _05021_/A VGND VGND VPWR VPWR _05020_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06971_ _06969_/Y _05293_/A _06970_/Y _06515_/A VGND VGND VPWR VPWR _06971_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09690_ _08370_/X input193/X _09698_/S VGND VGND VPWR VPWR _09690_/X sky130_fd_sc_hd__mux2_1
X_05922_ _10152_/Q _05919_/X _09577_/X _05920_/Y VGND VGND VPWR VPWR _10152_/D sky130_fd_sc_hd__a22o_1
X_08710_ _08710_/A _08831_/B VGND VGND VPWR VPWR _09162_/B sky130_fd_sc_hd__or2_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _08641_/A _08641_/B _08641_/C VGND VGND VPWR VPWR _08794_/B sky130_fd_sc_hd__or3_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05853_ _05854_/A VGND VGND VPWR VPWR _05853_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_04804_ _10283_/Q input80/X input79/X VGND VGND VPWR VPWR _09731_/A sky130_fd_sc_hd__mux2_2
X_08572_ _08582_/A _08685_/B _09012_/A _08563_/A _09011_/A VGND VGND VPWR VPWR _08572_/X
+ sky130_fd_sc_hd__o32a_1
X_05784_ _06327_/A VGND VGND VPWR VPWR _05874_/A sky130_fd_sc_hd__buf_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07523_ _07523_/A VGND VGND VPWR VPWR _07533_/B sky130_fd_sc_hd__clkbuf_2
X_07454_ _06759_/X _07451_/X _09741_/Q _07453_/X VGND VGND VPWR VPWR _09741_/D sky130_fd_sc_hd__o22a_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06405_ _06405_/A VGND VGND VPWR VPWR _06405_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07385_ _07383_/Y _06079_/B _07384_/Y _06312_/A VGND VGND VPWR VPWR _07385_/X sky130_fd_sc_hd__o22a_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06336_ _09941_/Q _06330_/X _09536_/A3 _06331_/Y VGND VGND VPWR VPWR _09941_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09124_ _09124_/A VGND VGND VPWR VPWR _09379_/B sky130_fd_sc_hd__inv_2
XFILLER_163_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09055_ _09277_/A _09055_/B VGND VGND VPWR VPWR _09058_/B sky130_fd_sc_hd__or2_2
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06267_ _06313_/A _06267_/B VGND VGND VPWR VPWR _06269_/A sky130_fd_sc_hd__or2_2
X_05218_ _09983_/Q VGND VGND VPWR VPWR _05218_/Y sky130_fd_sc_hd__clkinv_4
X_08006_ _08006_/A _10004_/Q VGND VGND VPWR VPWR _08045_/C sky130_fd_sc_hd__or2_1
XFILLER_190_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06198_ _08046_/A _07994_/B VGND VGND VPWR VPWR _08044_/A sky130_fd_sc_hd__or2_2
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05149_ _05149_/A _05329_/A VGND VGND VPWR VPWR _05603_/B sky130_fd_sc_hd__or2_1
X_09957_ _10288_/CLK _09957_/D repeater406/X VGND VGND VPWR VPWR _09957_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08908_ _08908_/A _08908_/B VGND VGND VPWR VPWR _09015_/B sky130_fd_sc_hd__or2_2
XFILLER_106_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09888_ _10397_/CLK _09888_/D repeater409/X VGND VGND VPWR VPWR _09888_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08839_ _08665_/Y _09096_/B _08838_/X VGND VGND VPWR VPWR _08839_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput172 wb_dat_i[16] VGND VGND VPWR VPWR _08357_/B sky130_fd_sc_hd__clkbuf_1
Xinput150 wb_adr_i[26] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_adr_i[7] VGND VGND VPWR VPWR _09236_/A sky130_fd_sc_hd__buf_4
X_10028_ _10411_/CLK _10028_/D repeater407/X VGND VGND VPWR VPWR _10028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput183 wb_dat_i[26] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[7] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07170_ input54/X _05114_/A _09768_/Q _05146_/Y VGND VGND VPWR VPWR _07170_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06121_ _06121_/A VGND VGND VPWR VPWR _06122_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_145_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06052_ _10071_/Q _06046_/X _09536_/A3 _06047_/Y VGND VGND VPWR VPWR _10071_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05003_ _10444_/Q _04995_/A _06684_/B1 _04996_/A VGND VGND VPWR VPWR _10444_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09811_ _09572_/A1 _09811_/D _06578_/X VGND VGND VPWR VPWR _09811_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09742_ _09752_/CLK _09742_/D VGND VGND VPWR VPWR _09742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06954_ _10361_/Q VGND VGND VPWR VPWR _06954_/Y sky130_fd_sc_hd__clkinv_4
X_05905_ _10161_/Q _05898_/A _09660_/A1 _05899_/A VGND VGND VPWR VPWR _10161_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06885_ _09838_/Q VGND VGND VPWR VPWR _06885_/Y sky130_fd_sc_hd__clkinv_2
X_09673_ _09799_/Q input58/X _09773_/Q VGND VGND VPWR VPWR _09673_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08624_ _08624_/A _09344_/A VGND VGND VPWR VPWR _08806_/A sky130_fd_sc_hd__or2_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05836_ _10202_/Q _05831_/X _06684_/B1 _05832_/Y VGND VGND VPWR VPWR _10202_/D sky130_fd_sc_hd__a22o_1
X_05767_ _10243_/Q _05763_/X _09580_/X _05765_/X VGND VGND VPWR VPWR _10243_/D sky130_fd_sc_hd__a22o_1
X_08555_ _08582_/A _08575_/A VGND VGND VPWR VPWR _08563_/A sky130_fd_sc_hd__or2_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07506_ _10329_/Q VGND VGND VPWR VPWR _07506_/Y sky130_fd_sc_hd__inv_2
X_05698_ _10283_/Q _05691_/A _09574_/X _05692_/A VGND VGND VPWR VPWR _10283_/D sky130_fd_sc_hd__a22o_1
X_08486_ _08905_/B VGND VGND VPWR VPWR _08921_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07437_ _09783_/Q VGND VGND VPWR VPWR _07438_/B sky130_fd_sc_hd__inv_2
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ _09863_/Q VGND VGND VPWR VPWR _07368_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09107_ _08849_/A _08810_/B _09103_/X _09106_/Y VGND VGND VPWR VPWR _09107_/X sky130_fd_sc_hd__o211a_1
X_06319_ _09952_/Q _06314_/X _09579_/X _06316_/X VGND VGND VPWR VPWR _09952_/D sky130_fd_sc_hd__a22o_1
X_07299_ _10056_/Q VGND VGND VPWR VPWR _07299_/Y sky130_fd_sc_hd__inv_2
X_09038_ _09432_/A _09425_/A _09038_/C VGND VGND VPWR VPWR _09040_/A sky130_fd_sc_hd__or3_1
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 input92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06670_ _06670_/A VGND VGND VPWR VPWR _06670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05621_ _10325_/Q _05616_/X _06684_/B1 _05617_/Y VGND VGND VPWR VPWR _10325_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05552_ _05552_/A VGND VGND VPWR VPWR _05553_/A sky130_fd_sc_hd__inv_2
X_08340_ _08340_/A VGND VGND VPWR VPWR _08341_/B sky130_fd_sc_hd__inv_2
X_05483_ _05483_/A VGND VGND VPWR VPWR _05483_/X sky130_fd_sc_hd__clkbuf_1
X_08271_ _07409_/Y _08213_/X _07365_/Y _08214_/X VGND VGND VPWR VPWR _08271_/X sky130_fd_sc_hd__o22a_1
XFILLER_177_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07222_ _09817_/Q VGND VGND VPWR VPWR _07222_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07153_ _10499_/Q VGND VGND VPWR VPWR _07153_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06104_ _10040_/Q _06097_/X _09658_/A1 _06099_/X VGND VGND VPWR VPWR _10040_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07084_ _09950_/Q VGND VGND VPWR VPWR _09477_/A sky130_fd_sc_hd__inv_6
XFILLER_172_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06035_ _10081_/Q _06026_/A _09536_/A3 _06027_/A VGND VGND VPWR VPWR _10081_/D sky130_fd_sc_hd__a22o_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07986_ _06986_/Y _07825_/A _06909_/Y _07827_/A _07985_/X VGND VGND VPWR VPWR _07987_/D
+ sky130_fd_sc_hd__o221a_1
X_09725_ _10291_/Q _09503_/A VGND VGND VPWR VPWR _09725_/Z sky130_fd_sc_hd__ebufn_1
X_06937_ _10093_/Q VGND VGND VPWR VPWR _06937_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09656_ _10428_/Q _06759_/X _09680_/S VGND VGND VPWR VPWR _09656_/X sky130_fd_sc_hd__mux2_1
X_08607_ _08457_/X _08461_/X _08606_/X VGND VGND VPWR VPWR _08608_/B sky130_fd_sc_hd__o21ai_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06868_ _09952_/Q VGND VGND VPWR VPWR _06868_/Y sky130_fd_sc_hd__inv_2
X_09587_ _10314_/Q _09580_/X _09699_/S VGND VGND VPWR VPWR _09587_/X sky130_fd_sc_hd__mux2_1
X_05819_ _10211_/Q _05810_/A _09659_/A1 _05811_/A VGND VGND VPWR VPWR _10211_/D sky130_fd_sc_hd__a22o_1
X_06799_ _09939_/Q VGND VGND VPWR VPWR _06799_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08538_ _08929_/A VGND VGND VPWR VPWR _08934_/A sky130_fd_sc_hd__buf_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _08695_/A VGND VGND VPWR VPWR _09295_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10500_ _10500_/CLK _10500_/D repeater407/X VGND VGND VPWR VPWR _10500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10431_ _10471_/CLK _10431_/D repeater409/X VGND VGND VPWR VPWR _10431_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10362_ _10364_/CLK _10362_/D repeater410/X VGND VGND VPWR VPWR _10362_/Q sky130_fd_sc_hd__dfrtp_1
X_10293_ _10296_/CLK _10293_/D repeater402/X VGND VGND VPWR VPWR _10293_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_8_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10254_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07840_ _06752_/Y _07794_/X _06753_/Y _07795_/X VGND VGND VPWR VPWR _07840_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07771_ _06886_/Y _07768_/X _06858_/Y _07769_/X _07770_/X VGND VGND VPWR VPWR _07775_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09510_ _09510_/A VGND VGND VPWR VPWR _09510_/X sky130_fd_sc_hd__clkbuf_1
X_06722_ _09901_/Q VGND VGND VPWR VPWR _06722_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_04983_ _10458_/Q _04980_/X _09581_/X _04982_/X VGND VGND VPWR VPWR _10458_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06653_ _06655_/A VGND VGND VPWR VPWR _06654_/A sky130_fd_sc_hd__clkbuf_1
X_09441_ _09441_/A VGND VGND VPWR VPWR _09441_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09372_ _09372_/A _09372_/B _09372_/C VGND VGND VPWR VPWR _09372_/X sky130_fd_sc_hd__or3_1
X_06584_ _06584_/A VGND VGND VPWR VPWR _06584_/X sky130_fd_sc_hd__clkbuf_1
X_05604_ _05605_/A VGND VGND VPWR VPWR _05604_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08323_ _06993_/Y _08207_/A _06928_/Y _08208_/A VGND VGND VPWR VPWR _08323_/X sky130_fd_sc_hd__o22a_1
X_05535_ _10374_/Q _05529_/X _09545_/A1 _05531_/X VGND VGND VPWR VPWR _10374_/D sky130_fd_sc_hd__a22o_1
XFILLER_165_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08254_ _05345_/Y _08211_/X _07881_/A _08212_/X _08253_/X VGND VGND VPWR VPWR _08255_/D
+ sky130_fd_sc_hd__o221a_1
X_05466_ _09694_/X _05449_/X _10393_/Q _05451_/X VGND VGND VPWR VPWR _10393_/D sky130_fd_sc_hd__a22o_1
X_05397_ _05397_/A VGND VGND VPWR VPWR _05398_/A sky130_fd_sc_hd__inv_2
X_07205_ _07200_/Y _05761_/A _07201_/Y _05838_/A _07204_/X VGND VGND VPWR VPWR _07218_/B
+ sky130_fd_sc_hd__o221a_1
X_08185_ _06811_/Y _08184_/X _06793_/Y _08158_/X VGND VGND VPWR VPWR _08185_/X sky130_fd_sc_hd__o22a_1
XFILLER_180_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07136_ _07134_/Y _05253_/A _07135_/Y _05575_/A VGND VGND VPWR VPWR _07136_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07067_ _10389_/Q VGND VGND VPWR VPWR _07067_/Y sky130_fd_sc_hd__clkinv_2
Xoutput262 _09724_/Z VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_2
X_06018_ _10093_/Q _06012_/X _09547_/A1 _06014_/X VGND VGND VPWR VPWR _10093_/D sky130_fd_sc_hd__a22o_1
Xoutput251 _09714_/Z VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__buf_2
Xoutput240 _09462_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_2
Xoutput273 _09563_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput295 _10442_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_2
Xoutput284 _07492_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_2
X_07969_ _06998_/Y _07794_/A _06949_/Y _07795_/A VGND VGND VPWR VPWR _07969_/X sky130_fd_sc_hd__o22a_1
X_09708_ _09708_/A _09469_/A VGND VGND VPWR VPWR _09708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09639_ _10425_/Q _07030_/X _09680_/S VGND VGND VPWR VPWR _09639_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10414_ _04807_/A1 _10414_/D _05411_/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfrtp_1
XFILLER_143_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10345_ _10349_/CLK _10345_/D repeater405/X VGND VGND VPWR VPWR _10345_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10276_ _10405_/CLK _10276_/D hold41/X VGND VGND VPWR VPWR _10276_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ _05310_/Y _06053_/A _05312_/Y _05740_/B _05319_/X VGND VGND VPWR VPWR _05321_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05251_ _10149_/Q VGND VGND VPWR VPWR _05251_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05182_ _05172_/Y _06024_/B _05175_/Y _06045_/B _05181_/X VGND VGND VPWR VPWR _05182_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09990_ _10006_/CLK _09990_/D repeater407/X VGND VGND VPWR VPWR _09990_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08941_ _08941_/A _09068_/B _09287_/B VGND VGND VPWR VPWR _08945_/A sky130_fd_sc_hd__or3_1
X_08872_ _09415_/A _08872_/B VGND VGND VPWR VPWR _08872_/X sky130_fd_sc_hd__or2_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07823_ _07823_/A _07932_/B VGND VGND VPWR VPWR _07823_/X sky130_fd_sc_hd__or2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04966_ _04967_/A VGND VGND VPWR VPWR _04966_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07754_ _10034_/Q VGND VGND VPWR VPWR _07754_/Y sky130_fd_sc_hd__inv_2
X_07685_ _07233_/Y _07652_/X _07282_/Y _07653_/X VGND VGND VPWR VPWR _07685_/X sky130_fd_sc_hd__o22a_1
X_06705_ _06705_/A VGND VGND VPWR VPWR _06705_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06636_ _06637_/A VGND VGND VPWR VPWR _06636_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_04897_ _10488_/Q _04888_/A _09659_/A1 _04889_/A VGND VGND VPWR VPWR _10488_/D sky130_fd_sc_hd__a22o_1
X_09424_ _09450_/A _09424_/B VGND VGND VPWR VPWR _09424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09355_ _08665_/Y _09096_/B _09021_/B _09070_/D _09288_/D VGND VGND VPWR VPWR _09387_/D
+ sky130_fd_sc_hd__a2111o_4
X_06567_ _06567_/A VGND VGND VPWR VPWR _09814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05518_ _05518_/A VGND VGND VPWR VPWR _05519_/A sky130_fd_sc_hd__clkbuf_1
X_06498_ _09852_/Q _06495_/X _09577_/X _06496_/Y VGND VGND VPWR VPWR _09852_/D sky130_fd_sc_hd__a22o_1
X_08306_ _07141_/Y _08205_/A _07060_/Y _08206_/A _08305_/X VGND VGND VPWR VPWR _08309_/C
+ sky130_fd_sc_hd__o221a_1
X_09286_ _09286_/A _09286_/B _09286_/C VGND VGND VPWR VPWR _09442_/D sky130_fd_sc_hd__or3_1
XFILLER_193_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05449_ _05450_/A VGND VGND VPWR VPWR _05449_/X sky130_fd_sc_hd__clkbuf_2
X_08237_ _08237_/A _08237_/B _08237_/C _08237_/D VGND VGND VPWR VPWR _08238_/D sky130_fd_sc_hd__and4_2
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08168_ _06881_/Y _08086_/X _06899_/Y _08087_/X _08167_/X VGND VGND VPWR VPWR _08171_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07119_ _09958_/Q VGND VGND VPWR VPWR _07119_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08099_ _08099_/A _08099_/B _08099_/C _08099_/D VGND VGND VPWR VPWR _08099_/Y sky130_fd_sc_hd__nand4_4
X_10130_ _10353_/CLK _10130_/D repeater403/X VGND VGND VPWR VPWR _10130_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10061_ _10062_/CLK _10061_/D repeater405/X VGND VGND VPWR VPWR _10061_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10157_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10310_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10510_/CLK _10328_/D _05034_/A VGND VGND VPWR VPWR _10328_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10290_/CLK _10259_/D repeater402/X VGND VGND VPWR VPWR _10259_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04820_ _09663_/X _05201_/C _05213_/B VGND VGND VPWR VPWR _05155_/A sky130_fd_sc_hd__or3_2
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07470_ _09797_/Q VGND VGND VPWR VPWR _07470_/Y sky130_fd_sc_hd__inv_2
X_06421_ _06417_/X _09625_/X _09650_/X _09887_/Q VGND VGND VPWR VPWR _09887_/D sky130_fd_sc_hd__o22a_1
XFILLER_61_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06352_ _06353_/A VGND VGND VPWR VPWR _06352_/X sky130_fd_sc_hd__clkbuf_2
X_09140_ _09273_/A _09384_/C _09140_/C VGND VGND VPWR VPWR _09142_/A sky130_fd_sc_hd__or3_1
X_06283_ _09973_/Q _06281_/X _09578_/X _06282_/Y VGND VGND VPWR VPWR _09973_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05303_ _05305_/A _05355_/A VGND VGND VPWR VPWR _05761_/A sky130_fd_sc_hd__or2_2
X_09071_ _09262_/A _09084_/B _08947_/A VGND VGND VPWR VPWR _09289_/C sky130_fd_sc_hd__o21ai_1
X_08022_ _05294_/Y _08188_/A _05308_/A _08189_/A VGND VGND VPWR VPWR _08022_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05234_ _07881_/A _06279_/A _05232_/Y _06303_/A VGND VGND VPWR VPWR _05234_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05165_ _05165_/A VGND VGND VPWR VPWR _09677_/S sky130_fd_sc_hd__buf_12
X_09973_ _10283_/CLK _09973_/D repeater406/X VGND VGND VPWR VPWR _09973_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05096_ _10451_/Q _05089_/X _10437_/Q _05091_/X _05095_/X VGND VGND VPWR VPWR _05108_/C
+ sky130_fd_sc_hd__a221o_1
X_08924_ _08938_/A _08927_/B VGND VGND VPWR VPWR _09370_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08855_ _08855_/A _09057_/B VGND VGND VPWR VPWR _09076_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08786_ _08786_/A _08786_/B VGND VGND VPWR VPWR _08864_/A sky130_fd_sc_hd__or2_1
X_07806_ _07806_/A VGND VGND VPWR VPWR _07806_/X sky130_fd_sc_hd__buf_2
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05998_ _10104_/Q _05994_/X _09576_/X _05995_/Y VGND VGND VPWR VPWR _10104_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07737_ _07016_/Y _07656_/X _06936_/Y _07657_/X _07736_/X VGND VGND VPWR VPWR _07743_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_169_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04949_ _09678_/X _04947_/Y _09536_/A3 _10471_/Q _04948_/X VGND VGND VPWR VPWR _10471_/D
+ sky130_fd_sc_hd__a32o_1
X_07668_ _07829_/A VGND VGND VPWR VPWR _07668_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09407_ _09407_/A _09407_/B _09407_/C _09407_/D VGND VGND VPWR VPWR _09439_/D sky130_fd_sc_hd__or4_1
XFILLER_111_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07599_ _05328_/Y _07532_/A _05241_/Y _07811_/A _07598_/X VGND VGND VPWR VPWR _07615_/A
+ sky130_fd_sc_hd__o221a_1
X_06619_ _06619_/A VGND VGND VPWR VPWR _06619_/X sky130_fd_sc_hd__clkbuf_1
X_09338_ _09109_/A _09336_/X _09048_/X _09337_/Y VGND VGND VPWR VPWR _09341_/B sky130_fd_sc_hd__o22ai_2
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09269_ _09269_/A VGND VGND VPWR VPWR _09400_/B sky130_fd_sc_hd__inv_2
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10113_ _10371_/CLK _10113_/D repeater405/X VGND VGND VPWR VPWR _10113_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10044_ _10404_/CLK _10044_/D repeater410/X VGND VGND VPWR VPWR _10044_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR net399_2/A
+ sky130_fd_sc_hd__clkbuf_2
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _07504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06970_ _09837_/Q VGND VGND VPWR VPWR _06970_/Y sky130_fd_sc_hd__clkinv_4
X_05921_ _10153_/Q _05919_/X _09578_/X _05920_/Y VGND VGND VPWR VPWR _10153_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08640_ _08640_/A _08781_/B VGND VGND VPWR VPWR _08645_/A sky130_fd_sc_hd__or2_4
X_05852_ _05896_/A _05852_/B VGND VGND VPWR VPWR _05854_/A sky130_fd_sc_hd__or2_2
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08571_ _08634_/B _08884_/A _08571_/C _08888_/A VGND VGND VPWR VPWR _09011_/A sky130_fd_sc_hd__or4_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05783_ _06679_/A VGND VGND VPWR VPWR _06327_/A sky130_fd_sc_hd__clkbuf_4
X_07522_ _07758_/A VGND VGND VPWR VPWR _07523_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07453_ _07453_/A VGND VGND VPWR VPWR _07453_/X sky130_fd_sc_hd__clkbuf_2
X_06404_ _06404_/A VGND VGND VPWR VPWR _06405_/A sky130_fd_sc_hd__inv_2
X_09123_ _09262_/A _09099_/X _09120_/X _09122_/Y VGND VGND VPWR VPWR _09123_/X sky130_fd_sc_hd__o211a_1
XFILLER_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07384_ _09948_/Q VGND VGND VPWR VPWR _07384_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06335_ _09942_/Q _06330_/X _06684_/B1 _06331_/Y VGND VGND VPWR VPWR _09942_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09054_ _09057_/B _09053_/X _08911_/X VGND VGND VPWR VPWR _09055_/B sky130_fd_sc_hd__o21a_1
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06266_ _06266_/A VGND VGND VPWR VPWR _06267_/B sky130_fd_sc_hd__buf_2
XFILLER_190_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05217_ _05336_/A _05355_/B VGND VGND VPWR VPWR _06266_/A sky130_fd_sc_hd__or2_4
X_08005_ _05265_/Y _08219_/A _05354_/Y _08220_/A _08004_/X VGND VGND VPWR VPWR _08050_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_150_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06197_ _10002_/Q VGND VGND VPWR VPWR _07994_/B sky130_fd_sc_hd__inv_2
XFILLER_171_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05148_ _05148_/A VGND VGND VPWR VPWR _05329_/A sky130_fd_sc_hd__buf_4
X_09956_ _10288_/CLK _09956_/D repeater406/X VGND VGND VPWR VPWR _09956_/Q sky130_fd_sc_hd__dfrtp_1
X_05079_ _06108_/B VGND VGND VPWR VPWR _05080_/A sky130_fd_sc_hd__inv_2
X_08907_ _09012_/A _08933_/A _09016_/D VGND VGND VPWR VPWR _08919_/B sky130_fd_sc_hd__o21ai_1
X_09887_ _10397_/CLK _09887_/D repeater409/X VGND VGND VPWR VPWR _09887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08838_ _08838_/A _09068_/A _09287_/A _09339_/B VGND VGND VPWR VPWR _08838_/X sky130_fd_sc_hd__or4_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater392 _09578_/X VGND VGND VPWR VPWR _09545_/A1 sky130_fd_sc_hd__buf_12
X_08769_ _08822_/B VGND VGND VPWR VPWR _08853_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput151 wb_adr_i[27] VGND VGND VPWR VPWR _06460_/A sky130_fd_sc_hd__clkbuf_1
Xinput140 wb_adr_i[17] VGND VGND VPWR VPWR _08399_/A sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_adr_i[8] VGND VGND VPWR VPWR _08405_/D sky130_fd_sc_hd__clkbuf_1
X_10027_ _10411_/CLK _10027_/D repeater407/X VGND VGND VPWR VPWR _10027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput184 wb_dat_i[27] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[17] VGND VGND VPWR VPWR _08359_/B sky130_fd_sc_hd__clkbuf_1
Xinput195 wb_dat_i[8] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06120_ _06327_/A VGND VGND VPWR VPWR _06304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06051_ _10072_/Q _06046_/X _06684_/B1 _06047_/Y VGND VGND VPWR VPWR _10072_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05002_ _10445_/Q _04995_/A _06683_/B1 _04996_/A VGND VGND VPWR VPWR _10445_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09810_ _10406_/CLK _09810_/D _06584_/X VGND VGND VPWR VPWR _09810_/Q sky130_fd_sc_hd__dfrtp_1
X_09741_ _09781_/CLK _09741_/D VGND VGND VPWR VPWR _09741_/Q sky130_fd_sc_hd__dfxtp_1
X_06953_ _06948_/Y _05728_/B _06949_/Y _06635_/B _06952_/X VGND VGND VPWR VPWR _06960_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05904_ _10162_/Q _05897_/X _09550_/A0 _05899_/X VGND VGND VPWR VPWR _10162_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06884_ _06882_/Y _06439_/B _06883_/Y _06291_/B VGND VGND VPWR VPWR _06884_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09672_ _09671_/X _10395_/Q _10299_/Q VGND VGND VPWR VPWR _09672_/X sky130_fd_sc_hd__mux2_2
X_08623_ _08766_/B VGND VGND VPWR VPWR _09145_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05835_ _10203_/Q _05831_/X _06683_/B1 _05832_/Y VGND VGND VPWR VPWR _10203_/D sky130_fd_sc_hd__a22o_1
X_05766_ _10244_/Q _05763_/X _09581_/X _05765_/X VGND VGND VPWR VPWR _10244_/D sky130_fd_sc_hd__a22o_1
X_08554_ _08490_/A _08546_/Y _08553_/X VGND VGND VPWR VPWR _08554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _07505_/A hold40/X VGND VGND VPWR VPWR _07505_/Y sky130_fd_sc_hd__nor2_2
X_08485_ _08485_/A _08492_/B _08492_/C VGND VGND VPWR VPWR _08905_/B sky130_fd_sc_hd__or3_4
X_05697_ _10284_/Q _05690_/X hold46/X _05692_/X VGND VGND VPWR VPWR _10284_/D sky130_fd_sc_hd__a22o_1
XFILLER_167_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07436_ _05367_/X _07427_/A _09750_/Q _07428_/A VGND VGND VPWR VPWR _09750_/D sky130_fd_sc_hd__o22a_1
X_07367_ _07362_/Y _06251_/B _07363_/Y _06290_/A _07366_/X VGND VGND VPWR VPWR _07374_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ _09104_/Y _09105_/Y _08815_/Y VGND VGND VPWR VPWR _09106_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06318_ _09953_/Q _06314_/X _09580_/X _06316_/X VGND VGND VPWR VPWR _09953_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09037_ _08999_/A _08385_/B _08980_/B _09036_/X VGND VGND VPWR VPWR _09038_/C sky130_fd_sc_hd__a31o_1
X_07298_ _10108_/Q VGND VGND VPWR VPWR _07298_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06249_ _09988_/Q _06203_/A _06245_/B _06147_/X VGND VGND VPWR VPWR _09988_/D sky130_fd_sc_hd__o22a_1
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09939_ _10310_/CLK _09939_/D repeater404/X VGND VGND VPWR VPWR _09939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _10513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05620_ _10326_/Q _05616_/X _06683_/B1 _05617_/Y VGND VGND VPWR VPWR _10326_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05551_ _05552_/A VGND VGND VPWR VPWR _05551_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05482_ _05497_/A VGND VGND VPWR VPWR _05483_/A sky130_fd_sc_hd__clkbuf_1
X_08270_ _07352_/Y _08205_/X _07343_/Y _08206_/X _08269_/X VGND VGND VPWR VPWR _08273_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07221_ _10400_/Q VGND VGND VPWR VPWR _07221_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_164_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07152_ _10368_/Q VGND VGND VPWR VPWR _07152_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06103_ _10041_/Q _06097_/X _09545_/A1 _06099_/X VGND VGND VPWR VPWR _10041_/D sky130_fd_sc_hd__a22o_1
X_07083_ _09972_/Q VGND VGND VPWR VPWR _07957_/A sky130_fd_sc_hd__inv_4
XFILLER_172_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06034_ _10082_/Q _06026_/A _06684_/B1 _06027_/A VGND VGND VPWR VPWR _10082_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07985_ _06964_/Y _07828_/A _07024_/Y _07829_/A VGND VGND VPWR VPWR _07985_/X sky130_fd_sc_hd__o22a_1
X_09724_ _10290_/Q _09501_/A VGND VGND VPWR VPWR _09724_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06936_ _10041_/Q VGND VGND VPWR VPWR _06936_/Y sky130_fd_sc_hd__clkinv_4
X_06867_ _07770_/A _06267_/B _06863_/Y _05808_/B _06866_/X VGND VGND VPWR VPWR _06880_/B
+ sky130_fd_sc_hd__o221a_1
X_09655_ _08352_/Y _09813_/Q _09770_/Q VGND VGND VPWR VPWR _09655_/X sky130_fd_sc_hd__mux2_1
X_05818_ _10212_/Q _05810_/A _09661_/A1 _05811_/A VGND VGND VPWR VPWR _10212_/D sky130_fd_sc_hd__a22o_1
X_08606_ _08457_/X _09218_/A _08605_/Y VGND VGND VPWR VPWR _08606_/X sky130_fd_sc_hd__o21ba_1
XFILLER_55_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09586_ _10310_/Q _09660_/A1 _09699_/S VGND VGND VPWR VPWR _09586_/X sky130_fd_sc_hd__mux2_1
X_06798_ _10349_/Q VGND VGND VPWR VPWR _06798_/Y sky130_fd_sc_hd__inv_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08537_ _08640_/A _08556_/B _08537_/C _09236_/A VGND VGND VPWR VPWR _08929_/A sky130_fd_sc_hd__or4_4
XFILLER_151_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05749_ _05794_/A _05749_/B VGND VGND VPWR VPWR _05751_/A sky130_fd_sc_hd__or2_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _09046_/A VGND VGND VPWR VPWR _08491_/C sky130_fd_sc_hd__inv_2
X_07419_ _07419_/A _07419_/B _07419_/C _07419_/D VGND VGND VPWR VPWR _07419_/X sky130_fd_sc_hd__and4_4
XFILLER_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08399_ _08399_/A _08399_/B _08399_/C _08399_/D VGND VGND VPWR VPWR _08641_/A sky130_fd_sc_hd__nand4_1
XFILLER_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _10471_/CLK _10430_/D repeater409/X VGND VGND VPWR VPWR _10430_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10361_ _10364_/CLK _10361_/D repeater410/X VGND VGND VPWR VPWR _10361_/Q sky130_fd_sc_hd__dfrtp_1
X_10292_ _10296_/CLK _10292_/D repeater402/X VGND VGND VPWR VPWR _10292_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07770_ _07770_/A _07770_/B VGND VGND VPWR VPWR _07770_/X sky130_fd_sc_hd__or2_1
X_04982_ _04982_/A VGND VGND VPWR VPWR _04982_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06721_ _06716_/Y _06154_/B _06717_/Y _06096_/B _06720_/X VGND VGND VPWR VPWR _06740_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09440_ _09440_/A VGND VGND VPWR VPWR _09440_/X sky130_fd_sc_hd__clkbuf_1
X_06652_ _06652_/A VGND VGND VPWR VPWR _06652_/X sky130_fd_sc_hd__clkbuf_1
X_09371_ _09371_/A _09371_/B _09371_/C _08560_/X VGND VGND VPWR VPWR _09439_/C sky130_fd_sc_hd__or4b_2
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06583_ _06591_/A VGND VGND VPWR VPWR _06584_/A sky130_fd_sc_hd__clkbuf_1
X_05603_ _05603_/A _05603_/B VGND VGND VPWR VPWR _05605_/A sky130_fd_sc_hd__or2_2
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08322_ _06974_/Y _08199_/A _06996_/Y _08200_/A _08321_/X VGND VGND VPWR VPWR _08327_/B
+ sky130_fd_sc_hd__o221a_1
X_05534_ _10375_/Q _05529_/X _09579_/X _05531_/X VGND VGND VPWR VPWR _10375_/D sky130_fd_sc_hd__a22o_1
X_08253_ _05208_/Y _08213_/X _05232_/Y _08214_/X VGND VGND VPWR VPWR _08253_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05465_ _05465_/A VGND VGND VPWR VPWR _05465_/X sky130_fd_sc_hd__clkbuf_1
X_07204_ _07202_/Y _05527_/A _07203_/Y _06329_/B VGND VGND VPWR VPWR _07204_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05396_ _05397_/A VGND VGND VPWR VPWR _05396_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08184_ _08184_/A VGND VGND VPWR VPWR _08184_/X sky130_fd_sc_hd__buf_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07135_ _10346_/Q VGND VGND VPWR VPWR _07135_/Y sky130_fd_sc_hd__clkinv_2
X_07066_ _10240_/Q VGND VGND VPWR VPWR _09509_/A sky130_fd_sc_hd__inv_4
XFILLER_161_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput230 _09512_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_06017_ _10094_/Q _06012_/X _09579_/X _06014_/X VGND VGND VPWR VPWR _10094_/D sky130_fd_sc_hd__a22o_1
Xoutput252 _09715_/Z VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput241 _09464_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput274 _09564_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_2
Xoutput263 _09725_/Z VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_2
Xoutput285 _09571_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_2
Xoutput296 _10469_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_2
XFILLER_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07968_ _06974_/Y _07627_/A _06955_/Y _07788_/A _07967_/X VGND VGND VPWR VPWR _07977_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09707_ _09707_/A _09467_/A VGND VGND VPWR VPWR _09707_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_74_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06919_ _10463_/Q _06689_/A input30/X _05129_/A VGND VGND VPWR VPWR _06919_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07899_ _07388_/Y _07806_/X _07414_/Y _07807_/X VGND VGND VPWR VPWR _07899_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09638_ _10426_/Q _06906_/X _09680_/S VGND VGND VPWR VPWR _09638_/X sky130_fd_sc_hd__mux2_1
X_09569_ _07504_/Y input90/X input76/X VGND VGND VPWR VPWR _09569_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10413_ _04807_/A1 _10413_/D _05414_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_1
XFILLER_139_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10344_ _10349_/CLK _10344_/D repeater404/X VGND VGND VPWR VPWR _10344_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10275_ _10405_/CLK _10275_/D repeater410/X VGND VGND VPWR VPWR _10275_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05250_ _05355_/A _05361_/B VGND VGND VPWR VPWR _06537_/A sky130_fd_sc_hd__or2_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05181_ _05336_/A _05139_/B _05179_/Y _05180_/Y _04915_/A VGND VGND VPWR VPWR _05181_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08940_ _09020_/A _08957_/B VGND VGND VPWR VPWR _09287_/B sky130_fd_sc_hd__nor2_1
X_08871_ _08996_/A _09271_/A _08871_/C VGND VGND VPWR VPWR _08872_/B sky130_fd_sc_hd__or3_1
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07822_ _07983_/B VGND VGND VPWR VPWR _07932_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07753_ _06857_/Y _07632_/X _06887_/Y _07633_/X _07752_/X VGND VGND VPWR VPWR _07761_/B
+ sky130_fd_sc_hd__o221a_2
X_04965_ _04993_/A _05085_/A VGND VGND VPWR VPWR _04967_/A sky130_fd_sc_hd__or2_2
X_04896_ _10489_/Q _04888_/A _09661_/A1 _04889_/A VGND VGND VPWR VPWR _10489_/D sky130_fd_sc_hd__a22o_1
X_07684_ _07684_/A _07684_/B _07684_/C _07684_/D VGND VGND VPWR VPWR _07695_/B sky130_fd_sc_hd__and4_1
X_06704_ _06704_/A VGND VGND VPWR VPWR _06704_/X sky130_fd_sc_hd__buf_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06635_ _06635_/A _06635_/B VGND VGND VPWR VPWR _06637_/A sky130_fd_sc_hd__or2_2
X_09423_ _09048_/X _09336_/X _08810_/B _09337_/Y _09422_/Y VGND VGND VPWR VPWR _09424_/B
+ sky130_fd_sc_hd__o221ai_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09354_ _09354_/A _09354_/B _09354_/C _09354_/D VGND VGND VPWR VPWR _09443_/A sky130_fd_sc_hd__or4_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08305_ _07151_/Y _08207_/A _07150_/Y _08208_/A VGND VGND VPWR VPWR _08305_/X sky130_fd_sc_hd__o22a_1
X_06566_ _09655_/X _09814_/Q _06575_/S VGND VGND VPWR VPWR _06567_/A sky130_fd_sc_hd__mux2_1
X_05517_ _05517_/A VGND VGND VPWR VPWR _10380_/D sky130_fd_sc_hd__clkbuf_1
X_06497_ _09853_/Q _06495_/X _09578_/X _06496_/Y VGND VGND VPWR VPWR _09853_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09285_ _09285_/A _09285_/B _09285_/C VGND VGND VPWR VPWR _09354_/D sky130_fd_sc_hd__or3_1
X_05448_ _09786_/Q _08356_/A VGND VGND VPWR VPWR _05450_/A sky130_fd_sc_hd__or2_4
XFILLER_176_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08236_ _06742_/Y _08211_/X _07854_/A _08212_/X _08235_/X VGND VGND VPWR VPWR _08237_/D
+ sky130_fd_sc_hd__o221a_1
X_08167_ _06864_/Y _08088_/X _06897_/Y _08089_/X VGND VGND VPWR VPWR _08167_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07118_ _09493_/A _05138_/A _09495_/A _05928_/B VGND VGND VPWR VPWR _07118_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05379_ _05379_/A VGND VGND VPWR VPWR _05379_/X sky130_fd_sc_hd__clkbuf_1
X_08098_ _08098_/A _08098_/B _08098_/C _08098_/D VGND VGND VPWR VPWR _08099_/D sky130_fd_sc_hd__and4_2
XFILLER_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_csclk clkbuf_leaf_7_csclk/A VGND VGND VPWR VPWR _10184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07049_ _10332_/Q VGND VGND VPWR VPWR _07049_/Y sky130_fd_sc_hd__inv_2
X_10060_ _10062_/CLK _10060_/D repeater405/X VGND VGND VPWR VPWR _10060_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10327_ _10336_/CLK _10327_/D repeater409/X VGND VGND VPWR VPWR _10327_/Q sky130_fd_sc_hd__dfstp_2
X_10258_ _10290_/CLK _10258_/D repeater402/X VGND VGND VPWR VPWR _10258_/Q sky130_fd_sc_hd__dfstp_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10189_ _10224_/CLK _10189_/D repeater405/X VGND VGND VPWR VPWR _10189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06420_ _06417_/X _09627_/X _09650_/X _09888_/Q VGND VGND VPWR VPWR _09888_/D sky130_fd_sc_hd__o22a_1
XFILLER_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06351_ _06472_/A _06351_/B VGND VGND VPWR VPWR _06353_/A sky130_fd_sc_hd__or2_2
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06282_ _06282_/A VGND VGND VPWR VPWR _06282_/Y sky130_fd_sc_hd__inv_2
X_05302_ _10237_/Q VGND VGND VPWR VPWR _05302_/Y sky130_fd_sc_hd__clkinv_4
X_09070_ _09070_/A _09442_/C _09287_/C _09070_/D VGND VGND VPWR VPWR _09074_/A sky130_fd_sc_hd__or4_1
XFILLER_147_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05233_ _05359_/A _05349_/B VGND VGND VPWR VPWR _06303_/A sky130_fd_sc_hd__or2_1
X_08021_ _08044_/A _08043_/B _08038_/C VGND VGND VPWR VPWR _08189_/A sky130_fd_sc_hd__or3_4
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05164_ _05318_/A _05164_/B VGND VGND VPWR VPWR _05165_/A sky130_fd_sc_hd__or2_1
X_09972_ _10283_/CLK _09972_/D repeater406/X VGND VGND VPWR VPWR _09972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05095_ _10467_/Q _04959_/Y _10107_/Q _05094_/Y VGND VGND VPWR VPWR _05095_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08923_ _08923_/A _08943_/A VGND VGND VPWR VPWR _09388_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08854_ _08854_/A _09357_/A VGND VGND VPWR VPWR _08856_/A sky130_fd_sc_hd__or2_1
X_05997_ _10105_/Q _05994_/X _09550_/A0 _05995_/Y VGND VGND VPWR VPWR _10105_/D sky130_fd_sc_hd__a22o_1
X_08785_ _09229_/A _09145_/B VGND VGND VPWR VPWR _09271_/A sky130_fd_sc_hd__nor2_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07805_ _07805_/A VGND VGND VPWR VPWR _07805_/X sky130_fd_sc_hd__buf_2
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_04948_ _05031_/A _04948_/B VGND VGND VPWR VPWR _04948_/X sky130_fd_sc_hd__or2_1
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07736_ _07003_/Y _07658_/X _07735_/Y _07659_/X VGND VGND VPWR VPWR _07736_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07667_ _07828_/A VGND VGND VPWR VPWR _07667_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04879_ _05651_/A VGND VGND VPWR VPWR _05806_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09406_ _09204_/A _08911_/X _09016_/D _08572_/X VGND VGND VPWR VPWR _09407_/B sky130_fd_sc_hd__o211ai_2
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07598_ _05221_/Y _07812_/A _05335_/Y _07653_/A VGND VGND VPWR VPWR _07598_/X sky130_fd_sc_hd__o22a_1
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06618_ _06666_/A VGND VGND VPWR VPWR _06619_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09337_ _09337_/A _09337_/B VGND VGND VPWR VPWR _09337_/Y sky130_fd_sc_hd__nor2_1
X_06549_ _09820_/Q _06540_/A _09659_/A1 _06541_/A VGND VGND VPWR VPWR _09820_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09268_ _09092_/A _08645_/A _09093_/A _08482_/A _09267_/Y VGND VGND VPWR VPWR _09269_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08219_ _08219_/A VGND VGND VPWR VPWR _08219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ _08527_/Y _09002_/Y _09379_/A _09075_/B VGND VGND VPWR VPWR _09311_/D sky130_fd_sc_hd__a211o_1
XFILLER_134_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10112_ _10482_/CLK _10112_/D repeater405/X VGND VGND VPWR VPWR _10112_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10043_ _10404_/CLK _10043_/D repeater410/X VGND VGND VPWR VPWR _10043_/Q sky130_fd_sc_hd__dfrtp_1
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_4 _05357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05920_ _05920_/A VGND VGND VPWR VPWR _05920_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05851_ _05851_/A VGND VGND VPWR VPWR _05852_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08570_ _08685_/B _08570_/B VGND VGND VPWR VPWR _08570_/X sky130_fd_sc_hd__or2_1
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05782_ _10232_/Q _05776_/X _09659_/A1 _05777_/Y VGND VGND VPWR VPWR _10232_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07521_ _07564_/C _07596_/B VGND VGND VPWR VPWR _07758_/A sky130_fd_sc_hd__or2_1
XFILLER_47_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07452_ _07452_/A VGND VGND VPWR VPWR _07453_/A sky130_fd_sc_hd__inv_2
XFILLER_62_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06403_ _06404_/A VGND VGND VPWR VPWR _06403_/X sky130_fd_sc_hd__clkbuf_2
X_07383_ _10051_/Q VGND VGND VPWR VPWR _07383_/Y sky130_fd_sc_hd__clkinv_4
X_06334_ _09943_/Q _06330_/X _06683_/B1 _06331_/Y VGND VGND VPWR VPWR _09943_/D sky130_fd_sc_hd__a22o_1
X_09122_ _09339_/C VGND VGND VPWR VPWR _09122_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09053_ _09083_/B _09056_/C VGND VGND VPWR VPWR _09053_/X sky130_fd_sc_hd__or2_1
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06265_ _06203_/Y _06259_/Y _06264_/Y _09982_/Q _06264_/A VGND VGND VPWR VPWR _09982_/D
+ sky130_fd_sc_hd__a32o_1
X_05216_ _09974_/Q VGND VGND VPWR VPWR _07606_/A sky130_fd_sc_hd__clkinv_2
X_08004_ _05184_/Y _08173_/A _05356_/Y _08174_/A VGND VGND VPWR VPWR _08004_/X sky130_fd_sc_hd__o22a_1
X_06196_ _10003_/Q VGND VGND VPWR VPWR _08046_/A sky130_fd_sc_hd__inv_2
X_05147_ _05142_/Y _05119_/Y _05144_/X _09766_/Q _05146_/Y VGND VGND VPWR VPWR _05183_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09955_ _10288_/CLK _09955_/D repeater406/X VGND VGND VPWR VPWR _09955_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05078_ _05160_/A _05100_/B VGND VGND VPWR VPWR _06108_/B sky130_fd_sc_hd__or2_1
X_08906_ _08911_/B _08906_/B VGND VGND VPWR VPWR _09016_/D sky130_fd_sc_hd__or2_2
XFILLER_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09886_ _09919_/CLK _09886_/D repeater409/X VGND VGND VPWR VPWR _09886_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _10283_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08837_ _08837_/A _08841_/B VGND VGND VPWR VPWR _09339_/B sky130_fd_sc_hd__nor2_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater393 _09578_/X VGND VGND VPWR VPWR _09547_/A1 sky130_fd_sc_hd__buf_12
X_08768_ _09085_/D _09102_/B _08768_/C VGND VGND VPWR VPWR _08822_/B sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_25_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _10491_/CLK sky130_fd_sc_hd__clkbuf_16
X_08699_ _08570_/B _08697_/B _08783_/A VGND VGND VPWR VPWR _08700_/D sky130_fd_sc_hd__a21oi_1
X_07719_ _06927_/Y _07622_/X _06937_/Y _07623_/X VGND VGND VPWR VPWR _07719_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput152 wb_adr_i[28] VGND VGND VPWR VPWR _06460_/B sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_adr_i[18] VGND VGND VPWR VPWR _08399_/D sky130_fd_sc_hd__clkbuf_1
Xinput130 usr2_vcc_pwrgood VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__buf_6
Xinput163 wb_adr_i[9] VGND VGND VPWR VPWR _08405_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10026_ _10411_/CLK _10026_/D repeater407/X VGND VGND VPWR VPWR _10026_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput185 wb_dat_i[28] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__clkbuf_1
Xinput174 wb_dat_i[18] VGND VGND VPWR VPWR _08361_/B sky130_fd_sc_hd__clkbuf_1
Xinput196 wb_dat_i[9] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06050_ _10073_/Q _06046_/X _06683_/B1 _06047_/Y VGND VGND VPWR VPWR _10073_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05001_ _10446_/Q _04994_/X _09658_/A1 _04996_/X VGND VGND VPWR VPWR _10446_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09740_ _09781_/CLK _09740_/D VGND VGND VPWR VPWR _09740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06952_ _06950_/Y _05851_/A _06951_/Y _05474_/B VGND VGND VPWR VPWR _06952_/X sky130_fd_sc_hd__o22a_2
.ends

