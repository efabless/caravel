magic
tech sky130A
timestamp 1638030917
<< viali >>
rect 1118 1572 1135 1589
rect 1348 1572 1365 1589
rect 1762 1572 1779 1589
rect 2222 1572 2239 1589
rect 2544 1572 2561 1589
rect 2682 1572 2699 1589
rect 2820 1572 2837 1589
rect 3004 1572 3021 1589
rect 3280 1572 3297 1589
rect 3418 1572 3435 1589
rect 3556 1572 3573 1589
rect 3694 1572 3711 1589
rect 3832 1572 3849 1589
rect 3970 1572 3987 1589
rect 4108 1572 4125 1589
rect 4246 1572 4263 1589
rect 4384 1572 4401 1589
rect 4568 1572 4585 1589
rect 4844 1572 4861 1589
rect 4982 1572 4999 1589
rect 5396 1572 5413 1589
rect 5672 1572 5689 1589
rect 6086 1572 6103 1589
rect 6362 1572 6379 1589
rect 6638 1572 6655 1589
rect 6776 1572 6793 1589
rect 6914 1572 6931 1589
rect 7190 1572 7207 1589
rect 7604 1572 7621 1589
rect 7880 1572 7897 1589
rect 8432 1572 8449 1589
rect 8846 1572 8863 1589
rect 9260 1572 9277 1589
rect 9720 1572 9737 1589
rect 10134 1572 10151 1589
rect 10686 1572 10703 1589
rect 11284 1572 11301 1589
rect 11836 1572 11853 1589
rect 12434 1572 12451 1589
rect 13124 1572 13141 1589
rect 13722 1572 13739 1589
rect 14274 1572 14291 1589
rect 14872 1572 14889 1589
rect 15424 1572 15441 1589
rect 15976 1572 15993 1589
rect 16436 1572 16453 1589
rect 16988 1572 17005 1589
rect 17586 1572 17603 1589
rect 18276 1572 18293 1589
rect 18874 1572 18891 1589
rect 19426 1572 19443 1589
rect 20024 1572 20041 1589
rect 20576 1572 20593 1589
rect 21312 1572 21329 1589
rect 21726 1572 21743 1589
rect 22140 1572 22157 1589
rect 22600 1572 22617 1589
rect 23888 1572 23905 1589
rect 24348 1572 24365 1589
rect 24486 1572 24503 1589
rect 24624 1572 24641 1589
rect 24762 1572 24779 1589
rect 24900 1572 24917 1589
rect 25176 1572 25193 1589
rect 25452 1572 25469 1589
rect 25590 1572 25607 1589
rect 25866 1572 25883 1589
rect 26142 1572 26159 1589
rect 26280 1572 26297 1589
rect 26602 1572 26619 1589
rect 26878 1572 26895 1589
rect 27016 1572 27033 1589
rect 27292 1572 27309 1589
rect 27568 1572 27585 1589
rect 27890 1572 27907 1589
rect 28304 1572 28321 1589
rect 28580 1572 28597 1589
rect 29040 1572 29057 1589
rect 29454 1572 29471 1589
rect 29868 1572 29885 1589
rect 30328 1572 30345 1589
rect 30604 1572 30621 1589
rect 31018 1572 31035 1589
rect 31294 1572 31311 1589
rect 31754 1572 31771 1589
rect 32582 1572 32599 1589
rect 33180 1572 33197 1589
rect 33318 1572 33335 1589
rect 33548 1572 33565 1589
rect 33686 1572 33703 1589
rect 33824 1572 33841 1589
rect 1486 1538 1503 1555
rect 8570 1538 8587 1555
rect 8984 1538 9001 1555
rect 9536 1538 9553 1555
rect 9996 1538 10013 1555
rect 10548 1538 10565 1555
rect 11146 1538 11163 1555
rect 11698 1538 11715 1555
rect 12112 1538 12129 1555
rect 12710 1538 12727 1555
rect 13584 1538 13601 1555
rect 14136 1538 14153 1555
rect 15010 1538 15027 1555
rect 15562 1538 15579 1555
rect 16160 1538 16177 1555
rect 16712 1538 16729 1555
rect 17264 1538 17281 1555
rect 18000 1538 18017 1555
rect 18736 1538 18753 1555
rect 19288 1538 19305 1555
rect 19840 1538 19857 1555
rect 20438 1538 20455 1555
rect 21450 1538 21467 1555
rect 22002 1538 22019 1555
rect 22738 1538 22755 1555
rect 25314 1538 25331 1555
rect 26004 1538 26021 1555
rect 26740 1538 26757 1555
rect 27154 1538 27171 1555
rect 27430 1538 27447 1555
rect 27752 1538 27769 1555
rect 28718 1538 28735 1555
rect 29178 1538 29195 1555
rect 29592 1538 29609 1555
rect 30006 1538 30023 1555
rect 30466 1538 30483 1555
rect 30880 1538 30897 1555
rect 31432 1538 31449 1555
rect 31892 1538 31909 1555
rect 32444 1538 32461 1555
rect 33042 1538 33059 1555
rect 1532 1504 1549 1521
rect 4706 1504 4723 1521
rect 5258 1504 5275 1521
rect 5534 1504 5551 1521
rect 5856 1504 5873 1521
rect 6224 1504 6241 1521
rect 6500 1504 6517 1521
rect 7466 1504 7483 1521
rect 7742 1504 7759 1521
rect 8018 1504 8035 1521
rect 8708 1504 8725 1521
rect 9122 1504 9139 1521
rect 9858 1504 9875 1521
rect 10410 1504 10427 1521
rect 11008 1504 11025 1521
rect 11422 1504 11439 1521
rect 11974 1504 11991 1521
rect 12572 1504 12589 1521
rect 13262 1504 13279 1521
rect 13860 1504 13877 1521
rect 14412 1504 14429 1521
rect 15148 1504 15165 1521
rect 15700 1504 15717 1521
rect 16298 1504 16315 1521
rect 16850 1504 16867 1521
rect 17448 1504 17465 1521
rect 18138 1504 18155 1521
rect 18414 1504 18431 1521
rect 19012 1504 19029 1521
rect 19564 1504 19581 1521
rect 20162 1504 20179 1521
rect 20714 1504 20731 1521
rect 21128 1504 21145 1521
rect 21588 1504 21605 1521
rect 22278 1504 22295 1521
rect 22876 1504 22893 1521
rect 24026 1504 24043 1521
rect 25728 1504 25745 1521
rect 26464 1504 26481 1521
rect 28166 1504 28183 1521
rect 28442 1504 28459 1521
rect 28856 1504 28873 1521
rect 29316 1504 29333 1521
rect 29730 1504 29747 1521
rect 30144 1504 30161 1521
rect 30742 1504 30759 1521
rect 31156 1504 31173 1521
rect 31616 1504 31633 1521
rect 32168 1504 32185 1521
rect 32720 1504 32737 1521
rect 32996 1504 33013 1521
rect 1808 1470 1825 1487
rect 2084 1470 2101 1487
rect 2360 1470 2377 1487
rect 5120 1470 5137 1487
rect 7328 1470 7345 1487
rect 8156 1470 8173 1487
rect 9398 1470 9415 1487
rect 10272 1470 10289 1487
rect 10824 1470 10841 1487
rect 11560 1470 11577 1487
rect 12296 1470 12313 1487
rect 12848 1470 12865 1487
rect 12986 1470 13003 1487
rect 13400 1470 13417 1487
rect 13998 1470 14015 1487
rect 14550 1470 14567 1487
rect 14688 1470 14705 1487
rect 15286 1470 15303 1487
rect 15838 1470 15855 1487
rect 16574 1470 16591 1487
rect 17126 1470 17143 1487
rect 17724 1470 17741 1487
rect 17862 1470 17879 1487
rect 18552 1470 18569 1487
rect 19150 1470 19167 1487
rect 19702 1470 19719 1487
rect 20300 1470 20317 1487
rect 20852 1470 20869 1487
rect 20990 1470 21007 1487
rect 21864 1470 21881 1487
rect 22416 1470 22433 1487
rect 28028 1470 28045 1487
rect 32030 1470 32047 1487
rect 32306 1470 32323 1487
rect 1394 1232 1411 1249
rect 1762 1232 1779 1249
rect 2084 1232 2101 1249
rect 2636 1232 2653 1249
rect 3142 1232 3159 1249
rect 5948 1232 5965 1249
rect 14412 1232 14429 1249
rect 18276 1232 18293 1249
rect 20852 1232 20869 1249
rect 22140 1232 22157 1249
rect 22646 1232 22663 1249
rect 22784 1232 22801 1249
rect 22922 1232 22939 1249
rect 23060 1232 23077 1249
rect 23198 1232 23215 1249
rect 23336 1232 23353 1249
rect 23474 1232 23491 1249
rect 23612 1232 23629 1249
rect 24026 1232 24043 1249
rect 24164 1232 24181 1249
rect 32490 1232 32507 1249
rect 32720 1232 32737 1249
rect 32996 1232 33013 1249
rect 33134 1232 33151 1249
rect 33272 1232 33289 1249
rect 1532 1198 1549 1215
rect 2774 1198 2791 1215
rect 3280 1198 3297 1215
rect 2222 1164 2239 1181
rect 2498 1164 2515 1181
rect 1256 1130 1273 1147
rect 1808 1130 1825 1147
rect 2360 1130 2377 1147
rect 2912 1130 2929 1147
rect 1072 1028 1089 1045
rect 1946 1028 1963 1045
rect 2084 1028 2101 1045
rect 3280 1028 3297 1045
rect 3418 1028 3435 1045
rect 2222 994 2239 1011
rect 2912 994 2929 1011
rect 1118 960 1135 977
rect 2360 960 2377 977
rect 3050 960 3067 977
rect 23060 960 23077 977
rect 1348 926 1365 943
rect 1394 926 1411 943
rect 1532 926 1549 943
rect 1670 926 1687 943
rect 1808 926 1825 943
rect 2498 926 2515 943
rect 2636 926 2653 943
rect 2774 926 2791 943
rect 3648 926 3665 943
rect 4936 926 4953 943
rect 6086 926 6103 943
rect 7052 926 7069 943
rect 8432 926 8449 943
rect 10134 926 10151 943
rect 11100 926 11117 943
rect 12526 926 12543 943
rect 14642 926 14659 943
rect 15746 926 15763 943
rect 16298 926 16315 943
rect 22186 926 22203 943
rect 22784 926 22801 943
rect 26142 926 26159 943
rect 13906 688 13923 705
rect 20208 688 20225 705
rect 23474 688 23491 705
rect 26142 688 26159 705
rect 1072 654 1089 671
rect 1532 654 1549 671
rect 2360 654 2377 671
rect 2774 654 2791 671
rect 2912 654 2929 671
rect 3602 654 3619 671
rect 3924 654 3941 671
rect 5074 654 5091 671
rect 5994 654 6011 671
rect 6776 654 6793 671
rect 7190 654 7207 671
rect 8156 654 8173 671
rect 8754 654 8771 671
rect 9168 654 9185 671
rect 9996 654 10013 671
rect 10410 654 10427 671
rect 10824 654 10841 671
rect 11514 654 11531 671
rect 12112 654 12129 671
rect 12802 654 12819 671
rect 13354 654 13371 671
rect 14044 654 14061 671
rect 14596 654 14613 671
rect 15194 654 15211 671
rect 15884 654 15901 671
rect 16574 654 16591 671
rect 16988 654 17005 671
rect 17448 654 17465 671
rect 17724 654 17741 671
rect 18276 654 18293 671
rect 18736 654 18753 671
rect 19150 654 19167 671
rect 19564 654 19581 671
rect 20346 654 20363 671
rect 20898 654 20915 671
rect 21450 654 21467 671
rect 22186 654 22203 671
rect 22600 654 22617 671
rect 23198 654 23215 671
rect 23888 654 23905 671
rect 24302 654 24319 671
rect 24854 654 24871 671
rect 25176 654 25193 671
rect 25590 654 25607 671
rect 26464 654 26481 671
rect 27016 654 27033 671
rect 27890 654 27907 671
rect 1256 620 1273 637
rect 2222 620 2239 637
rect 3050 620 3067 637
rect 3464 620 3481 637
rect 4062 620 4079 637
rect 4384 620 4401 637
rect 4706 620 4723 637
rect 5350 620 5367 637
rect 5626 620 5643 637
rect 6224 620 6241 637
rect 6638 620 6655 637
rect 7328 620 7345 637
rect 7604 620 7621 637
rect 8616 620 8633 637
rect 9306 620 9323 637
rect 9858 620 9875 637
rect 10272 620 10289 637
rect 10686 620 10703 637
rect 11238 620 11255 637
rect 11790 620 11807 637
rect 12296 620 12313 637
rect 12664 620 12681 637
rect 13216 620 13233 637
rect 13768 620 13785 637
rect 14458 620 14475 637
rect 14918 620 14935 637
rect 15332 620 15349 637
rect 15608 620 15625 637
rect 16436 620 16453 637
rect 16850 620 16867 637
rect 17264 620 17281 637
rect 18138 620 18155 637
rect 18552 620 18569 637
rect 19012 620 19029 637
rect 19426 620 19443 637
rect 20070 620 20087 637
rect 20484 620 20501 637
rect 20760 620 20777 637
rect 21772 620 21789 637
rect 22922 620 22939 637
rect 23336 620 23353 637
rect 23612 620 23629 637
rect 24164 620 24181 637
rect 24716 620 24733 637
rect 25314 620 25331 637
rect 26280 620 26297 637
rect 26740 620 26757 637
rect 27154 620 27171 637
rect 27430 620 27447 637
rect 28028 620 28045 637
rect 934 586 951 603
rect 1210 586 1227 603
rect 1394 586 1411 603
rect 1670 586 1687 603
rect 1808 586 1825 603
rect 2084 586 2101 603
rect 2498 586 2515 603
rect 2636 586 2653 603
rect 3326 586 3343 603
rect 3786 586 3803 603
rect 4246 586 4263 603
rect 4568 586 4585 603
rect 4844 586 4861 603
rect 5212 586 5229 603
rect 5488 586 5505 603
rect 5856 586 5873 603
rect 6362 586 6379 603
rect 6500 586 6517 603
rect 6914 586 6931 603
rect 7466 586 7483 603
rect 7742 586 7759 603
rect 7880 586 7897 603
rect 8018 586 8035 603
rect 8432 586 8449 603
rect 8892 586 8909 603
rect 9030 586 9047 603
rect 9444 586 9461 603
rect 9720 586 9737 603
rect 10134 586 10151 603
rect 10548 586 10565 603
rect 11008 586 11025 603
rect 11376 586 11393 603
rect 11652 586 11669 603
rect 11974 586 11991 603
rect 12434 586 12451 603
rect 12940 586 12957 603
rect 13078 586 13095 603
rect 13584 586 13601 603
rect 14182 586 14199 603
rect 14320 586 14337 603
rect 15056 586 15073 603
rect 15470 586 15487 603
rect 15746 586 15763 603
rect 16160 586 16177 603
rect 16298 586 16315 603
rect 16712 586 16729 603
rect 17126 586 17143 603
rect 17586 586 17603 603
rect 17862 586 17879 603
rect 18000 586 18017 603
rect 18414 586 18431 603
rect 18874 586 18891 603
rect 19288 586 19305 603
rect 19702 586 19719 603
rect 19840 586 19857 603
rect 20622 586 20639 603
rect 21036 586 21053 603
rect 21312 586 21329 603
rect 21588 586 21605 603
rect 21910 586 21927 603
rect 22048 586 22065 603
rect 22324 586 22341 603
rect 22738 586 22755 603
rect 23060 586 23077 603
rect 24026 586 24043 603
rect 24440 586 24457 603
rect 24578 586 24595 603
rect 24992 586 25009 603
rect 25452 586 25469 603
rect 25728 586 25745 603
rect 25866 586 25883 603
rect 26004 586 26021 603
rect 26602 586 26619 603
rect 26878 586 26895 603
rect 27292 586 27309 603
rect 27568 586 27585 603
rect 27752 586 27769 603
rect 28166 586 28183 603
<< metal1 >>
rect 329 1704 332 1730
rect 358 1724 361 1730
rect 3411 1724 3414 1730
rect 358 1710 3414 1724
rect 358 1704 361 1710
rect 3411 1704 3414 1710
rect 3440 1704 3443 1730
rect 835 1670 838 1696
rect 864 1690 867 1696
rect 2951 1690 2954 1696
rect 864 1676 2954 1690
rect 864 1670 867 1676
rect 2951 1670 2954 1676
rect 2980 1670 2983 1696
rect 12427 1670 12430 1696
rect 12456 1690 12459 1696
rect 12933 1690 12936 1696
rect 12456 1676 12936 1690
rect 12456 1670 12459 1676
rect 12933 1670 12936 1676
rect 12962 1670 12965 1696
rect 644 1645 34408 1656
rect 644 1619 6631 1645
rect 6657 1619 12631 1645
rect 12657 1619 18631 1645
rect 18657 1619 24631 1645
rect 24657 1619 30631 1645
rect 30657 1619 34408 1645
rect 644 1608 34408 1619
rect 697 1568 700 1594
rect 726 1588 729 1594
rect 1112 1589 1141 1592
rect 1112 1588 1118 1589
rect 726 1574 1118 1588
rect 726 1568 729 1574
rect 1112 1572 1118 1574
rect 1135 1572 1141 1589
rect 1112 1569 1141 1572
rect 1342 1589 1371 1592
rect 1342 1572 1348 1589
rect 1365 1588 1371 1589
rect 1663 1588 1666 1594
rect 1365 1574 1666 1588
rect 1365 1572 1371 1574
rect 1342 1569 1371 1572
rect 1663 1568 1666 1574
rect 1692 1568 1695 1594
rect 1756 1589 1785 1592
rect 1756 1572 1762 1589
rect 1779 1588 1785 1589
rect 1801 1588 1804 1594
rect 1779 1574 1804 1588
rect 1779 1572 1785 1574
rect 1756 1569 1785 1572
rect 1801 1568 1804 1574
rect 1830 1568 1833 1594
rect 2031 1568 2034 1594
rect 2060 1588 2063 1594
rect 2216 1589 2245 1592
rect 2216 1588 2222 1589
rect 2060 1574 2222 1588
rect 2060 1568 2063 1574
rect 2216 1572 2222 1574
rect 2239 1572 2245 1589
rect 2216 1569 2245 1572
rect 2491 1568 2494 1594
rect 2520 1588 2523 1594
rect 2538 1589 2567 1592
rect 2538 1588 2544 1589
rect 2520 1574 2544 1588
rect 2520 1568 2523 1574
rect 2538 1572 2544 1574
rect 2561 1572 2567 1589
rect 2538 1569 2567 1572
rect 2629 1568 2632 1594
rect 2658 1588 2661 1594
rect 2676 1589 2705 1592
rect 2676 1588 2682 1589
rect 2658 1574 2682 1588
rect 2658 1568 2661 1574
rect 2676 1572 2682 1574
rect 2699 1572 2705 1589
rect 2676 1569 2705 1572
rect 2767 1568 2770 1594
rect 2796 1588 2799 1594
rect 2814 1589 2843 1592
rect 2814 1588 2820 1589
rect 2796 1574 2820 1588
rect 2796 1568 2799 1574
rect 2814 1572 2820 1574
rect 2837 1572 2843 1589
rect 2814 1569 2843 1572
rect 2905 1568 2908 1594
rect 2934 1588 2937 1594
rect 2998 1589 3027 1592
rect 2998 1588 3004 1589
rect 2934 1574 3004 1588
rect 2934 1568 2937 1574
rect 2998 1572 3004 1574
rect 3021 1572 3027 1589
rect 2998 1569 3027 1572
rect 3181 1568 3184 1594
rect 3210 1588 3213 1594
rect 3274 1589 3303 1592
rect 3274 1588 3280 1589
rect 3210 1574 3280 1588
rect 3210 1568 3213 1574
rect 3274 1572 3280 1574
rect 3297 1572 3303 1589
rect 3274 1569 3303 1572
rect 3319 1568 3322 1594
rect 3348 1588 3351 1594
rect 3412 1589 3441 1592
rect 3412 1588 3418 1589
rect 3348 1574 3418 1588
rect 3348 1568 3351 1574
rect 3412 1572 3418 1574
rect 3435 1572 3441 1589
rect 3412 1569 3441 1572
rect 3457 1568 3460 1594
rect 3486 1588 3489 1594
rect 3550 1589 3579 1592
rect 3550 1588 3556 1589
rect 3486 1574 3556 1588
rect 3486 1568 3489 1574
rect 3550 1572 3556 1574
rect 3573 1572 3579 1589
rect 3687 1588 3690 1594
rect 3667 1574 3690 1588
rect 3550 1569 3579 1572
rect 3687 1568 3690 1574
rect 3716 1568 3719 1594
rect 3733 1568 3736 1594
rect 3762 1588 3765 1594
rect 3826 1589 3855 1592
rect 3826 1588 3832 1589
rect 3762 1574 3832 1588
rect 3762 1568 3765 1574
rect 3826 1572 3832 1574
rect 3849 1572 3855 1589
rect 3826 1569 3855 1572
rect 3871 1568 3874 1594
rect 3900 1588 3903 1594
rect 3964 1589 3993 1592
rect 3964 1588 3970 1589
rect 3900 1574 3970 1588
rect 3900 1568 3903 1574
rect 3964 1572 3970 1574
rect 3987 1572 3993 1589
rect 3964 1569 3993 1572
rect 4009 1568 4012 1594
rect 4038 1588 4041 1594
rect 4102 1589 4131 1592
rect 4102 1588 4108 1589
rect 4038 1574 4108 1588
rect 4038 1568 4041 1574
rect 4102 1572 4108 1574
rect 4125 1572 4131 1589
rect 4102 1569 4131 1572
rect 4147 1568 4150 1594
rect 4176 1588 4179 1594
rect 4240 1589 4269 1592
rect 4240 1588 4246 1589
rect 4176 1574 4246 1588
rect 4176 1568 4179 1574
rect 4240 1572 4246 1574
rect 4263 1572 4269 1589
rect 4240 1569 4269 1572
rect 4285 1568 4288 1594
rect 4314 1588 4317 1594
rect 4378 1589 4407 1592
rect 4378 1588 4384 1589
rect 4314 1574 4384 1588
rect 4314 1568 4317 1574
rect 4378 1572 4384 1574
rect 4401 1572 4407 1589
rect 4378 1569 4407 1572
rect 4423 1568 4426 1594
rect 4452 1588 4455 1594
rect 4562 1589 4591 1592
rect 4562 1588 4568 1589
rect 4452 1574 4568 1588
rect 4452 1568 4455 1574
rect 4562 1572 4568 1574
rect 4585 1572 4591 1589
rect 4837 1588 4840 1594
rect 4817 1574 4840 1588
rect 4562 1569 4591 1572
rect 4837 1568 4840 1574
rect 4866 1568 4869 1594
rect 4883 1568 4886 1594
rect 4912 1588 4915 1594
rect 4976 1589 5005 1592
rect 4976 1588 4982 1589
rect 4912 1574 4982 1588
rect 4912 1568 4915 1574
rect 4976 1572 4982 1574
rect 4999 1572 5005 1589
rect 4976 1569 5005 1572
rect 5251 1568 5254 1594
rect 5280 1588 5283 1594
rect 5390 1589 5419 1592
rect 5390 1588 5396 1589
rect 5280 1574 5396 1588
rect 5280 1568 5283 1574
rect 5390 1572 5396 1574
rect 5413 1572 5419 1589
rect 5390 1569 5419 1572
rect 5527 1568 5530 1594
rect 5556 1588 5559 1594
rect 5666 1589 5695 1592
rect 5666 1588 5672 1589
rect 5556 1574 5672 1588
rect 5556 1568 5559 1574
rect 5666 1572 5672 1574
rect 5689 1572 5695 1589
rect 5666 1569 5695 1572
rect 5941 1568 5944 1594
rect 5970 1588 5973 1594
rect 6080 1589 6109 1592
rect 6080 1588 6086 1589
rect 5970 1574 6086 1588
rect 5970 1568 5973 1574
rect 6080 1572 6086 1574
rect 6103 1572 6109 1589
rect 6080 1569 6109 1572
rect 6217 1568 6220 1594
rect 6246 1588 6249 1594
rect 6356 1589 6385 1592
rect 6356 1588 6362 1589
rect 6246 1574 6362 1588
rect 6246 1568 6249 1574
rect 6356 1572 6362 1574
rect 6379 1572 6385 1589
rect 6356 1569 6385 1572
rect 6493 1568 6496 1594
rect 6522 1588 6525 1594
rect 6632 1589 6661 1592
rect 6632 1588 6638 1589
rect 6522 1574 6638 1588
rect 6522 1568 6525 1574
rect 6632 1572 6638 1574
rect 6655 1572 6661 1589
rect 6632 1569 6661 1572
rect 6723 1568 6726 1594
rect 6752 1588 6755 1594
rect 6770 1589 6799 1592
rect 6770 1588 6776 1589
rect 6752 1574 6776 1588
rect 6752 1568 6755 1574
rect 6770 1572 6776 1574
rect 6793 1572 6799 1589
rect 6907 1588 6910 1594
rect 6887 1574 6910 1588
rect 6770 1569 6799 1572
rect 6907 1568 6910 1574
rect 6936 1568 6939 1594
rect 7045 1568 7048 1594
rect 7074 1588 7077 1594
rect 7184 1589 7213 1592
rect 7184 1588 7190 1589
rect 7074 1574 7190 1588
rect 7074 1568 7077 1574
rect 7184 1572 7190 1574
rect 7207 1572 7213 1589
rect 7184 1569 7213 1572
rect 7321 1568 7324 1594
rect 7350 1588 7353 1594
rect 7598 1589 7627 1592
rect 7598 1588 7604 1589
rect 7350 1574 7604 1588
rect 7350 1568 7353 1574
rect 7598 1572 7604 1574
rect 7621 1572 7627 1589
rect 7598 1569 7627 1572
rect 7643 1568 7646 1594
rect 7672 1588 7675 1594
rect 7874 1589 7903 1592
rect 7874 1588 7880 1589
rect 7672 1574 7880 1588
rect 7672 1568 7675 1574
rect 7874 1572 7880 1574
rect 7897 1572 7903 1589
rect 7874 1569 7903 1572
rect 8011 1568 8014 1594
rect 8040 1588 8043 1594
rect 8426 1589 8455 1592
rect 8426 1588 8432 1589
rect 8040 1574 8432 1588
rect 8040 1568 8043 1574
rect 8426 1572 8432 1574
rect 8449 1572 8455 1589
rect 8426 1569 8455 1572
rect 8471 1568 8474 1594
rect 8500 1588 8503 1594
rect 8840 1589 8869 1592
rect 8840 1588 8846 1589
rect 8500 1574 8846 1588
rect 8500 1568 8503 1574
rect 8840 1572 8846 1574
rect 8863 1572 8869 1589
rect 8840 1569 8869 1572
rect 8885 1568 8888 1594
rect 8914 1588 8917 1594
rect 9254 1589 9283 1592
rect 9254 1588 9260 1589
rect 8914 1574 9260 1588
rect 8914 1568 8917 1574
rect 9254 1572 9260 1574
rect 9277 1572 9283 1589
rect 9254 1569 9283 1572
rect 9299 1568 9302 1594
rect 9328 1588 9331 1594
rect 9714 1589 9743 1592
rect 9714 1588 9720 1589
rect 9328 1574 9720 1588
rect 9328 1568 9331 1574
rect 9714 1572 9720 1574
rect 9737 1572 9743 1589
rect 9714 1569 9743 1572
rect 9759 1568 9762 1594
rect 9788 1588 9791 1594
rect 10128 1589 10157 1592
rect 10128 1588 10134 1589
rect 9788 1574 10134 1588
rect 9788 1568 9791 1574
rect 10128 1572 10134 1574
rect 10151 1572 10157 1589
rect 10128 1569 10157 1572
rect 10219 1568 10222 1594
rect 10248 1588 10251 1594
rect 10680 1589 10709 1592
rect 10680 1588 10686 1589
rect 10248 1574 10686 1588
rect 10248 1568 10251 1574
rect 10680 1572 10686 1574
rect 10703 1572 10709 1589
rect 10680 1569 10709 1572
rect 10771 1568 10774 1594
rect 10800 1588 10803 1594
rect 11278 1589 11307 1592
rect 11278 1588 11284 1589
rect 10800 1574 11284 1588
rect 10800 1568 10803 1574
rect 11278 1572 11284 1574
rect 11301 1572 11307 1589
rect 11278 1569 11307 1572
rect 11323 1568 11326 1594
rect 11352 1588 11355 1594
rect 11830 1589 11859 1592
rect 11830 1588 11836 1589
rect 11352 1574 11836 1588
rect 11352 1568 11355 1574
rect 11830 1572 11836 1574
rect 11853 1572 11859 1589
rect 11830 1569 11859 1572
rect 11875 1568 11878 1594
rect 11904 1588 11907 1594
rect 12428 1589 12457 1592
rect 12428 1588 12434 1589
rect 11904 1574 12434 1588
rect 11904 1568 11907 1574
rect 12428 1572 12434 1574
rect 12451 1572 12457 1589
rect 12428 1569 12457 1572
rect 12565 1568 12568 1594
rect 12594 1588 12597 1594
rect 13118 1589 13147 1592
rect 13118 1588 13124 1589
rect 12594 1574 13124 1588
rect 12594 1568 12597 1574
rect 13118 1572 13124 1574
rect 13141 1572 13147 1589
rect 13118 1569 13147 1572
rect 13163 1568 13166 1594
rect 13192 1588 13195 1594
rect 13716 1589 13745 1592
rect 13716 1588 13722 1589
rect 13192 1574 13722 1588
rect 13192 1568 13195 1574
rect 13716 1572 13722 1574
rect 13739 1572 13745 1589
rect 13716 1569 13745 1572
rect 13807 1568 13810 1594
rect 13836 1588 13839 1594
rect 14268 1589 14297 1592
rect 14268 1588 14274 1589
rect 13836 1574 14274 1588
rect 13836 1568 13839 1574
rect 14268 1572 14274 1574
rect 14291 1572 14297 1589
rect 14268 1569 14297 1572
rect 14359 1568 14362 1594
rect 14388 1588 14391 1594
rect 14866 1589 14895 1592
rect 14866 1588 14872 1589
rect 14388 1574 14872 1588
rect 14388 1568 14391 1574
rect 14866 1572 14872 1574
rect 14889 1572 14895 1589
rect 14866 1569 14895 1572
rect 14911 1568 14914 1594
rect 14940 1588 14943 1594
rect 15418 1589 15447 1592
rect 15418 1588 15424 1589
rect 14940 1574 15424 1588
rect 14940 1568 14943 1574
rect 15418 1572 15424 1574
rect 15441 1572 15447 1589
rect 15418 1569 15447 1572
rect 15463 1568 15466 1594
rect 15492 1588 15495 1594
rect 15970 1589 15999 1592
rect 15970 1588 15976 1589
rect 15492 1574 15976 1588
rect 15492 1568 15495 1574
rect 15970 1572 15976 1574
rect 15993 1572 15999 1589
rect 15970 1569 15999 1572
rect 16015 1568 16018 1594
rect 16044 1588 16047 1594
rect 16430 1589 16459 1592
rect 16430 1588 16436 1589
rect 16044 1574 16436 1588
rect 16044 1568 16047 1574
rect 16430 1572 16436 1574
rect 16453 1572 16459 1589
rect 16430 1569 16459 1572
rect 16567 1568 16570 1594
rect 16596 1588 16599 1594
rect 16982 1589 17011 1592
rect 16982 1588 16988 1589
rect 16596 1574 16988 1588
rect 16596 1568 16599 1574
rect 16982 1572 16988 1574
rect 17005 1572 17011 1589
rect 16982 1569 17011 1572
rect 17027 1568 17030 1594
rect 17056 1588 17059 1594
rect 17580 1589 17609 1592
rect 17580 1588 17586 1589
rect 17056 1574 17586 1588
rect 17056 1568 17059 1574
rect 17580 1572 17586 1574
rect 17603 1572 17609 1589
rect 17580 1569 17609 1572
rect 17671 1568 17674 1594
rect 17700 1588 17703 1594
rect 18270 1589 18299 1592
rect 18270 1588 18276 1589
rect 17700 1574 18276 1588
rect 17700 1568 17703 1574
rect 18270 1572 18276 1574
rect 18293 1572 18299 1589
rect 18270 1569 18299 1572
rect 18361 1568 18364 1594
rect 18390 1588 18393 1594
rect 18868 1589 18897 1592
rect 18868 1588 18874 1589
rect 18390 1574 18874 1588
rect 18390 1568 18393 1574
rect 18868 1572 18874 1574
rect 18891 1572 18897 1589
rect 18868 1569 18897 1572
rect 18913 1568 18916 1594
rect 18942 1588 18945 1594
rect 19420 1589 19449 1592
rect 19420 1588 19426 1589
rect 18942 1574 19426 1588
rect 18942 1568 18945 1574
rect 19420 1572 19426 1574
rect 19443 1572 19449 1589
rect 19420 1569 19449 1572
rect 19465 1568 19468 1594
rect 19494 1588 19497 1594
rect 20018 1589 20047 1592
rect 20018 1588 20024 1589
rect 19494 1574 20024 1588
rect 19494 1568 19497 1574
rect 20018 1572 20024 1574
rect 20041 1572 20047 1589
rect 20018 1569 20047 1572
rect 20063 1568 20066 1594
rect 20092 1588 20095 1594
rect 20570 1589 20599 1592
rect 20570 1588 20576 1589
rect 20092 1574 20576 1588
rect 20092 1568 20095 1574
rect 20570 1572 20576 1574
rect 20593 1572 20599 1589
rect 20570 1569 20599 1572
rect 20615 1568 20618 1594
rect 20644 1588 20647 1594
rect 20644 1574 20822 1588
rect 20644 1568 20647 1574
rect 1480 1555 1509 1558
rect 1480 1538 1486 1555
rect 1503 1554 1509 1555
rect 2077 1554 2080 1560
rect 1503 1540 2080 1554
rect 1503 1538 1509 1540
rect 1480 1535 1509 1538
rect 2077 1534 2080 1540
rect 2106 1534 2109 1560
rect 5113 1534 5116 1560
rect 5142 1554 5145 1560
rect 5142 1540 5274 1554
rect 5142 1534 5145 1540
rect 145 1500 148 1526
rect 174 1520 177 1526
rect 1526 1521 1555 1524
rect 1526 1520 1532 1521
rect 174 1506 1532 1520
rect 174 1500 177 1506
rect 1526 1504 1532 1506
rect 1549 1504 1555 1521
rect 1526 1501 1555 1504
rect 4561 1500 4564 1526
rect 4590 1520 4593 1526
rect 5260 1524 5274 1540
rect 8287 1534 8290 1560
rect 8316 1554 8319 1560
rect 8564 1555 8593 1558
rect 8564 1554 8570 1555
rect 8316 1540 8570 1554
rect 8316 1534 8319 1540
rect 8564 1538 8570 1540
rect 8587 1538 8593 1555
rect 8564 1535 8593 1538
rect 8609 1534 8612 1560
rect 8638 1554 8641 1560
rect 8978 1555 9007 1558
rect 8978 1554 8984 1555
rect 8638 1540 8984 1554
rect 8638 1534 8641 1540
rect 8978 1538 8984 1540
rect 9001 1538 9007 1555
rect 8978 1535 9007 1538
rect 9161 1534 9164 1560
rect 9190 1554 9193 1560
rect 9530 1555 9559 1558
rect 9530 1554 9536 1555
rect 9190 1540 9536 1554
rect 9190 1534 9193 1540
rect 9530 1538 9536 1540
rect 9553 1538 9559 1555
rect 9530 1535 9559 1538
rect 9575 1534 9578 1560
rect 9604 1554 9607 1560
rect 9990 1555 10019 1558
rect 9990 1554 9996 1555
rect 9604 1540 9996 1554
rect 9604 1534 9607 1540
rect 9990 1538 9996 1540
rect 10013 1538 10019 1555
rect 9990 1535 10019 1538
rect 10081 1534 10084 1560
rect 10110 1554 10113 1560
rect 10542 1555 10571 1558
rect 10542 1554 10548 1555
rect 10110 1540 10548 1554
rect 10110 1534 10113 1540
rect 10542 1538 10548 1540
rect 10565 1538 10571 1555
rect 10542 1535 10571 1538
rect 10633 1534 10636 1560
rect 10662 1554 10665 1560
rect 11140 1555 11169 1558
rect 11140 1554 11146 1555
rect 10662 1540 11146 1554
rect 10662 1534 10665 1540
rect 11140 1538 11146 1540
rect 11163 1538 11169 1555
rect 11140 1535 11169 1538
rect 11185 1534 11188 1560
rect 11214 1554 11217 1560
rect 11692 1555 11721 1558
rect 11692 1554 11698 1555
rect 11214 1540 11698 1554
rect 11214 1534 11217 1540
rect 11692 1538 11698 1540
rect 11715 1538 11721 1555
rect 11692 1535 11721 1538
rect 11737 1534 11740 1560
rect 11766 1554 11769 1560
rect 12106 1555 12135 1558
rect 12106 1554 12112 1555
rect 11766 1540 12112 1554
rect 11766 1534 11769 1540
rect 12106 1538 12112 1540
rect 12129 1538 12135 1555
rect 12106 1535 12135 1538
rect 12151 1534 12154 1560
rect 12180 1554 12183 1560
rect 12704 1555 12733 1558
rect 12704 1554 12710 1555
rect 12180 1540 12710 1554
rect 12180 1534 12183 1540
rect 12704 1538 12710 1540
rect 12727 1538 12733 1555
rect 12704 1535 12733 1538
rect 12979 1534 12982 1560
rect 13008 1554 13011 1560
rect 13578 1555 13607 1558
rect 13578 1554 13584 1555
rect 13008 1540 13584 1554
rect 13008 1534 13011 1540
rect 13578 1538 13584 1540
rect 13601 1538 13607 1555
rect 13578 1535 13607 1538
rect 13623 1534 13626 1560
rect 13652 1554 13655 1560
rect 14130 1555 14159 1558
rect 14130 1554 14136 1555
rect 13652 1540 14136 1554
rect 13652 1534 13655 1540
rect 14130 1538 14136 1540
rect 14153 1538 14159 1555
rect 14130 1535 14159 1538
rect 14497 1534 14500 1560
rect 14526 1554 14529 1560
rect 15004 1555 15033 1558
rect 15004 1554 15010 1555
rect 14526 1540 15010 1554
rect 14526 1534 14529 1540
rect 15004 1538 15010 1540
rect 15027 1538 15033 1555
rect 15004 1535 15033 1538
rect 15049 1534 15052 1560
rect 15078 1554 15081 1560
rect 15556 1555 15585 1558
rect 15556 1554 15562 1555
rect 15078 1540 15562 1554
rect 15078 1534 15081 1540
rect 15556 1538 15562 1540
rect 15579 1538 15585 1555
rect 15556 1535 15585 1538
rect 15877 1534 15880 1560
rect 15906 1554 15909 1560
rect 16154 1555 16183 1558
rect 16154 1554 16160 1555
rect 15906 1540 16160 1554
rect 15906 1534 15909 1540
rect 16154 1538 16160 1540
rect 16177 1538 16183 1555
rect 16154 1535 16183 1538
rect 16199 1534 16202 1560
rect 16228 1554 16231 1560
rect 16706 1555 16735 1558
rect 16706 1554 16712 1555
rect 16228 1540 16712 1554
rect 16228 1534 16231 1540
rect 16706 1538 16712 1540
rect 16729 1538 16735 1555
rect 16706 1535 16735 1538
rect 16751 1534 16754 1560
rect 16780 1554 16783 1560
rect 17258 1555 17287 1558
rect 17258 1554 17264 1555
rect 16780 1540 17264 1554
rect 16780 1534 16783 1540
rect 17258 1538 17264 1540
rect 17281 1538 17287 1555
rect 17258 1535 17287 1538
rect 17395 1534 17398 1560
rect 17424 1554 17427 1560
rect 17994 1555 18023 1558
rect 17994 1554 18000 1555
rect 17424 1540 18000 1554
rect 17424 1534 17427 1540
rect 17994 1538 18000 1540
rect 18017 1538 18023 1555
rect 17994 1535 18023 1538
rect 18223 1534 18226 1560
rect 18252 1554 18255 1560
rect 18730 1555 18759 1558
rect 18730 1554 18736 1555
rect 18252 1540 18736 1554
rect 18252 1534 18255 1540
rect 18730 1538 18736 1540
rect 18753 1538 18759 1555
rect 18730 1535 18759 1538
rect 18775 1534 18778 1560
rect 18804 1554 18807 1560
rect 19282 1555 19311 1558
rect 19282 1554 19288 1555
rect 18804 1540 19288 1554
rect 18804 1534 18807 1540
rect 19282 1538 19288 1540
rect 19305 1538 19311 1555
rect 19282 1535 19311 1538
rect 19327 1534 19330 1560
rect 19356 1554 19359 1560
rect 19834 1555 19863 1558
rect 19834 1554 19840 1555
rect 19356 1540 19840 1554
rect 19356 1534 19359 1540
rect 19834 1538 19840 1540
rect 19857 1538 19863 1555
rect 19834 1535 19863 1538
rect 19879 1534 19882 1560
rect 19908 1554 19911 1560
rect 20432 1555 20461 1558
rect 20432 1554 20438 1555
rect 19908 1540 20438 1554
rect 19908 1534 19911 1540
rect 20432 1538 20438 1540
rect 20455 1538 20461 1555
rect 20432 1535 20461 1538
rect 4700 1521 4729 1524
rect 4700 1520 4706 1521
rect 4590 1506 4706 1520
rect 4590 1500 4593 1506
rect 4700 1504 4706 1506
rect 4723 1504 4729 1521
rect 4700 1501 4729 1504
rect 5252 1521 5281 1524
rect 5252 1504 5258 1521
rect 5275 1504 5281 1521
rect 5527 1520 5530 1526
rect 5507 1506 5530 1520
rect 5252 1501 5281 1504
rect 5527 1500 5530 1506
rect 5556 1500 5559 1526
rect 5665 1500 5668 1526
rect 5694 1520 5697 1526
rect 5850 1521 5879 1524
rect 5850 1520 5856 1521
rect 5694 1506 5856 1520
rect 5694 1500 5697 1506
rect 5850 1504 5856 1506
rect 5873 1504 5879 1521
rect 6217 1520 6220 1526
rect 6197 1506 6220 1520
rect 5850 1501 5879 1504
rect 6217 1500 6220 1506
rect 6246 1500 6249 1526
rect 6355 1500 6358 1526
rect 6384 1520 6387 1526
rect 6494 1521 6523 1524
rect 6494 1520 6500 1521
rect 6384 1506 6500 1520
rect 6384 1500 6387 1506
rect 6494 1504 6500 1506
rect 6517 1504 6523 1521
rect 6494 1501 6523 1504
rect 7183 1500 7186 1526
rect 7212 1520 7215 1526
rect 7460 1521 7489 1524
rect 7460 1520 7466 1521
rect 7212 1506 7466 1520
rect 7212 1500 7215 1506
rect 7460 1504 7466 1506
rect 7483 1504 7489 1521
rect 7460 1501 7489 1504
rect 7597 1500 7600 1526
rect 7626 1520 7629 1526
rect 7736 1521 7765 1524
rect 7736 1520 7742 1521
rect 7626 1506 7742 1520
rect 7626 1500 7629 1506
rect 7736 1504 7742 1506
rect 7759 1504 7765 1521
rect 7736 1501 7765 1504
rect 7781 1500 7784 1526
rect 7810 1520 7813 1526
rect 8012 1521 8041 1524
rect 8012 1520 8018 1521
rect 7810 1506 8018 1520
rect 7810 1500 7813 1506
rect 8012 1504 8018 1506
rect 8035 1504 8041 1521
rect 8012 1501 8041 1504
rect 8333 1500 8336 1526
rect 8362 1520 8365 1526
rect 8702 1521 8731 1524
rect 8702 1520 8708 1521
rect 8362 1506 8708 1520
rect 8362 1500 8365 1506
rect 8702 1504 8708 1506
rect 8725 1504 8731 1521
rect 8702 1501 8731 1504
rect 8747 1500 8750 1526
rect 8776 1520 8779 1526
rect 9116 1521 9145 1524
rect 9116 1520 9122 1521
rect 8776 1506 9122 1520
rect 8776 1500 8779 1506
rect 9116 1504 9122 1506
rect 9139 1504 9145 1521
rect 9116 1501 9145 1504
rect 9437 1500 9440 1526
rect 9466 1520 9469 1526
rect 9852 1521 9881 1524
rect 9852 1520 9858 1521
rect 9466 1506 9858 1520
rect 9466 1500 9469 1506
rect 9852 1504 9858 1506
rect 9875 1504 9881 1521
rect 9852 1501 9881 1504
rect 9943 1500 9946 1526
rect 9972 1520 9975 1526
rect 10404 1521 10433 1524
rect 10404 1520 10410 1521
rect 9972 1506 10410 1520
rect 9972 1500 9975 1506
rect 10404 1504 10410 1506
rect 10427 1504 10433 1521
rect 10404 1501 10433 1504
rect 10495 1500 10498 1526
rect 10524 1520 10527 1526
rect 11002 1521 11031 1524
rect 11002 1520 11008 1521
rect 10524 1506 11008 1520
rect 10524 1500 10527 1506
rect 11002 1504 11008 1506
rect 11025 1504 11031 1521
rect 11002 1501 11031 1504
rect 11047 1500 11050 1526
rect 11076 1520 11079 1526
rect 11416 1521 11445 1524
rect 11416 1520 11422 1521
rect 11076 1506 11422 1520
rect 11076 1500 11079 1506
rect 11416 1504 11422 1506
rect 11439 1504 11445 1521
rect 11416 1501 11445 1504
rect 11461 1500 11464 1526
rect 11490 1520 11493 1526
rect 11968 1521 11997 1524
rect 11968 1520 11974 1521
rect 11490 1506 11974 1520
rect 11490 1500 11493 1506
rect 11968 1504 11974 1506
rect 11991 1504 11997 1521
rect 11968 1501 11997 1504
rect 12013 1500 12016 1526
rect 12042 1520 12045 1526
rect 12566 1521 12595 1524
rect 12566 1520 12572 1521
rect 12042 1506 12572 1520
rect 12042 1500 12045 1506
rect 12566 1504 12572 1506
rect 12589 1504 12595 1521
rect 12566 1501 12595 1504
rect 12749 1500 12752 1526
rect 12778 1520 12781 1526
rect 13256 1521 13285 1524
rect 13256 1520 13262 1521
rect 12778 1506 13262 1520
rect 12778 1500 12781 1506
rect 13256 1504 13262 1506
rect 13279 1504 13285 1521
rect 13256 1501 13285 1504
rect 13301 1500 13304 1526
rect 13330 1520 13333 1526
rect 13854 1521 13883 1524
rect 13854 1520 13860 1521
rect 13330 1506 13860 1520
rect 13330 1500 13333 1506
rect 13854 1504 13860 1506
rect 13877 1504 13883 1521
rect 13854 1501 13883 1504
rect 13899 1500 13902 1526
rect 13928 1520 13931 1526
rect 14406 1521 14435 1524
rect 14406 1520 14412 1521
rect 13928 1506 14412 1520
rect 13928 1500 13931 1506
rect 14406 1504 14412 1506
rect 14429 1504 14435 1521
rect 14406 1501 14435 1504
rect 14635 1500 14638 1526
rect 14664 1520 14667 1526
rect 15142 1521 15171 1524
rect 15142 1520 15148 1521
rect 14664 1506 15148 1520
rect 14664 1500 14667 1506
rect 15142 1504 15148 1506
rect 15165 1504 15171 1521
rect 15142 1501 15171 1504
rect 15187 1500 15190 1526
rect 15216 1520 15219 1526
rect 15694 1521 15723 1524
rect 15694 1520 15700 1521
rect 15216 1506 15700 1520
rect 15216 1500 15219 1506
rect 15694 1504 15700 1506
rect 15717 1504 15723 1521
rect 15694 1501 15723 1504
rect 15923 1500 15926 1526
rect 15952 1520 15955 1526
rect 16292 1521 16321 1524
rect 16292 1520 16298 1521
rect 15952 1506 16298 1520
rect 15952 1500 15955 1506
rect 16292 1504 16298 1506
rect 16315 1504 16321 1521
rect 16292 1501 16321 1504
rect 16337 1500 16340 1526
rect 16366 1520 16369 1526
rect 16844 1521 16873 1524
rect 16844 1520 16850 1521
rect 16366 1506 16850 1520
rect 16366 1500 16369 1506
rect 16844 1504 16850 1506
rect 16867 1504 16873 1521
rect 16844 1501 16873 1504
rect 16889 1500 16892 1526
rect 16918 1520 16921 1526
rect 17442 1521 17471 1524
rect 17442 1520 17448 1521
rect 16918 1506 17448 1520
rect 16918 1500 16921 1506
rect 17442 1504 17448 1506
rect 17465 1504 17471 1521
rect 17442 1501 17471 1504
rect 17533 1500 17536 1526
rect 17562 1520 17565 1526
rect 18132 1521 18161 1524
rect 18132 1520 18138 1521
rect 17562 1506 18138 1520
rect 17562 1500 17565 1506
rect 18132 1504 18138 1506
rect 18155 1504 18161 1521
rect 18408 1521 18437 1524
rect 18408 1520 18414 1521
rect 18132 1501 18161 1504
rect 18186 1506 18414 1520
rect 7 1466 10 1492
rect 36 1486 39 1492
rect 1802 1487 1831 1490
rect 1802 1486 1808 1487
rect 36 1472 1808 1486
rect 36 1466 39 1472
rect 1802 1470 1808 1472
rect 1825 1470 1831 1487
rect 2077 1486 2080 1492
rect 2057 1472 2080 1486
rect 1802 1467 1831 1470
rect 2077 1466 2080 1472
rect 2106 1466 2109 1492
rect 2354 1487 2383 1490
rect 2354 1470 2360 1487
rect 2377 1470 2383 1487
rect 2354 1467 2383 1470
rect 283 1432 286 1458
rect 312 1452 315 1458
rect 2362 1452 2376 1467
rect 4975 1466 4978 1492
rect 5004 1486 5007 1492
rect 5114 1487 5143 1490
rect 5114 1486 5120 1487
rect 5004 1472 5120 1486
rect 5004 1466 5007 1472
rect 5114 1470 5120 1472
rect 5137 1470 5143 1487
rect 5114 1467 5143 1470
rect 6953 1466 6956 1492
rect 6982 1486 6985 1492
rect 7322 1487 7351 1490
rect 7322 1486 7328 1487
rect 6982 1472 7328 1486
rect 6982 1466 6985 1472
rect 7322 1470 7328 1472
rect 7345 1470 7351 1487
rect 7322 1467 7351 1470
rect 7873 1466 7876 1492
rect 7902 1486 7905 1492
rect 8150 1487 8179 1490
rect 8150 1486 8156 1487
rect 7902 1472 8156 1486
rect 7902 1466 7905 1472
rect 8150 1470 8156 1472
rect 8173 1470 8179 1487
rect 8150 1467 8179 1470
rect 8977 1466 8980 1492
rect 9006 1486 9009 1492
rect 9392 1487 9421 1490
rect 9392 1486 9398 1487
rect 9006 1472 9398 1486
rect 9006 1466 9009 1472
rect 9392 1470 9398 1472
rect 9415 1470 9421 1487
rect 9392 1467 9421 1470
rect 9805 1466 9808 1492
rect 9834 1486 9837 1492
rect 10266 1487 10295 1490
rect 10266 1486 10272 1487
rect 9834 1472 10272 1486
rect 9834 1466 9837 1472
rect 10266 1470 10272 1472
rect 10289 1470 10295 1487
rect 10266 1467 10295 1470
rect 10357 1466 10360 1492
rect 10386 1486 10389 1492
rect 10818 1487 10847 1490
rect 10818 1486 10824 1487
rect 10386 1472 10824 1486
rect 10386 1466 10389 1472
rect 10818 1470 10824 1472
rect 10841 1470 10847 1487
rect 10818 1467 10847 1470
rect 11093 1466 11096 1492
rect 11122 1486 11125 1492
rect 11554 1487 11583 1490
rect 11554 1486 11560 1487
rect 11122 1472 11560 1486
rect 11122 1466 11125 1472
rect 11554 1470 11560 1472
rect 11577 1470 11583 1487
rect 11554 1467 11583 1470
rect 11783 1466 11786 1492
rect 11812 1486 11815 1492
rect 12290 1487 12319 1490
rect 12290 1486 12296 1487
rect 11812 1472 12296 1486
rect 11812 1466 11815 1472
rect 12290 1470 12296 1472
rect 12313 1470 12319 1487
rect 12290 1467 12319 1470
rect 12427 1466 12430 1492
rect 12456 1486 12459 1492
rect 12842 1487 12871 1490
rect 12842 1486 12848 1487
rect 12456 1472 12848 1486
rect 12456 1466 12459 1472
rect 12842 1470 12848 1472
rect 12865 1470 12871 1487
rect 12842 1467 12871 1470
rect 12933 1466 12936 1492
rect 12962 1486 12965 1492
rect 12980 1487 13009 1490
rect 12980 1486 12986 1487
rect 12962 1472 12986 1486
rect 12962 1466 12965 1472
rect 12980 1470 12986 1472
rect 13003 1470 13009 1487
rect 13394 1487 13423 1490
rect 13394 1486 13400 1487
rect 12980 1467 13009 1470
rect 13103 1472 13400 1486
rect 312 1438 2376 1452
rect 312 1432 315 1438
rect 12887 1432 12890 1458
rect 12916 1452 12919 1458
rect 13103 1452 13117 1472
rect 13394 1470 13400 1472
rect 13417 1470 13423 1487
rect 13394 1467 13423 1470
rect 13439 1466 13442 1492
rect 13468 1486 13471 1492
rect 13992 1487 14021 1490
rect 13992 1486 13998 1487
rect 13468 1472 13998 1486
rect 13468 1466 13471 1472
rect 13992 1470 13998 1472
rect 14015 1470 14021 1487
rect 13992 1467 14021 1470
rect 14037 1466 14040 1492
rect 14066 1486 14069 1492
rect 14544 1487 14573 1490
rect 14544 1486 14550 1487
rect 14066 1472 14550 1486
rect 14066 1466 14069 1472
rect 14544 1470 14550 1472
rect 14567 1470 14573 1487
rect 14544 1467 14573 1470
rect 14682 1487 14711 1490
rect 14682 1470 14688 1487
rect 14705 1470 14711 1487
rect 14682 1467 14711 1470
rect 12916 1438 13117 1452
rect 12916 1432 12919 1438
rect 14083 1432 14086 1458
rect 14112 1452 14115 1458
rect 14690 1452 14704 1467
rect 14773 1466 14776 1492
rect 14802 1486 14805 1492
rect 15280 1487 15309 1490
rect 15280 1486 15286 1487
rect 14802 1472 15286 1486
rect 14802 1466 14805 1472
rect 15280 1470 15286 1472
rect 15303 1470 15309 1487
rect 15280 1467 15309 1470
rect 15325 1466 15328 1492
rect 15354 1486 15357 1492
rect 15832 1487 15861 1490
rect 15832 1486 15838 1487
rect 15354 1472 15838 1486
rect 15354 1466 15357 1472
rect 15832 1470 15838 1472
rect 15855 1470 15861 1487
rect 15832 1467 15861 1470
rect 16061 1466 16064 1492
rect 16090 1486 16093 1492
rect 16568 1487 16597 1490
rect 16568 1486 16574 1487
rect 16090 1472 16574 1486
rect 16090 1466 16093 1472
rect 16568 1470 16574 1472
rect 16591 1470 16597 1487
rect 16568 1467 16597 1470
rect 16613 1466 16616 1492
rect 16642 1486 16645 1492
rect 17120 1487 17149 1490
rect 17120 1486 17126 1487
rect 16642 1472 17126 1486
rect 16642 1466 16645 1472
rect 17120 1470 17126 1472
rect 17143 1470 17149 1487
rect 17120 1467 17149 1470
rect 17257 1466 17260 1492
rect 17286 1486 17289 1492
rect 17718 1487 17747 1490
rect 17718 1486 17724 1487
rect 17286 1472 17724 1486
rect 17286 1466 17289 1472
rect 17718 1470 17724 1472
rect 17741 1470 17747 1487
rect 17718 1467 17747 1470
rect 17856 1487 17885 1490
rect 17856 1470 17862 1487
rect 17879 1470 17885 1487
rect 17856 1467 17885 1470
rect 14112 1438 14704 1452
rect 14112 1432 14115 1438
rect 17303 1432 17306 1458
rect 17332 1452 17335 1458
rect 17864 1452 17878 1467
rect 17947 1466 17950 1492
rect 17976 1486 17979 1492
rect 18186 1486 18200 1506
rect 18408 1504 18414 1506
rect 18431 1504 18437 1521
rect 18408 1501 18437 1504
rect 18499 1500 18502 1526
rect 18528 1520 18531 1526
rect 19006 1521 19035 1524
rect 19006 1520 19012 1521
rect 18528 1506 19012 1520
rect 18528 1500 18531 1506
rect 19006 1504 19012 1506
rect 19029 1504 19035 1521
rect 19006 1501 19035 1504
rect 19051 1500 19054 1526
rect 19080 1520 19083 1526
rect 19558 1521 19587 1524
rect 19558 1520 19564 1521
rect 19080 1506 19564 1520
rect 19080 1500 19083 1506
rect 19558 1504 19564 1506
rect 19581 1504 19587 1521
rect 19558 1501 19587 1504
rect 19603 1500 19606 1526
rect 19632 1520 19635 1526
rect 20156 1521 20185 1524
rect 20156 1520 20162 1521
rect 19632 1506 20162 1520
rect 19632 1500 19635 1506
rect 20156 1504 20162 1506
rect 20179 1504 20185 1521
rect 20156 1501 20185 1504
rect 20201 1500 20204 1526
rect 20230 1520 20233 1526
rect 20708 1521 20737 1524
rect 20708 1520 20714 1521
rect 20230 1506 20714 1520
rect 20230 1500 20233 1506
rect 20708 1504 20714 1506
rect 20731 1504 20737 1521
rect 20808 1520 20822 1574
rect 20845 1568 20848 1594
rect 20874 1588 20877 1594
rect 21306 1589 21335 1592
rect 21306 1588 21312 1589
rect 20874 1574 21312 1588
rect 20874 1568 20877 1574
rect 21306 1572 21312 1574
rect 21329 1572 21335 1589
rect 21306 1569 21335 1572
rect 21397 1568 21400 1594
rect 21426 1588 21429 1594
rect 21720 1589 21749 1592
rect 21720 1588 21726 1589
rect 21426 1574 21726 1588
rect 21426 1568 21429 1574
rect 21720 1572 21726 1574
rect 21743 1572 21749 1589
rect 21720 1569 21749 1572
rect 21765 1568 21768 1594
rect 21794 1588 21797 1594
rect 22134 1589 22163 1592
rect 22134 1588 22140 1589
rect 21794 1574 22140 1588
rect 21794 1568 21797 1574
rect 22134 1572 22140 1574
rect 22157 1572 22163 1589
rect 22134 1569 22163 1572
rect 22225 1568 22228 1594
rect 22254 1588 22257 1594
rect 22594 1589 22623 1592
rect 22594 1588 22600 1589
rect 22254 1574 22600 1588
rect 22254 1568 22257 1574
rect 22594 1572 22600 1574
rect 22617 1572 22623 1589
rect 22594 1569 22623 1572
rect 23743 1568 23746 1594
rect 23772 1588 23775 1594
rect 23882 1589 23911 1592
rect 23882 1588 23888 1589
rect 23772 1574 23888 1588
rect 23772 1568 23775 1574
rect 23882 1572 23888 1574
rect 23905 1572 23911 1589
rect 23882 1569 23911 1572
rect 24295 1568 24298 1594
rect 24324 1588 24327 1594
rect 24342 1589 24371 1592
rect 24342 1588 24348 1589
rect 24324 1574 24348 1588
rect 24324 1568 24327 1574
rect 24342 1572 24348 1574
rect 24365 1572 24371 1589
rect 24342 1569 24371 1572
rect 24433 1568 24436 1594
rect 24462 1588 24465 1594
rect 24480 1589 24509 1592
rect 24480 1588 24486 1589
rect 24462 1574 24486 1588
rect 24462 1568 24465 1574
rect 24480 1572 24486 1574
rect 24503 1572 24509 1589
rect 24480 1569 24509 1572
rect 24571 1568 24574 1594
rect 24600 1588 24603 1594
rect 24618 1589 24647 1592
rect 24618 1588 24624 1589
rect 24600 1574 24624 1588
rect 24600 1568 24603 1574
rect 24618 1572 24624 1574
rect 24641 1572 24647 1589
rect 24618 1569 24647 1572
rect 24709 1568 24712 1594
rect 24738 1588 24741 1594
rect 24756 1589 24785 1592
rect 24756 1588 24762 1589
rect 24738 1574 24762 1588
rect 24738 1568 24741 1574
rect 24756 1572 24762 1574
rect 24779 1572 24785 1589
rect 24756 1569 24785 1572
rect 24847 1568 24850 1594
rect 24876 1588 24879 1594
rect 24894 1589 24923 1592
rect 24894 1588 24900 1589
rect 24876 1574 24900 1588
rect 24876 1568 24879 1574
rect 24894 1572 24900 1574
rect 24917 1572 24923 1589
rect 24894 1569 24923 1572
rect 24985 1568 24988 1594
rect 25014 1588 25017 1594
rect 25170 1589 25199 1592
rect 25170 1588 25176 1589
rect 25014 1574 25176 1588
rect 25014 1568 25017 1574
rect 25170 1572 25176 1574
rect 25193 1572 25199 1589
rect 25170 1569 25199 1572
rect 25261 1568 25264 1594
rect 25290 1588 25293 1594
rect 25446 1589 25475 1592
rect 25446 1588 25452 1589
rect 25290 1574 25452 1588
rect 25290 1568 25293 1574
rect 25446 1572 25452 1574
rect 25469 1572 25475 1589
rect 25446 1569 25475 1572
rect 25537 1568 25540 1594
rect 25566 1588 25569 1594
rect 25584 1589 25613 1592
rect 25584 1588 25590 1589
rect 25566 1574 25590 1588
rect 25566 1568 25569 1574
rect 25584 1572 25590 1574
rect 25607 1572 25613 1589
rect 25584 1569 25613 1572
rect 25675 1568 25678 1594
rect 25704 1588 25707 1594
rect 25860 1589 25889 1592
rect 25860 1588 25866 1589
rect 25704 1574 25866 1588
rect 25704 1568 25707 1574
rect 25860 1572 25866 1574
rect 25883 1572 25889 1589
rect 25860 1569 25889 1572
rect 25951 1568 25954 1594
rect 25980 1588 25983 1594
rect 26136 1589 26165 1592
rect 26136 1588 26142 1589
rect 25980 1574 26142 1588
rect 25980 1568 25983 1574
rect 26136 1572 26142 1574
rect 26159 1572 26165 1589
rect 26136 1569 26165 1572
rect 26227 1568 26230 1594
rect 26256 1588 26259 1594
rect 26274 1589 26303 1592
rect 26274 1588 26280 1589
rect 26256 1574 26280 1588
rect 26256 1568 26259 1574
rect 26274 1572 26280 1574
rect 26297 1572 26303 1589
rect 26274 1569 26303 1572
rect 26365 1568 26368 1594
rect 26394 1588 26397 1594
rect 26596 1589 26625 1592
rect 26596 1588 26602 1589
rect 26394 1574 26602 1588
rect 26394 1568 26397 1574
rect 26596 1572 26602 1574
rect 26619 1572 26625 1589
rect 26596 1569 26625 1572
rect 26641 1568 26644 1594
rect 26670 1588 26673 1594
rect 26872 1589 26901 1592
rect 26872 1588 26878 1589
rect 26670 1574 26878 1588
rect 26670 1568 26673 1574
rect 26872 1572 26878 1574
rect 26895 1572 26901 1589
rect 26872 1569 26901 1572
rect 26917 1568 26920 1594
rect 26946 1588 26949 1594
rect 27010 1589 27039 1592
rect 27010 1588 27016 1589
rect 26946 1574 27016 1588
rect 26946 1568 26949 1574
rect 27010 1572 27016 1574
rect 27033 1572 27039 1589
rect 27010 1569 27039 1572
rect 27055 1568 27058 1594
rect 27084 1588 27087 1594
rect 27286 1589 27315 1592
rect 27286 1588 27292 1589
rect 27084 1574 27292 1588
rect 27084 1568 27087 1574
rect 27286 1572 27292 1574
rect 27309 1572 27315 1589
rect 27286 1569 27315 1572
rect 27331 1568 27334 1594
rect 27360 1588 27363 1594
rect 27562 1589 27591 1592
rect 27562 1588 27568 1589
rect 27360 1574 27568 1588
rect 27360 1568 27363 1574
rect 27562 1572 27568 1574
rect 27585 1572 27591 1589
rect 27562 1569 27591 1572
rect 27699 1568 27702 1594
rect 27728 1588 27731 1594
rect 27884 1589 27913 1592
rect 27884 1588 27890 1589
rect 27728 1574 27890 1588
rect 27728 1568 27731 1574
rect 27884 1572 27890 1574
rect 27907 1572 27913 1589
rect 27884 1569 27913 1572
rect 28021 1568 28024 1594
rect 28050 1588 28053 1594
rect 28298 1589 28327 1592
rect 28298 1588 28304 1589
rect 28050 1574 28304 1588
rect 28050 1568 28053 1574
rect 28298 1572 28304 1574
rect 28321 1572 28327 1589
rect 28298 1569 28327 1572
rect 28343 1568 28346 1594
rect 28372 1588 28375 1594
rect 28574 1589 28603 1592
rect 28574 1588 28580 1589
rect 28372 1574 28580 1588
rect 28372 1568 28375 1574
rect 28574 1572 28580 1574
rect 28597 1572 28603 1589
rect 28574 1569 28603 1572
rect 28757 1568 28760 1594
rect 28786 1588 28789 1594
rect 29034 1589 29063 1592
rect 29034 1588 29040 1589
rect 28786 1574 29040 1588
rect 28786 1568 28789 1574
rect 29034 1572 29040 1574
rect 29057 1572 29063 1589
rect 29034 1569 29063 1572
rect 29125 1568 29128 1594
rect 29154 1588 29157 1594
rect 29448 1589 29477 1592
rect 29448 1588 29454 1589
rect 29154 1574 29454 1588
rect 29154 1568 29157 1574
rect 29448 1572 29454 1574
rect 29471 1572 29477 1589
rect 29448 1569 29477 1572
rect 29539 1568 29542 1594
rect 29568 1588 29571 1594
rect 29862 1589 29891 1592
rect 29862 1588 29868 1589
rect 29568 1574 29868 1588
rect 29568 1568 29571 1574
rect 29862 1572 29868 1574
rect 29885 1572 29891 1589
rect 29862 1569 29891 1572
rect 29953 1568 29956 1594
rect 29982 1588 29985 1594
rect 30322 1589 30351 1592
rect 30322 1588 30328 1589
rect 29982 1574 30328 1588
rect 29982 1568 29985 1574
rect 30322 1572 30328 1574
rect 30345 1572 30351 1589
rect 30322 1569 30351 1572
rect 30367 1568 30370 1594
rect 30396 1588 30399 1594
rect 30598 1589 30627 1592
rect 30598 1588 30604 1589
rect 30396 1574 30604 1588
rect 30396 1568 30399 1574
rect 30598 1572 30604 1574
rect 30621 1572 30627 1589
rect 30598 1569 30627 1572
rect 30689 1568 30692 1594
rect 30718 1588 30721 1594
rect 31012 1589 31041 1592
rect 31012 1588 31018 1589
rect 30718 1574 31018 1588
rect 30718 1568 30721 1574
rect 31012 1572 31018 1574
rect 31035 1572 31041 1589
rect 31012 1569 31041 1572
rect 31057 1568 31060 1594
rect 31086 1588 31089 1594
rect 31288 1589 31317 1592
rect 31288 1588 31294 1589
rect 31086 1574 31294 1588
rect 31086 1568 31089 1574
rect 31288 1572 31294 1574
rect 31311 1572 31317 1589
rect 31288 1569 31317 1572
rect 31333 1568 31336 1594
rect 31362 1588 31365 1594
rect 31748 1589 31777 1592
rect 31748 1588 31754 1589
rect 31362 1574 31754 1588
rect 31362 1568 31365 1574
rect 31748 1572 31754 1574
rect 31771 1572 31777 1589
rect 31748 1569 31777 1572
rect 32161 1568 32164 1594
rect 32190 1588 32193 1594
rect 32576 1589 32605 1592
rect 32576 1588 32582 1589
rect 32190 1574 32582 1588
rect 32190 1568 32193 1574
rect 32576 1572 32582 1574
rect 32599 1572 32605 1589
rect 32576 1569 32605 1572
rect 32851 1568 32854 1594
rect 32880 1588 32883 1594
rect 33174 1589 33203 1592
rect 33174 1588 33180 1589
rect 32880 1574 33180 1588
rect 32880 1568 32883 1574
rect 33174 1572 33180 1574
rect 33197 1572 33203 1589
rect 33174 1569 33203 1572
rect 33265 1568 33268 1594
rect 33294 1588 33297 1594
rect 33312 1589 33341 1592
rect 33312 1588 33318 1589
rect 33294 1574 33318 1588
rect 33294 1568 33297 1574
rect 33312 1572 33318 1574
rect 33335 1572 33341 1589
rect 33541 1588 33544 1594
rect 33521 1574 33544 1588
rect 33312 1569 33341 1572
rect 33541 1568 33544 1574
rect 33570 1568 33573 1594
rect 33680 1589 33709 1592
rect 33680 1572 33686 1589
rect 33703 1588 33709 1589
rect 33725 1588 33728 1594
rect 33703 1574 33728 1588
rect 33703 1572 33709 1574
rect 33680 1569 33709 1572
rect 33725 1568 33728 1574
rect 33754 1568 33757 1594
rect 33817 1588 33820 1594
rect 33797 1574 33820 1588
rect 33817 1568 33820 1574
rect 33846 1568 33849 1594
rect 20983 1534 20986 1560
rect 21012 1554 21015 1560
rect 21444 1555 21473 1558
rect 21444 1554 21450 1555
rect 21012 1540 21450 1554
rect 21012 1534 21015 1540
rect 21444 1538 21450 1540
rect 21467 1538 21473 1555
rect 21444 1535 21473 1538
rect 21535 1534 21538 1560
rect 21564 1554 21567 1560
rect 21996 1555 22025 1558
rect 21996 1554 22002 1555
rect 21564 1540 22002 1554
rect 21564 1534 21567 1540
rect 21996 1538 22002 1540
rect 22019 1538 22025 1555
rect 21996 1535 22025 1538
rect 22363 1534 22366 1560
rect 22392 1554 22395 1560
rect 22732 1555 22761 1558
rect 22732 1554 22738 1555
rect 22392 1540 22738 1554
rect 22392 1534 22395 1540
rect 22732 1538 22738 1540
rect 22755 1538 22761 1555
rect 22732 1535 22761 1538
rect 25123 1534 25126 1560
rect 25152 1554 25155 1560
rect 25308 1555 25337 1558
rect 25308 1554 25314 1555
rect 25152 1540 25314 1554
rect 25152 1534 25155 1540
rect 25308 1538 25314 1540
rect 25331 1538 25337 1555
rect 25308 1535 25337 1538
rect 25813 1534 25816 1560
rect 25842 1554 25845 1560
rect 25998 1555 26027 1558
rect 25998 1554 26004 1555
rect 25842 1540 26004 1554
rect 25842 1534 25845 1540
rect 25998 1538 26004 1540
rect 26021 1538 26027 1555
rect 25998 1535 26027 1538
rect 26503 1534 26506 1560
rect 26532 1554 26535 1560
rect 26734 1555 26763 1558
rect 26734 1554 26740 1555
rect 26532 1540 26740 1554
rect 26532 1534 26535 1540
rect 26734 1538 26740 1540
rect 26757 1538 26763 1555
rect 26734 1535 26763 1538
rect 26963 1534 26966 1560
rect 26992 1554 26995 1560
rect 27148 1555 27177 1558
rect 27148 1554 27154 1555
rect 26992 1540 27154 1554
rect 26992 1534 26995 1540
rect 27148 1538 27154 1540
rect 27171 1538 27177 1555
rect 27148 1535 27177 1538
rect 27193 1534 27196 1560
rect 27222 1554 27225 1560
rect 27424 1555 27453 1558
rect 27424 1554 27430 1555
rect 27222 1540 27430 1554
rect 27222 1534 27225 1540
rect 27424 1538 27430 1540
rect 27447 1538 27453 1555
rect 27424 1535 27453 1538
rect 27469 1534 27472 1560
rect 27498 1554 27501 1560
rect 27746 1555 27775 1558
rect 27746 1554 27752 1555
rect 27498 1540 27752 1554
rect 27498 1534 27501 1540
rect 27746 1538 27752 1540
rect 27769 1538 27775 1555
rect 27746 1535 27775 1538
rect 28481 1534 28484 1560
rect 28510 1554 28513 1560
rect 28712 1555 28741 1558
rect 28712 1554 28718 1555
rect 28510 1540 28718 1554
rect 28510 1534 28513 1540
rect 28712 1538 28718 1540
rect 28735 1538 28741 1555
rect 28712 1535 28741 1538
rect 28987 1534 28990 1560
rect 29016 1554 29019 1560
rect 29172 1555 29201 1558
rect 29172 1554 29178 1555
rect 29016 1540 29178 1554
rect 29016 1534 29019 1540
rect 29172 1538 29178 1540
rect 29195 1538 29201 1555
rect 29172 1535 29201 1538
rect 29263 1534 29266 1560
rect 29292 1554 29295 1560
rect 29586 1555 29615 1558
rect 29586 1554 29592 1555
rect 29292 1540 29592 1554
rect 29292 1534 29295 1540
rect 29586 1538 29592 1540
rect 29609 1538 29615 1555
rect 29586 1535 29615 1538
rect 29677 1534 29680 1560
rect 29706 1554 29709 1560
rect 30000 1555 30029 1558
rect 30000 1554 30006 1555
rect 29706 1540 30006 1554
rect 29706 1534 29709 1540
rect 30000 1538 30006 1540
rect 30023 1538 30029 1555
rect 30000 1535 30029 1538
rect 30091 1534 30094 1560
rect 30120 1554 30123 1560
rect 30460 1555 30489 1558
rect 30460 1554 30466 1555
rect 30120 1540 30466 1554
rect 30120 1534 30123 1540
rect 30460 1538 30466 1540
rect 30483 1538 30489 1555
rect 30460 1535 30489 1538
rect 30505 1534 30508 1560
rect 30534 1554 30537 1560
rect 30874 1555 30903 1558
rect 30874 1554 30880 1555
rect 30534 1540 30880 1554
rect 30534 1534 30537 1540
rect 30874 1538 30880 1540
rect 30897 1538 30903 1555
rect 30874 1535 30903 1538
rect 31103 1534 31106 1560
rect 31132 1554 31135 1560
rect 31426 1555 31455 1558
rect 31426 1554 31432 1555
rect 31132 1540 31432 1554
rect 31132 1534 31135 1540
rect 31426 1538 31432 1540
rect 31449 1538 31455 1555
rect 31426 1535 31455 1538
rect 31471 1534 31474 1560
rect 31500 1554 31503 1560
rect 31886 1555 31915 1558
rect 31886 1554 31892 1555
rect 31500 1540 31892 1554
rect 31500 1534 31503 1540
rect 31886 1538 31892 1540
rect 31909 1538 31915 1555
rect 31886 1535 31915 1538
rect 32023 1534 32026 1560
rect 32052 1554 32055 1560
rect 32438 1555 32467 1558
rect 32438 1554 32444 1555
rect 32052 1540 32444 1554
rect 32052 1534 32055 1540
rect 32438 1538 32444 1540
rect 32461 1538 32467 1555
rect 32438 1535 32467 1538
rect 32621 1534 32624 1560
rect 32650 1554 32653 1560
rect 33036 1555 33065 1558
rect 33036 1554 33042 1555
rect 32650 1540 33042 1554
rect 32650 1534 32653 1540
rect 33036 1538 33042 1540
rect 33059 1538 33065 1555
rect 33036 1535 33065 1538
rect 21122 1521 21151 1524
rect 21122 1520 21128 1521
rect 20808 1506 21128 1520
rect 20708 1501 20737 1504
rect 21122 1504 21128 1506
rect 21145 1504 21151 1521
rect 21122 1501 21151 1504
rect 21167 1500 21170 1526
rect 21196 1520 21199 1526
rect 21582 1521 21611 1524
rect 21582 1520 21588 1521
rect 21196 1506 21588 1520
rect 21196 1500 21199 1506
rect 21582 1504 21588 1506
rect 21605 1504 21611 1521
rect 21582 1501 21611 1504
rect 21811 1500 21814 1526
rect 21840 1520 21843 1526
rect 22272 1521 22301 1524
rect 22272 1520 22278 1521
rect 21840 1506 22278 1520
rect 21840 1500 21843 1506
rect 22272 1504 22278 1506
rect 22295 1504 22301 1521
rect 22272 1501 22301 1504
rect 22501 1500 22504 1526
rect 22530 1520 22533 1526
rect 22870 1521 22899 1524
rect 22870 1520 22876 1521
rect 22530 1506 22876 1520
rect 22530 1500 22533 1506
rect 22870 1504 22876 1506
rect 22893 1504 22899 1521
rect 22870 1501 22899 1504
rect 23881 1500 23884 1526
rect 23910 1520 23913 1526
rect 24020 1521 24049 1524
rect 24020 1520 24026 1521
rect 23910 1506 24026 1520
rect 23910 1500 23913 1506
rect 24020 1504 24026 1506
rect 24043 1504 24049 1521
rect 24020 1501 24049 1504
rect 25583 1500 25586 1526
rect 25612 1520 25615 1526
rect 25722 1521 25751 1524
rect 25722 1520 25728 1521
rect 25612 1506 25728 1520
rect 25612 1500 25615 1506
rect 25722 1504 25728 1506
rect 25745 1504 25751 1521
rect 25722 1501 25751 1504
rect 26273 1500 26276 1526
rect 26302 1520 26305 1526
rect 26458 1521 26487 1524
rect 26458 1520 26464 1521
rect 26302 1506 26464 1520
rect 26302 1500 26305 1506
rect 26458 1504 26464 1506
rect 26481 1504 26487 1521
rect 26458 1501 26487 1504
rect 27883 1500 27886 1526
rect 27912 1520 27915 1526
rect 28160 1521 28189 1524
rect 28160 1520 28166 1521
rect 27912 1506 28166 1520
rect 27912 1500 27915 1506
rect 28160 1504 28166 1506
rect 28183 1504 28189 1521
rect 28160 1501 28189 1504
rect 28297 1500 28300 1526
rect 28326 1520 28329 1526
rect 28436 1521 28465 1524
rect 28436 1520 28442 1521
rect 28326 1506 28442 1520
rect 28326 1500 28329 1506
rect 28436 1504 28442 1506
rect 28459 1504 28465 1521
rect 28436 1501 28465 1504
rect 28573 1500 28576 1526
rect 28602 1520 28605 1526
rect 28850 1521 28879 1524
rect 28850 1520 28856 1521
rect 28602 1506 28856 1520
rect 28602 1500 28605 1506
rect 28850 1504 28856 1506
rect 28873 1504 28879 1521
rect 28850 1501 28879 1504
rect 29033 1500 29036 1526
rect 29062 1520 29065 1526
rect 29310 1521 29339 1524
rect 29310 1520 29316 1521
rect 29062 1506 29316 1520
rect 29062 1500 29065 1506
rect 29310 1504 29316 1506
rect 29333 1504 29339 1521
rect 29310 1501 29339 1504
rect 29401 1500 29404 1526
rect 29430 1520 29433 1526
rect 29724 1521 29753 1524
rect 29724 1520 29730 1521
rect 29430 1506 29730 1520
rect 29430 1500 29433 1506
rect 29724 1504 29730 1506
rect 29747 1504 29753 1521
rect 29724 1501 29753 1504
rect 29815 1500 29818 1526
rect 29844 1520 29847 1526
rect 30138 1521 30167 1524
rect 30138 1520 30144 1521
rect 29844 1506 30144 1520
rect 29844 1500 29847 1506
rect 30138 1504 30144 1506
rect 30161 1504 30167 1521
rect 30138 1501 30167 1504
rect 30413 1500 30416 1526
rect 30442 1520 30445 1526
rect 30736 1521 30765 1524
rect 30736 1520 30742 1521
rect 30442 1506 30742 1520
rect 30442 1500 30445 1506
rect 30736 1504 30742 1506
rect 30759 1504 30765 1521
rect 30736 1501 30765 1504
rect 30781 1500 30784 1526
rect 30810 1520 30813 1526
rect 31150 1521 31179 1524
rect 31150 1520 31156 1521
rect 30810 1506 31156 1520
rect 30810 1500 30813 1506
rect 31150 1504 31156 1506
rect 31173 1504 31179 1521
rect 31150 1501 31179 1504
rect 31195 1500 31198 1526
rect 31224 1520 31227 1526
rect 31610 1521 31639 1524
rect 31610 1520 31616 1521
rect 31224 1506 31616 1520
rect 31224 1500 31227 1506
rect 31610 1504 31616 1506
rect 31633 1504 31639 1521
rect 31610 1501 31639 1504
rect 31793 1500 31796 1526
rect 31822 1520 31825 1526
rect 32162 1521 32191 1524
rect 32162 1520 32168 1521
rect 31822 1506 32168 1520
rect 31822 1500 31825 1506
rect 32162 1504 32168 1506
rect 32185 1504 32191 1521
rect 32162 1501 32191 1504
rect 32345 1500 32348 1526
rect 32374 1520 32377 1526
rect 32714 1521 32743 1524
rect 32714 1520 32720 1521
rect 32374 1506 32720 1520
rect 32374 1500 32377 1506
rect 32714 1504 32720 1506
rect 32737 1504 32743 1521
rect 32714 1501 32743 1504
rect 32990 1521 33019 1524
rect 32990 1504 32996 1521
rect 33013 1520 33019 1521
rect 33955 1520 33958 1526
rect 33013 1506 33958 1520
rect 33013 1504 33019 1506
rect 32990 1501 33019 1504
rect 33955 1500 33958 1506
rect 33984 1500 33987 1526
rect 17976 1472 18200 1486
rect 18546 1487 18575 1490
rect 17976 1466 17979 1472
rect 18546 1470 18552 1487
rect 18569 1470 18575 1487
rect 18546 1467 18575 1470
rect 17332 1438 17878 1452
rect 17332 1432 17335 1438
rect 17993 1432 17996 1458
rect 18022 1452 18025 1458
rect 18554 1452 18568 1467
rect 18683 1466 18686 1492
rect 18712 1486 18715 1492
rect 19144 1487 19173 1490
rect 19144 1486 19150 1487
rect 18712 1472 19150 1486
rect 18712 1466 18715 1472
rect 19144 1470 19150 1472
rect 19167 1470 19173 1487
rect 19144 1467 19173 1470
rect 19189 1466 19192 1492
rect 19218 1486 19221 1492
rect 19696 1487 19725 1490
rect 19696 1486 19702 1487
rect 19218 1472 19702 1486
rect 19218 1466 19221 1472
rect 19696 1470 19702 1472
rect 19719 1470 19725 1487
rect 19696 1467 19725 1470
rect 19741 1466 19744 1492
rect 19770 1486 19773 1492
rect 20294 1487 20323 1490
rect 20294 1486 20300 1487
rect 19770 1472 20300 1486
rect 19770 1466 19773 1472
rect 20294 1470 20300 1472
rect 20317 1470 20323 1487
rect 20294 1467 20323 1470
rect 20339 1466 20342 1492
rect 20368 1486 20371 1492
rect 20846 1487 20875 1490
rect 20846 1486 20852 1487
rect 20368 1472 20852 1486
rect 20368 1466 20371 1472
rect 20846 1470 20852 1472
rect 20869 1470 20875 1487
rect 20846 1467 20875 1470
rect 20984 1487 21013 1490
rect 20984 1470 20990 1487
rect 21007 1470 21013 1487
rect 20984 1467 21013 1470
rect 18022 1438 18568 1452
rect 18022 1432 18025 1438
rect 20431 1432 20434 1458
rect 20460 1452 20463 1458
rect 20992 1452 21006 1467
rect 21443 1466 21446 1492
rect 21472 1486 21475 1492
rect 21858 1487 21887 1490
rect 21858 1486 21864 1487
rect 21472 1472 21864 1486
rect 21472 1466 21475 1472
rect 21858 1470 21864 1472
rect 21881 1470 21887 1487
rect 21858 1467 21887 1470
rect 21949 1466 21952 1492
rect 21978 1486 21981 1492
rect 22410 1487 22439 1490
rect 22410 1486 22416 1487
rect 21978 1472 22416 1486
rect 21978 1466 21981 1472
rect 22410 1470 22416 1472
rect 22433 1470 22439 1487
rect 22410 1467 22439 1470
rect 27745 1466 27748 1492
rect 27774 1486 27777 1492
rect 28022 1487 28051 1490
rect 28022 1486 28028 1487
rect 27774 1472 28028 1486
rect 27774 1466 27777 1472
rect 28022 1470 28028 1472
rect 28045 1470 28051 1487
rect 28022 1467 28051 1470
rect 31747 1466 31750 1492
rect 31776 1486 31779 1492
rect 32024 1487 32053 1490
rect 32024 1486 32030 1487
rect 31776 1472 32030 1486
rect 31776 1466 31779 1472
rect 32024 1470 32030 1472
rect 32047 1470 32053 1487
rect 32024 1467 32053 1470
rect 32300 1487 32329 1490
rect 32300 1470 32306 1487
rect 32323 1470 32329 1487
rect 32300 1467 32329 1470
rect 20460 1438 21006 1452
rect 20460 1432 20463 1438
rect 31885 1432 31888 1458
rect 31914 1452 31917 1458
rect 32308 1452 32322 1467
rect 31914 1438 32322 1452
rect 31914 1432 31917 1438
rect 467 1398 470 1424
rect 496 1418 499 1424
rect 2813 1418 2816 1424
rect 496 1404 2816 1418
rect 496 1398 499 1404
rect 2813 1398 2816 1404
rect 2842 1398 2845 1424
rect 644 1373 34408 1384
rect 644 1347 3631 1373
rect 3657 1347 9631 1373
rect 9657 1347 15631 1373
rect 15657 1347 21631 1373
rect 21657 1347 27631 1373
rect 27657 1347 33631 1373
rect 33657 1347 34408 1373
rect 644 1336 34408 1347
rect 1479 1262 1482 1288
rect 1508 1282 1511 1288
rect 1508 1268 2100 1282
rect 1508 1262 1511 1268
rect 973 1228 976 1254
rect 1002 1248 1005 1254
rect 1388 1249 1417 1252
rect 1388 1248 1394 1249
rect 1002 1234 1394 1248
rect 1002 1228 1005 1234
rect 1388 1232 1394 1234
rect 1411 1232 1417 1249
rect 1388 1229 1417 1232
rect 1756 1249 1785 1252
rect 1756 1232 1762 1249
rect 1779 1248 1785 1249
rect 1939 1248 1942 1254
rect 1779 1234 1942 1248
rect 1779 1232 1785 1234
rect 1756 1229 1785 1232
rect 1939 1228 1942 1234
rect 1968 1228 1971 1254
rect 2086 1252 2100 1268
rect 2078 1249 2107 1252
rect 2078 1232 2084 1249
rect 2101 1232 2107 1249
rect 2078 1229 2107 1232
rect 2215 1228 2218 1254
rect 2244 1248 2247 1254
rect 2630 1249 2659 1252
rect 2630 1248 2636 1249
rect 2244 1234 2636 1248
rect 2244 1228 2247 1234
rect 2630 1232 2636 1234
rect 2653 1232 2659 1249
rect 2630 1229 2659 1232
rect 3043 1228 3046 1254
rect 3072 1248 3075 1254
rect 3136 1249 3165 1252
rect 3136 1248 3142 1249
rect 3072 1234 3142 1248
rect 3072 1228 3075 1234
rect 3136 1232 3142 1234
rect 3159 1232 3165 1249
rect 3136 1229 3165 1232
rect 5803 1228 5806 1254
rect 5832 1248 5835 1254
rect 5942 1249 5971 1252
rect 5942 1248 5948 1249
rect 5832 1234 5948 1248
rect 5832 1228 5835 1234
rect 5942 1232 5948 1234
rect 5965 1232 5971 1249
rect 5942 1229 5971 1232
rect 14221 1228 14224 1254
rect 14250 1248 14253 1254
rect 14406 1249 14435 1252
rect 14406 1248 14412 1249
rect 14250 1234 14412 1248
rect 14250 1228 14253 1234
rect 14406 1232 14412 1234
rect 14429 1232 14435 1249
rect 14406 1229 14435 1232
rect 18085 1228 18088 1254
rect 18114 1248 18117 1254
rect 18270 1249 18299 1252
rect 18270 1248 18276 1249
rect 18114 1234 18276 1248
rect 18114 1228 18117 1234
rect 18270 1232 18276 1234
rect 18293 1232 18299 1249
rect 18270 1229 18299 1232
rect 20707 1228 20710 1254
rect 20736 1248 20739 1254
rect 20846 1249 20875 1252
rect 20846 1248 20852 1249
rect 20736 1234 20852 1248
rect 20736 1228 20739 1234
rect 20846 1232 20852 1234
rect 20869 1232 20875 1249
rect 20846 1229 20875 1232
rect 22087 1228 22090 1254
rect 22116 1248 22119 1254
rect 22134 1249 22163 1252
rect 22134 1248 22140 1249
rect 22116 1234 22140 1248
rect 22116 1228 22119 1234
rect 22134 1232 22140 1234
rect 22157 1232 22163 1249
rect 22639 1248 22642 1254
rect 22619 1234 22642 1248
rect 22134 1229 22163 1232
rect 22639 1228 22642 1234
rect 22668 1228 22671 1254
rect 22777 1228 22780 1254
rect 22806 1248 22809 1254
rect 22915 1248 22918 1254
rect 22806 1234 22828 1248
rect 22895 1234 22918 1248
rect 22806 1228 22809 1234
rect 22915 1228 22918 1234
rect 22944 1228 22947 1254
rect 23053 1248 23056 1254
rect 23033 1234 23056 1248
rect 23053 1228 23056 1234
rect 23082 1228 23085 1254
rect 23191 1248 23194 1254
rect 23171 1234 23194 1248
rect 23191 1228 23194 1234
rect 23220 1228 23223 1254
rect 23329 1248 23332 1254
rect 23309 1234 23332 1248
rect 23329 1228 23332 1234
rect 23358 1228 23361 1254
rect 23467 1248 23470 1254
rect 23447 1234 23470 1248
rect 23467 1228 23470 1234
rect 23496 1228 23499 1254
rect 23605 1248 23608 1254
rect 23585 1234 23608 1248
rect 23605 1228 23608 1234
rect 23634 1228 23637 1254
rect 24019 1248 24022 1254
rect 23999 1234 24022 1248
rect 24019 1228 24022 1234
rect 24048 1228 24051 1254
rect 24157 1248 24160 1254
rect 24137 1234 24160 1248
rect 24157 1228 24160 1234
rect 24186 1228 24189 1254
rect 32437 1228 32440 1254
rect 32466 1248 32469 1254
rect 32484 1249 32513 1252
rect 32484 1248 32490 1249
rect 32466 1234 32490 1248
rect 32466 1228 32469 1234
rect 32484 1232 32490 1234
rect 32507 1232 32513 1249
rect 32713 1248 32716 1254
rect 32693 1234 32716 1248
rect 32484 1229 32513 1232
rect 32713 1228 32716 1234
rect 32742 1228 32745 1254
rect 32989 1248 32992 1254
rect 32969 1234 32992 1248
rect 32989 1228 32992 1234
rect 33018 1228 33021 1254
rect 33127 1248 33130 1254
rect 33107 1234 33130 1248
rect 33127 1228 33130 1234
rect 33156 1228 33159 1254
rect 33266 1249 33295 1252
rect 33266 1232 33272 1249
rect 33289 1248 33295 1249
rect 33403 1248 33406 1254
rect 33289 1234 33406 1248
rect 33289 1232 33295 1234
rect 33266 1229 33295 1232
rect 33403 1228 33406 1234
rect 33432 1228 33435 1254
rect 1249 1194 1252 1220
rect 1278 1214 1281 1220
rect 1526 1215 1555 1218
rect 1526 1214 1532 1215
rect 1278 1200 1532 1214
rect 1278 1194 1281 1200
rect 1526 1198 1532 1200
rect 1549 1198 1555 1215
rect 1526 1195 1555 1198
rect 1893 1194 1896 1220
rect 1922 1214 1925 1220
rect 1922 1200 2284 1214
rect 1922 1194 1925 1200
rect 1111 1160 1114 1186
rect 1140 1180 1143 1186
rect 1663 1180 1666 1186
rect 1140 1166 1666 1180
rect 1140 1160 1143 1166
rect 1663 1160 1666 1166
rect 1692 1160 1695 1186
rect 1847 1160 1850 1186
rect 1876 1180 1879 1186
rect 1876 1166 1916 1180
rect 1876 1160 1879 1166
rect 421 1126 424 1152
rect 450 1146 453 1152
rect 1250 1147 1279 1150
rect 1250 1146 1256 1147
rect 450 1132 1256 1146
rect 450 1126 453 1132
rect 1250 1130 1256 1132
rect 1273 1130 1279 1147
rect 1250 1127 1279 1130
rect 1387 1126 1390 1152
rect 1416 1146 1419 1152
rect 1755 1146 1758 1152
rect 1416 1132 1758 1146
rect 1416 1126 1419 1132
rect 1755 1126 1758 1132
rect 1784 1126 1787 1152
rect 1801 1126 1804 1152
rect 1830 1146 1833 1152
rect 1902 1146 1916 1166
rect 1985 1160 1988 1186
rect 2014 1180 2017 1186
rect 2216 1181 2245 1184
rect 2216 1180 2222 1181
rect 2014 1166 2222 1180
rect 2014 1160 2017 1166
rect 2216 1164 2222 1166
rect 2239 1164 2245 1181
rect 2270 1180 2284 1200
rect 2353 1194 2356 1220
rect 2382 1214 2385 1220
rect 2768 1215 2797 1218
rect 2768 1214 2774 1215
rect 2382 1200 2774 1214
rect 2382 1194 2385 1200
rect 2768 1198 2774 1200
rect 2791 1198 2797 1215
rect 2768 1195 2797 1198
rect 2905 1194 2908 1220
rect 2934 1214 2937 1220
rect 3274 1215 3303 1218
rect 3274 1214 3280 1215
rect 2934 1200 3280 1214
rect 2934 1194 2937 1200
rect 3274 1198 3280 1200
rect 3297 1198 3303 1215
rect 3274 1195 3303 1198
rect 2492 1181 2521 1184
rect 2492 1180 2498 1181
rect 2270 1166 2498 1180
rect 2216 1161 2245 1164
rect 2492 1164 2498 1166
rect 2515 1164 2521 1181
rect 2492 1161 2521 1164
rect 2354 1147 2383 1150
rect 2354 1146 2360 1147
rect 1830 1132 1852 1146
rect 1902 1132 2360 1146
rect 1830 1126 1833 1132
rect 2354 1130 2360 1132
rect 2377 1130 2383 1147
rect 2354 1127 2383 1130
rect 2859 1126 2862 1152
rect 2888 1146 2891 1152
rect 2906 1147 2935 1150
rect 2906 1146 2912 1147
rect 2888 1132 2912 1146
rect 2888 1126 2891 1132
rect 2906 1130 2912 1132
rect 2929 1130 2935 1147
rect 2906 1127 2935 1130
rect 644 1101 34408 1112
rect 644 1075 6631 1101
rect 6657 1075 12631 1101
rect 12657 1075 18631 1101
rect 18657 1075 24631 1101
rect 24657 1075 30631 1101
rect 30657 1075 34408 1101
rect 644 1064 34408 1075
rect 1066 1045 1095 1048
rect 1066 1028 1072 1045
rect 1089 1044 1095 1045
rect 1479 1044 1482 1050
rect 1089 1030 1482 1044
rect 1089 1028 1095 1030
rect 1066 1025 1095 1028
rect 1479 1024 1482 1030
rect 1508 1024 1511 1050
rect 1525 1024 1528 1050
rect 1554 1044 1557 1050
rect 1940 1045 1969 1048
rect 1940 1044 1946 1045
rect 1554 1030 1946 1044
rect 1554 1024 1557 1030
rect 1940 1028 1946 1030
rect 1963 1028 1969 1045
rect 1940 1025 1969 1028
rect 2078 1045 2107 1048
rect 2078 1028 2084 1045
rect 2101 1044 2107 1045
rect 2123 1044 2126 1050
rect 2101 1030 2126 1044
rect 2101 1028 2107 1030
rect 2078 1025 2107 1028
rect 2123 1024 2126 1030
rect 2152 1024 2155 1050
rect 2353 1024 2356 1050
rect 2382 1044 2385 1050
rect 3274 1045 3303 1048
rect 3274 1044 3280 1045
rect 2382 1030 3280 1044
rect 2382 1024 2385 1030
rect 3274 1028 3280 1030
rect 3297 1028 3303 1045
rect 3411 1044 3414 1050
rect 3391 1030 3414 1044
rect 3274 1025 3303 1028
rect 3411 1024 3414 1030
rect 3440 1024 3443 1050
rect 1387 990 1390 1016
rect 1416 1010 1419 1016
rect 2216 1011 2245 1014
rect 2216 1010 2222 1011
rect 1416 996 2222 1010
rect 1416 990 1419 996
rect 2216 994 2222 996
rect 2239 994 2245 1011
rect 2216 991 2245 994
rect 2767 990 2770 1016
rect 2796 1010 2799 1016
rect 2906 1011 2935 1014
rect 2906 1010 2912 1011
rect 2796 996 2912 1010
rect 2796 990 2799 996
rect 2906 994 2912 996
rect 2929 994 2935 1011
rect 2906 991 2935 994
rect 559 956 562 982
rect 588 976 591 982
rect 1112 977 1141 980
rect 1112 976 1118 977
rect 588 962 1118 976
rect 588 956 591 962
rect 1112 960 1118 962
rect 1135 960 1141 977
rect 1112 957 1141 960
rect 1166 962 1410 976
rect 697 888 700 914
rect 726 908 729 914
rect 1166 908 1180 962
rect 1396 946 1410 962
rect 1433 956 1436 982
rect 1462 976 1465 982
rect 2354 977 2383 980
rect 2354 976 2360 977
rect 1462 962 2360 976
rect 1462 956 1465 962
rect 2354 960 2360 962
rect 2377 960 2383 977
rect 2354 957 2383 960
rect 2675 956 2678 982
rect 2704 976 2707 982
rect 3044 977 3073 980
rect 3044 976 3050 977
rect 2704 962 3050 976
rect 2704 956 2707 962
rect 3044 960 3050 962
rect 3067 960 3073 977
rect 3044 957 3073 960
rect 22501 956 22504 982
rect 22530 976 22533 982
rect 23054 977 23083 980
rect 23054 976 23060 977
rect 22530 962 23060 976
rect 22530 956 22533 962
rect 23054 960 23060 962
rect 23077 960 23083 977
rect 23054 957 23083 960
rect 1342 943 1371 946
rect 1342 926 1348 943
rect 1365 926 1371 943
rect 1342 923 1371 926
rect 1388 943 1417 946
rect 1388 926 1394 943
rect 1411 926 1417 943
rect 1525 942 1528 948
rect 1505 928 1528 942
rect 1388 923 1417 926
rect 726 894 1180 908
rect 726 888 729 894
rect 1350 874 1364 923
rect 1525 922 1528 928
rect 1554 922 1557 948
rect 1663 942 1666 948
rect 1643 928 1666 942
rect 1663 922 1666 928
rect 1692 922 1695 948
rect 1755 922 1758 948
rect 1784 942 1787 948
rect 1802 943 1831 946
rect 1802 942 1808 943
rect 1784 928 1808 942
rect 1784 922 1787 928
rect 1802 926 1808 928
rect 1825 926 1831 943
rect 1802 923 1831 926
rect 2492 943 2521 946
rect 2492 926 2498 943
rect 2515 926 2521 943
rect 2492 923 2521 926
rect 1479 888 1482 914
rect 1508 908 1511 914
rect 2500 908 2514 923
rect 2583 922 2586 948
rect 2612 942 2615 948
rect 2630 943 2659 946
rect 2630 942 2636 943
rect 2612 928 2636 942
rect 2612 922 2615 928
rect 2630 926 2636 928
rect 2653 926 2659 943
rect 2630 923 2659 926
rect 2768 943 2797 946
rect 2768 926 2774 943
rect 2791 942 2797 943
rect 2951 942 2954 948
rect 2791 928 2954 942
rect 2791 926 2797 928
rect 2768 923 2797 926
rect 2951 922 2954 928
rect 2980 922 2983 948
rect 3457 922 3460 948
rect 3486 942 3489 948
rect 3642 943 3671 946
rect 3642 942 3648 943
rect 3486 928 3648 942
rect 3486 922 3489 928
rect 3642 926 3648 928
rect 3665 926 3671 943
rect 3642 923 3671 926
rect 4699 922 4702 948
rect 4728 942 4731 948
rect 4930 943 4959 946
rect 4930 942 4936 943
rect 4728 928 4936 942
rect 4728 922 4731 928
rect 4930 926 4936 928
rect 4953 926 4959 943
rect 4930 923 4959 926
rect 5803 922 5806 948
rect 5832 942 5835 948
rect 6080 943 6109 946
rect 6080 942 6086 943
rect 5832 928 6086 942
rect 5832 922 5835 928
rect 6080 926 6086 928
rect 6103 926 6109 943
rect 6080 923 6109 926
rect 6769 922 6772 948
rect 6798 942 6801 948
rect 7046 943 7075 946
rect 7046 942 7052 943
rect 6798 928 7052 942
rect 6798 922 6801 928
rect 7046 926 7052 928
rect 7069 926 7075 943
rect 7046 923 7075 926
rect 8057 922 8060 948
rect 8086 942 8089 948
rect 8426 943 8455 946
rect 8426 942 8432 943
rect 8086 928 8432 942
rect 8086 922 8089 928
rect 8426 926 8432 928
rect 8449 926 8455 943
rect 8426 923 8455 926
rect 9805 922 9808 948
rect 9834 942 9837 948
rect 10128 943 10157 946
rect 10128 942 10134 943
rect 9834 928 10134 942
rect 9834 922 9837 928
rect 10128 926 10134 928
rect 10151 926 10157 943
rect 10128 923 10157 926
rect 10771 922 10774 948
rect 10800 942 10803 948
rect 11094 943 11123 946
rect 11094 942 11100 943
rect 10800 928 11100 942
rect 10800 922 10803 928
rect 11094 926 11100 928
rect 11117 926 11123 943
rect 11094 923 11123 926
rect 12151 922 12154 948
rect 12180 942 12183 948
rect 12520 943 12549 946
rect 12520 942 12526 943
rect 12180 928 12526 942
rect 12180 922 12183 928
rect 12520 926 12526 928
rect 12543 926 12549 943
rect 12520 923 12549 926
rect 14221 922 14224 948
rect 14250 942 14253 948
rect 14636 943 14665 946
rect 14636 942 14642 943
rect 14250 928 14642 942
rect 14250 922 14253 928
rect 14636 926 14642 928
rect 14659 926 14665 943
rect 14636 923 14665 926
rect 15325 922 15328 948
rect 15354 942 15357 948
rect 15740 943 15769 946
rect 15740 942 15746 943
rect 15354 928 15746 942
rect 15354 922 15357 928
rect 15740 926 15746 928
rect 15763 926 15769 943
rect 15740 923 15769 926
rect 15877 922 15880 948
rect 15906 942 15909 948
rect 16292 943 16321 946
rect 16292 942 16298 943
rect 15906 928 16298 942
rect 15906 922 15909 928
rect 16292 926 16298 928
rect 16315 926 16321 943
rect 16292 923 16321 926
rect 21719 922 21722 948
rect 21748 942 21751 948
rect 22180 943 22209 946
rect 22180 942 22186 943
rect 21748 928 22186 942
rect 21748 922 21751 928
rect 22180 926 22186 928
rect 22203 926 22209 943
rect 22180 923 22209 926
rect 22225 922 22228 948
rect 22254 942 22257 948
rect 22778 943 22807 946
rect 22778 942 22784 943
rect 22254 928 22784 942
rect 22254 922 22257 928
rect 22778 926 22784 928
rect 22801 926 22807 943
rect 22778 923 22807 926
rect 25537 922 25540 948
rect 25566 942 25569 948
rect 26136 943 26165 946
rect 26136 942 26142 943
rect 25566 928 26142 942
rect 25566 922 25569 928
rect 26136 926 26142 928
rect 26159 926 26165 943
rect 26136 923 26165 926
rect 1508 894 2514 908
rect 1508 888 1511 894
rect 1939 874 1942 880
rect 1350 860 1942 874
rect 1939 854 1942 860
rect 1968 854 1971 880
rect 644 829 34408 840
rect 644 803 3631 829
rect 3657 803 9631 829
rect 9657 803 15631 829
rect 15657 803 21631 829
rect 21657 803 27631 829
rect 27657 803 33631 829
rect 33657 803 34408 829
rect 644 792 34408 803
rect 1111 684 1114 710
rect 1140 704 1143 710
rect 1140 690 1318 704
rect 1140 684 1143 690
rect 1066 671 1095 674
rect 1066 654 1072 671
rect 1089 670 1095 671
rect 1203 670 1206 676
rect 1089 656 1206 670
rect 1089 654 1095 656
rect 1066 651 1095 654
rect 1203 650 1206 656
rect 1232 650 1235 676
rect 1304 670 1318 690
rect 1571 684 1574 710
rect 1600 704 1603 710
rect 1801 704 1804 710
rect 1600 690 1804 704
rect 1600 684 1603 690
rect 1801 684 1804 690
rect 1830 684 1833 710
rect 13255 684 13258 710
rect 13284 704 13287 710
rect 13900 705 13929 708
rect 13900 704 13906 705
rect 13284 690 13906 704
rect 13284 684 13287 690
rect 13900 688 13906 690
rect 13923 688 13929 705
rect 13900 685 13929 688
rect 13945 684 13948 710
rect 13974 704 13977 710
rect 13974 690 14106 704
rect 13974 684 13977 690
rect 1526 671 1555 674
rect 1526 670 1532 671
rect 1304 656 1532 670
rect 1526 654 1532 656
rect 1549 654 1555 671
rect 1526 651 1555 654
rect 1893 650 1896 676
rect 1922 670 1925 676
rect 2354 671 2383 674
rect 2354 670 2360 671
rect 1922 656 2360 670
rect 1922 650 1925 656
rect 2354 654 2360 656
rect 2377 654 2383 671
rect 2354 651 2383 654
rect 2491 650 2494 676
rect 2520 670 2523 676
rect 2768 671 2797 674
rect 2768 670 2774 671
rect 2520 656 2774 670
rect 2520 650 2523 656
rect 2768 654 2774 656
rect 2791 654 2797 671
rect 2768 651 2797 654
rect 2813 650 2816 676
rect 2842 670 2845 676
rect 2906 671 2935 674
rect 2906 670 2912 671
rect 2842 656 2912 670
rect 2842 650 2845 656
rect 2906 654 2912 656
rect 2929 654 2935 671
rect 2906 651 2935 654
rect 3319 650 3322 676
rect 3348 670 3351 676
rect 3596 671 3625 674
rect 3596 670 3602 671
rect 3348 656 3602 670
rect 3348 650 3351 656
rect 3596 654 3602 656
rect 3619 654 3625 671
rect 3596 651 3625 654
rect 3733 650 3736 676
rect 3762 670 3765 676
rect 3918 671 3947 674
rect 3918 670 3924 671
rect 3762 656 3924 670
rect 3762 650 3765 656
rect 3918 654 3924 656
rect 3941 654 3947 671
rect 3918 651 3947 654
rect 4837 650 4840 676
rect 4866 670 4869 676
rect 5068 671 5097 674
rect 5068 670 5074 671
rect 4866 656 5074 670
rect 4866 650 4869 656
rect 5068 654 5074 656
rect 5091 654 5097 671
rect 5068 651 5097 654
rect 5665 650 5668 676
rect 5694 670 5697 676
rect 5988 671 6017 674
rect 5988 670 5994 671
rect 5694 656 5994 670
rect 5694 650 5697 656
rect 5988 654 5994 656
rect 6011 654 6017 671
rect 5988 651 6017 654
rect 6493 650 6496 676
rect 6522 670 6525 676
rect 6770 671 6799 674
rect 6770 670 6776 671
rect 6522 656 6776 670
rect 6522 650 6525 656
rect 6770 654 6776 656
rect 6793 654 6799 671
rect 6770 651 6799 654
rect 6907 650 6910 676
rect 6936 670 6939 676
rect 7184 671 7213 674
rect 7184 670 7190 671
rect 6936 656 7190 670
rect 6936 650 6939 656
rect 7184 654 7190 656
rect 7207 654 7213 671
rect 7184 651 7213 654
rect 7873 650 7876 676
rect 7902 670 7905 676
rect 8150 671 8179 674
rect 8150 670 8156 671
rect 7902 656 8156 670
rect 7902 650 7905 656
rect 8150 654 8156 656
rect 8173 654 8179 671
rect 8150 651 8179 654
rect 8425 650 8428 676
rect 8454 670 8457 676
rect 8748 671 8777 674
rect 8748 670 8754 671
rect 8454 656 8754 670
rect 8454 650 8457 656
rect 8748 654 8754 656
rect 8771 654 8777 671
rect 8748 651 8777 654
rect 8839 650 8842 676
rect 8868 670 8871 676
rect 9162 671 9191 674
rect 9162 670 9168 671
rect 8868 656 9168 670
rect 8868 650 8871 656
rect 9162 654 9168 656
rect 9185 654 9191 671
rect 9162 651 9191 654
rect 9713 650 9716 676
rect 9742 670 9745 676
rect 9990 671 10019 674
rect 9990 670 9996 671
rect 9742 656 9996 670
rect 9742 650 9745 656
rect 9990 654 9996 656
rect 10013 654 10019 671
rect 9990 651 10019 654
rect 10081 650 10084 676
rect 10110 670 10113 676
rect 10404 671 10433 674
rect 10404 670 10410 671
rect 10110 656 10410 670
rect 10110 650 10113 656
rect 10404 654 10410 656
rect 10427 654 10433 671
rect 10404 651 10433 654
rect 10495 650 10498 676
rect 10524 670 10527 676
rect 10818 671 10847 674
rect 10818 670 10824 671
rect 10524 656 10824 670
rect 10524 650 10527 656
rect 10818 654 10824 656
rect 10841 654 10847 671
rect 10818 651 10847 654
rect 11185 650 11188 676
rect 11214 670 11217 676
rect 11508 671 11537 674
rect 11508 670 11514 671
rect 11214 656 11514 670
rect 11214 650 11217 656
rect 11508 654 11514 656
rect 11531 654 11537 671
rect 11508 651 11537 654
rect 11737 650 11740 676
rect 11766 670 11769 676
rect 12106 671 12135 674
rect 12106 670 12112 671
rect 11766 656 12112 670
rect 11766 650 11769 656
rect 12106 654 12112 656
rect 12129 654 12135 671
rect 12106 651 12135 654
rect 12427 650 12430 676
rect 12456 670 12459 676
rect 12796 671 12825 674
rect 12796 670 12802 671
rect 12456 656 12802 670
rect 12456 650 12459 656
rect 12796 654 12802 656
rect 12819 654 12825 671
rect 12796 651 12825 654
rect 12979 650 12982 676
rect 13008 670 13011 676
rect 13348 671 13377 674
rect 13348 670 13354 671
rect 13008 656 13354 670
rect 13008 650 13011 656
rect 13348 654 13354 656
rect 13371 654 13377 671
rect 13348 651 13377 654
rect 13669 650 13672 676
rect 13698 670 13701 676
rect 14038 671 14067 674
rect 14038 670 14044 671
rect 13698 656 14044 670
rect 13698 650 13701 656
rect 14038 654 14044 656
rect 14061 654 14067 671
rect 14092 670 14106 690
rect 19465 684 19468 710
rect 19494 704 19497 710
rect 20202 705 20231 708
rect 20202 704 20208 705
rect 19494 690 20208 704
rect 19494 684 19497 690
rect 20202 688 20208 690
rect 20225 688 20231 705
rect 20202 685 20231 688
rect 20707 684 20710 710
rect 20736 704 20739 710
rect 20736 690 21006 704
rect 20736 684 20739 690
rect 14590 671 14619 674
rect 14590 670 14596 671
rect 14092 656 14596 670
rect 14038 651 14067 654
rect 14590 654 14596 656
rect 14613 654 14619 671
rect 14590 651 14619 654
rect 14773 650 14776 676
rect 14802 670 14805 676
rect 15188 671 15217 674
rect 15188 670 15194 671
rect 14802 656 15194 670
rect 14802 650 14805 656
rect 15188 654 15194 656
rect 15211 654 15217 671
rect 15188 651 15217 654
rect 15463 650 15466 676
rect 15492 670 15495 676
rect 15878 671 15907 674
rect 15878 670 15884 671
rect 15492 656 15884 670
rect 15492 650 15495 656
rect 15878 654 15884 656
rect 15901 654 15907 671
rect 15878 651 15907 654
rect 16153 650 16156 676
rect 16182 670 16185 676
rect 16568 671 16597 674
rect 16568 670 16574 671
rect 16182 656 16574 670
rect 16182 650 16185 656
rect 16568 654 16574 656
rect 16591 654 16597 671
rect 16568 651 16597 654
rect 16613 650 16616 676
rect 16642 670 16645 676
rect 16982 671 17011 674
rect 16982 670 16988 671
rect 16642 656 16988 670
rect 16642 650 16645 656
rect 16982 654 16988 656
rect 17005 654 17011 671
rect 16982 651 17011 654
rect 17027 650 17030 676
rect 17056 670 17059 676
rect 17442 671 17471 674
rect 17442 670 17448 671
rect 17056 656 17448 670
rect 17056 650 17059 656
rect 17442 654 17448 656
rect 17465 654 17471 671
rect 17718 671 17747 674
rect 17718 670 17724 671
rect 17442 651 17471 654
rect 17496 656 17724 670
rect 973 616 976 642
rect 1002 636 1005 642
rect 1250 637 1279 640
rect 1250 636 1256 637
rect 1002 622 1256 636
rect 1002 616 1005 622
rect 1250 620 1256 622
rect 1273 620 1279 637
rect 1617 636 1620 642
rect 1250 617 1279 620
rect 1350 622 1620 636
rect 927 602 930 608
rect 907 588 930 602
rect 927 582 930 588
rect 956 582 959 608
rect 1204 603 1233 606
rect 1204 586 1210 603
rect 1227 602 1233 603
rect 1350 602 1364 622
rect 1617 616 1620 622
rect 1646 616 1649 642
rect 1755 616 1758 642
rect 1784 636 1787 642
rect 2216 637 2245 640
rect 2216 636 2222 637
rect 1784 622 2222 636
rect 1784 616 1787 622
rect 2216 620 2222 622
rect 2239 620 2245 637
rect 2216 617 2245 620
rect 2261 616 2264 642
rect 2290 636 2293 642
rect 3044 637 3073 640
rect 3044 636 3050 637
rect 2290 622 3050 636
rect 2290 616 2293 622
rect 3044 620 3050 622
rect 3067 620 3073 637
rect 3044 617 3073 620
rect 3089 616 3092 642
rect 3118 636 3121 642
rect 3458 637 3487 640
rect 3458 636 3464 637
rect 3118 622 3464 636
rect 3118 616 3121 622
rect 3458 620 3464 622
rect 3481 620 3487 637
rect 3458 617 3487 620
rect 3871 616 3874 642
rect 3900 636 3903 642
rect 4056 637 4085 640
rect 4056 636 4062 637
rect 3900 622 4062 636
rect 3900 616 3903 622
rect 4056 620 4062 622
rect 4079 620 4085 637
rect 4056 617 4085 620
rect 4147 616 4150 642
rect 4176 636 4179 642
rect 4378 637 4407 640
rect 4378 636 4384 637
rect 4176 622 4384 636
rect 4176 616 4179 622
rect 4378 620 4384 622
rect 4401 620 4407 637
rect 4378 617 4407 620
rect 4423 616 4426 642
rect 4452 636 4455 642
rect 4700 637 4729 640
rect 4700 636 4706 637
rect 4452 622 4706 636
rect 4452 616 4455 622
rect 4700 620 4706 622
rect 4723 620 4729 637
rect 4700 617 4729 620
rect 5113 616 5116 642
rect 5142 636 5145 642
rect 5344 637 5373 640
rect 5344 636 5350 637
rect 5142 622 5350 636
rect 5142 616 5145 622
rect 5344 620 5350 622
rect 5367 620 5373 637
rect 5344 617 5373 620
rect 5389 616 5392 642
rect 5418 636 5421 642
rect 5620 637 5649 640
rect 5620 636 5626 637
rect 5418 622 5626 636
rect 5418 616 5421 622
rect 5620 620 5626 622
rect 5643 620 5649 637
rect 5620 617 5649 620
rect 5941 616 5944 642
rect 5970 636 5973 642
rect 6218 637 6247 640
rect 6218 636 6224 637
rect 5970 622 6224 636
rect 5970 616 5973 622
rect 6218 620 6224 622
rect 6241 620 6247 637
rect 6218 617 6247 620
rect 6401 616 6404 642
rect 6430 636 6433 642
rect 6632 637 6661 640
rect 6632 636 6638 637
rect 6430 622 6638 636
rect 6430 616 6433 622
rect 6632 620 6638 622
rect 6655 620 6661 637
rect 6632 617 6661 620
rect 7045 616 7048 642
rect 7074 636 7077 642
rect 7322 637 7351 640
rect 7322 636 7328 637
rect 7074 622 7328 636
rect 7074 616 7077 622
rect 7322 620 7328 622
rect 7345 620 7351 637
rect 7322 617 7351 620
rect 7367 616 7370 642
rect 7396 636 7399 642
rect 7598 637 7627 640
rect 7598 636 7604 637
rect 7396 622 7604 636
rect 7396 616 7399 622
rect 7598 620 7604 622
rect 7621 620 7627 637
rect 7598 617 7627 620
rect 7643 616 7646 642
rect 7672 636 7675 642
rect 7672 622 7896 636
rect 7672 616 7675 622
rect 1227 588 1364 602
rect 1227 586 1233 588
rect 1204 583 1233 586
rect 1387 582 1390 608
rect 1416 602 1419 608
rect 1663 602 1666 608
rect 1416 588 1438 602
rect 1643 588 1666 602
rect 1416 582 1419 588
rect 1663 582 1666 588
rect 1692 582 1695 608
rect 1709 582 1712 608
rect 1738 602 1741 608
rect 1802 603 1831 606
rect 1802 602 1808 603
rect 1738 588 1808 602
rect 1738 582 1741 588
rect 1802 586 1808 588
rect 1825 586 1831 603
rect 1802 583 1831 586
rect 1847 582 1850 608
rect 1876 602 1879 608
rect 2078 603 2107 606
rect 2078 602 2084 603
rect 1876 588 2084 602
rect 1876 582 1879 588
rect 2078 586 2084 588
rect 2101 586 2107 603
rect 2078 583 2107 586
rect 2123 582 2126 608
rect 2152 602 2155 608
rect 2492 603 2521 606
rect 2492 602 2498 603
rect 2152 588 2498 602
rect 2152 582 2155 588
rect 2492 586 2498 588
rect 2515 586 2521 603
rect 2492 583 2521 586
rect 2537 582 2540 608
rect 2566 602 2569 608
rect 2630 603 2659 606
rect 2630 602 2636 603
rect 2566 588 2636 602
rect 2566 582 2569 588
rect 2630 586 2636 588
rect 2653 586 2659 603
rect 2630 583 2659 586
rect 3181 582 3184 608
rect 3210 602 3213 608
rect 3320 603 3349 606
rect 3320 602 3326 603
rect 3210 588 3326 602
rect 3210 582 3213 588
rect 3320 586 3326 588
rect 3343 586 3349 603
rect 3320 583 3349 586
rect 3687 582 3690 608
rect 3716 602 3719 608
rect 3780 603 3809 606
rect 3780 602 3786 603
rect 3716 588 3786 602
rect 3716 582 3719 588
rect 3780 586 3786 588
rect 3803 586 3809 603
rect 3780 583 3809 586
rect 4009 582 4012 608
rect 4038 602 4041 608
rect 4240 603 4269 606
rect 4240 602 4246 603
rect 4038 588 4246 602
rect 4038 582 4041 588
rect 4240 586 4246 588
rect 4263 586 4269 603
rect 4240 583 4269 586
rect 4285 582 4288 608
rect 4314 602 4317 608
rect 4562 603 4591 606
rect 4562 602 4568 603
rect 4314 588 4568 602
rect 4314 582 4317 588
rect 4562 586 4568 588
rect 4585 586 4591 603
rect 4562 583 4591 586
rect 4607 582 4610 608
rect 4636 602 4639 608
rect 4838 603 4867 606
rect 4838 602 4844 603
rect 4636 588 4844 602
rect 4636 582 4639 588
rect 4838 586 4844 588
rect 4861 586 4867 603
rect 4838 583 4867 586
rect 4975 582 4978 608
rect 5004 602 5007 608
rect 5206 603 5235 606
rect 5206 602 5212 603
rect 5004 588 5212 602
rect 5004 582 5007 588
rect 5206 586 5212 588
rect 5229 586 5235 603
rect 5206 583 5235 586
rect 5251 582 5254 608
rect 5280 602 5283 608
rect 5482 603 5511 606
rect 5482 602 5488 603
rect 5280 588 5488 602
rect 5280 582 5283 588
rect 5482 586 5488 588
rect 5505 586 5511 603
rect 5482 583 5511 586
rect 5527 582 5530 608
rect 5556 602 5559 608
rect 5850 603 5879 606
rect 5850 602 5856 603
rect 5556 588 5856 602
rect 5556 582 5559 588
rect 5850 586 5856 588
rect 5873 586 5879 603
rect 5850 583 5879 586
rect 6079 582 6082 608
rect 6108 602 6111 608
rect 6356 603 6385 606
rect 6356 602 6362 603
rect 6108 588 6362 602
rect 6108 582 6111 588
rect 6356 586 6362 588
rect 6379 586 6385 603
rect 6356 583 6385 586
rect 6447 582 6450 608
rect 6476 602 6479 608
rect 6494 603 6523 606
rect 6494 602 6500 603
rect 6476 588 6500 602
rect 6476 582 6479 588
rect 6494 586 6500 588
rect 6517 586 6523 603
rect 6494 583 6523 586
rect 6723 582 6726 608
rect 6752 602 6755 608
rect 6908 603 6937 606
rect 6908 602 6914 603
rect 6752 588 6914 602
rect 6752 582 6755 588
rect 6908 586 6914 588
rect 6931 586 6937 603
rect 6908 583 6937 586
rect 7183 582 7186 608
rect 7212 602 7215 608
rect 7460 603 7489 606
rect 7460 602 7466 603
rect 7212 588 7466 602
rect 7212 582 7215 588
rect 7460 586 7466 588
rect 7483 586 7489 603
rect 7460 583 7489 586
rect 7505 582 7508 608
rect 7534 602 7537 608
rect 7882 606 7896 622
rect 8287 616 8290 642
rect 8316 636 8319 642
rect 8610 637 8639 640
rect 8610 636 8616 637
rect 8316 622 8616 636
rect 8316 616 8319 622
rect 8610 620 8616 622
rect 8633 620 8639 637
rect 8610 617 8639 620
rect 8701 616 8704 642
rect 8730 636 8733 642
rect 8730 622 8954 636
rect 8730 616 8733 622
rect 7736 603 7765 606
rect 7736 602 7742 603
rect 7534 588 7742 602
rect 7534 582 7537 588
rect 7736 586 7742 588
rect 7759 586 7765 603
rect 7736 583 7765 586
rect 7874 603 7903 606
rect 7874 586 7880 603
rect 7897 586 7903 603
rect 8011 602 8014 608
rect 7991 588 8014 602
rect 7874 583 7903 586
rect 8011 582 8014 588
rect 8040 582 8043 608
rect 8195 582 8198 608
rect 8224 602 8227 608
rect 8426 603 8455 606
rect 8426 602 8432 603
rect 8224 588 8432 602
rect 8224 582 8227 588
rect 8426 586 8432 588
rect 8449 586 8455 603
rect 8426 583 8455 586
rect 8563 582 8566 608
rect 8592 602 8595 608
rect 8886 603 8915 606
rect 8886 602 8892 603
rect 8592 588 8892 602
rect 8592 582 8595 588
rect 8886 586 8892 588
rect 8909 586 8915 603
rect 8940 602 8954 622
rect 8977 616 8980 642
rect 9006 636 9009 642
rect 9300 637 9329 640
rect 9300 636 9306 637
rect 9006 622 9306 636
rect 9006 616 9009 622
rect 9300 620 9306 622
rect 9323 620 9329 637
rect 9300 617 9329 620
rect 9529 616 9532 642
rect 9558 636 9561 642
rect 9852 637 9881 640
rect 9852 636 9858 637
rect 9558 622 9858 636
rect 9558 616 9561 622
rect 9852 620 9858 622
rect 9875 620 9881 637
rect 9852 617 9881 620
rect 9943 616 9946 642
rect 9972 636 9975 642
rect 10266 637 10295 640
rect 10266 636 10272 637
rect 9972 622 10272 636
rect 9972 616 9975 622
rect 10266 620 10272 622
rect 10289 620 10295 637
rect 10266 617 10295 620
rect 10357 616 10360 642
rect 10386 636 10389 642
rect 10680 637 10709 640
rect 10680 636 10686 637
rect 10386 622 10686 636
rect 10386 616 10389 622
rect 10680 620 10686 622
rect 10703 620 10709 637
rect 10680 617 10709 620
rect 10909 616 10912 642
rect 10938 636 10941 642
rect 11232 637 11261 640
rect 11232 636 11238 637
rect 10938 622 11238 636
rect 10938 616 10941 622
rect 11232 620 11238 622
rect 11255 620 11261 637
rect 11232 617 11261 620
rect 11323 616 11326 642
rect 11352 636 11355 642
rect 11352 622 11438 636
rect 11352 616 11355 622
rect 9024 603 9053 606
rect 9024 602 9030 603
rect 8940 588 9030 602
rect 8886 583 8915 586
rect 9024 586 9030 588
rect 9047 586 9053 603
rect 9024 583 9053 586
rect 9115 582 9118 608
rect 9144 602 9147 608
rect 9438 603 9467 606
rect 9438 602 9444 603
rect 9144 588 9444 602
rect 9144 582 9147 588
rect 9438 586 9444 588
rect 9461 586 9467 603
rect 9438 583 9467 586
rect 9483 582 9486 608
rect 9512 602 9515 608
rect 9714 603 9743 606
rect 9714 602 9720 603
rect 9512 588 9720 602
rect 9512 582 9515 588
rect 9714 586 9720 588
rect 9737 586 9743 603
rect 10127 602 10130 608
rect 10107 588 10130 602
rect 9714 583 9743 586
rect 10127 582 10130 588
rect 10156 582 10159 608
rect 10311 582 10314 608
rect 10340 602 10343 608
rect 10542 603 10571 606
rect 10542 602 10548 603
rect 10340 588 10548 602
rect 10340 582 10343 588
rect 10542 586 10548 588
rect 10565 586 10571 603
rect 10542 583 10571 586
rect 10633 582 10636 608
rect 10662 602 10665 608
rect 11002 603 11031 606
rect 11002 602 11008 603
rect 10662 588 11008 602
rect 10662 582 10665 588
rect 11002 586 11008 588
rect 11025 586 11031 603
rect 11002 583 11031 586
rect 11047 582 11050 608
rect 11076 602 11079 608
rect 11370 603 11399 606
rect 11370 602 11376 603
rect 11076 588 11376 602
rect 11076 582 11079 588
rect 11370 586 11376 588
rect 11393 586 11399 603
rect 11424 602 11438 622
rect 11461 616 11464 642
rect 11490 636 11493 642
rect 11784 637 11813 640
rect 11784 636 11790 637
rect 11490 622 11790 636
rect 11490 616 11493 622
rect 11784 620 11790 622
rect 11807 620 11813 637
rect 11784 617 11813 620
rect 11875 616 11878 642
rect 11904 636 11907 642
rect 12290 637 12319 640
rect 12290 636 12296 637
rect 11904 622 12296 636
rect 11904 616 11907 622
rect 12290 620 12296 622
rect 12313 620 12319 637
rect 12290 617 12319 620
rect 12335 616 12338 642
rect 12364 636 12367 642
rect 12658 637 12687 640
rect 12658 636 12664 637
rect 12364 622 12664 636
rect 12364 616 12367 622
rect 12658 620 12664 622
rect 12681 620 12687 637
rect 12658 617 12687 620
rect 12841 616 12844 642
rect 12870 636 12873 642
rect 13210 637 13239 640
rect 13210 636 13216 637
rect 12870 622 13216 636
rect 12870 616 12873 622
rect 13210 620 13216 622
rect 13233 620 13239 637
rect 13210 617 13239 620
rect 13393 616 13396 642
rect 13422 636 13425 642
rect 13762 637 13791 640
rect 13762 636 13768 637
rect 13422 622 13768 636
rect 13422 616 13425 622
rect 13762 620 13768 622
rect 13785 620 13791 637
rect 13762 617 13791 620
rect 13807 616 13810 642
rect 13836 636 13839 642
rect 13836 622 13968 636
rect 13836 616 13839 622
rect 11646 603 11675 606
rect 11646 602 11652 603
rect 11424 588 11652 602
rect 11370 583 11399 586
rect 11646 586 11652 588
rect 11669 586 11675 603
rect 11646 583 11675 586
rect 11691 582 11694 608
rect 11720 602 11723 608
rect 11968 603 11997 606
rect 11968 602 11974 603
rect 11720 588 11974 602
rect 11720 582 11723 588
rect 11968 586 11974 588
rect 11991 586 11997 603
rect 11968 583 11997 586
rect 12013 582 12016 608
rect 12042 602 12045 608
rect 12428 603 12457 606
rect 12428 602 12434 603
rect 12042 588 12434 602
rect 12042 582 12045 588
rect 12428 586 12434 588
rect 12451 586 12457 603
rect 12428 583 12457 586
rect 12565 582 12568 608
rect 12594 602 12597 608
rect 12934 603 12963 606
rect 12934 602 12940 603
rect 12594 588 12940 602
rect 12594 582 12597 588
rect 12934 586 12940 588
rect 12957 586 12963 603
rect 13071 602 13074 608
rect 13051 588 13074 602
rect 12934 583 12963 586
rect 13071 582 13074 588
rect 13100 582 13103 608
rect 13117 582 13120 608
rect 13146 602 13149 608
rect 13578 603 13607 606
rect 13578 602 13584 603
rect 13146 588 13584 602
rect 13146 582 13149 588
rect 13578 586 13584 588
rect 13601 586 13607 603
rect 13954 602 13968 622
rect 14083 616 14086 642
rect 14112 636 14115 642
rect 14452 637 14481 640
rect 14452 636 14458 637
rect 14112 622 14458 636
rect 14112 616 14115 622
rect 14452 620 14458 622
rect 14475 620 14481 637
rect 14452 617 14481 620
rect 14497 616 14500 642
rect 14526 636 14529 642
rect 14912 637 14941 640
rect 14912 636 14918 637
rect 14526 622 14918 636
rect 14526 616 14529 622
rect 14912 620 14918 622
rect 14935 620 14941 637
rect 14912 617 14941 620
rect 14957 616 14960 642
rect 14986 636 14989 642
rect 15326 637 15355 640
rect 15326 636 15332 637
rect 14986 622 15332 636
rect 14986 616 14989 622
rect 15326 620 15332 622
rect 15349 620 15355 637
rect 15602 637 15631 640
rect 15602 636 15608 637
rect 15326 617 15355 620
rect 15380 622 15608 636
rect 14176 603 14205 606
rect 14176 602 14182 603
rect 13954 588 14182 602
rect 13578 583 13607 586
rect 14176 586 14182 588
rect 14199 586 14205 603
rect 14313 602 14316 608
rect 14293 588 14316 602
rect 14176 583 14205 586
rect 14313 582 14316 588
rect 14342 582 14345 608
rect 14359 582 14362 608
rect 14388 602 14391 608
rect 15050 603 15079 606
rect 15050 602 15056 603
rect 14388 588 15056 602
rect 14388 582 14391 588
rect 15050 586 15056 588
rect 15073 586 15079 603
rect 15050 583 15079 586
rect 15187 582 15190 608
rect 15216 602 15219 608
rect 15380 602 15394 622
rect 15602 620 15608 622
rect 15625 620 15631 637
rect 15602 617 15631 620
rect 16015 616 16018 642
rect 16044 636 16047 642
rect 16430 637 16459 640
rect 16430 636 16436 637
rect 16044 622 16436 636
rect 16044 616 16047 622
rect 16430 620 16436 622
rect 16453 620 16459 637
rect 16430 617 16459 620
rect 16475 616 16478 642
rect 16504 636 16507 642
rect 16844 637 16873 640
rect 16844 636 16850 637
rect 16504 622 16850 636
rect 16504 616 16507 622
rect 16844 620 16850 622
rect 16867 620 16873 637
rect 16844 617 16873 620
rect 16889 616 16892 642
rect 16918 636 16921 642
rect 17258 637 17287 640
rect 17258 636 17264 637
rect 16918 622 17264 636
rect 16918 616 16921 622
rect 17258 620 17264 622
rect 17281 620 17287 637
rect 17258 617 17287 620
rect 17303 616 17306 642
rect 17332 636 17335 642
rect 17496 636 17510 656
rect 17718 654 17724 656
rect 17741 654 17747 671
rect 17718 651 17747 654
rect 17809 650 17812 676
rect 17838 670 17841 676
rect 18270 671 18299 674
rect 18270 670 18276 671
rect 17838 656 18276 670
rect 17838 650 17841 656
rect 18270 654 18276 656
rect 18293 654 18299 671
rect 18270 651 18299 654
rect 18315 650 18318 676
rect 18344 670 18347 676
rect 18730 671 18759 674
rect 18730 670 18736 671
rect 18344 656 18736 670
rect 18344 650 18347 656
rect 18730 654 18736 656
rect 18753 654 18759 671
rect 18730 651 18759 654
rect 18775 650 18778 676
rect 18804 670 18807 676
rect 19144 671 19173 674
rect 19144 670 19150 671
rect 18804 656 19150 670
rect 18804 650 18807 656
rect 19144 654 19150 656
rect 19167 654 19173 671
rect 19144 651 19173 654
rect 19189 650 19192 676
rect 19218 670 19221 676
rect 19558 671 19587 674
rect 19558 670 19564 671
rect 19218 656 19564 670
rect 19218 650 19221 656
rect 19558 654 19564 656
rect 19581 654 19587 671
rect 19558 651 19587 654
rect 19741 650 19744 676
rect 19770 670 19773 676
rect 20340 671 20369 674
rect 20340 670 20346 671
rect 19770 656 20346 670
rect 19770 650 19773 656
rect 20340 654 20346 656
rect 20363 654 20369 671
rect 20340 651 20369 654
rect 20385 650 20388 676
rect 20414 670 20417 676
rect 20892 671 20921 674
rect 20892 670 20898 671
rect 20414 656 20898 670
rect 20414 650 20417 656
rect 20892 654 20898 656
rect 20915 654 20921 671
rect 20992 670 21006 690
rect 22915 684 22918 710
rect 22944 704 22947 710
rect 23468 705 23497 708
rect 23468 704 23474 705
rect 22944 690 23474 704
rect 22944 684 22947 690
rect 23468 688 23474 690
rect 23491 688 23497 705
rect 23468 685 23497 688
rect 23697 684 23700 710
rect 23726 704 23729 710
rect 23726 690 23996 704
rect 23726 684 23729 690
rect 21444 671 21473 674
rect 21444 670 21450 671
rect 20992 656 21450 670
rect 20892 651 20921 654
rect 21444 654 21450 656
rect 21467 654 21473 671
rect 21444 651 21473 654
rect 21535 650 21538 676
rect 21564 670 21567 676
rect 22180 671 22209 674
rect 22180 670 22186 671
rect 21564 656 22186 670
rect 21564 650 21567 656
rect 22180 654 22186 656
rect 22203 654 22209 671
rect 22594 671 22623 674
rect 22594 670 22600 671
rect 22180 651 22209 654
rect 22234 656 22600 670
rect 17332 622 17510 636
rect 17332 616 17335 622
rect 17671 616 17674 642
rect 17700 636 17703 642
rect 18132 637 18161 640
rect 18132 636 18138 637
rect 17700 622 18138 636
rect 17700 616 17703 622
rect 18132 620 18138 622
rect 18155 620 18161 637
rect 18132 617 18161 620
rect 18177 616 18180 642
rect 18206 636 18209 642
rect 18546 637 18575 640
rect 18546 636 18552 637
rect 18206 622 18552 636
rect 18206 616 18209 622
rect 18546 620 18552 622
rect 18569 620 18575 637
rect 18546 617 18575 620
rect 18683 616 18686 642
rect 18712 636 18715 642
rect 19006 637 19035 640
rect 19006 636 19012 637
rect 18712 622 19012 636
rect 18712 616 18715 622
rect 19006 620 19012 622
rect 19029 620 19035 637
rect 19006 617 19035 620
rect 19051 616 19054 642
rect 19080 636 19083 642
rect 19420 637 19449 640
rect 19420 636 19426 637
rect 19080 622 19426 636
rect 19080 616 19083 622
rect 19420 620 19426 622
rect 19443 620 19449 637
rect 19420 617 19449 620
rect 19603 616 19606 642
rect 19632 636 19635 642
rect 20064 637 20093 640
rect 20064 636 20070 637
rect 19632 622 20070 636
rect 19632 616 19635 622
rect 20064 620 20070 622
rect 20087 620 20093 637
rect 20478 637 20507 640
rect 20478 636 20484 637
rect 20064 617 20093 620
rect 20118 622 20484 636
rect 15216 588 15394 602
rect 15216 582 15219 588
rect 15417 582 15420 608
rect 15446 602 15449 608
rect 15464 603 15493 606
rect 15464 602 15470 603
rect 15446 588 15470 602
rect 15446 582 15449 588
rect 15464 586 15470 588
rect 15487 586 15493 603
rect 15464 583 15493 586
rect 15509 582 15512 608
rect 15538 602 15541 608
rect 15740 603 15769 606
rect 15740 602 15746 603
rect 15538 588 15746 602
rect 15538 582 15541 588
rect 15740 586 15746 588
rect 15763 586 15769 603
rect 15740 583 15769 586
rect 15785 582 15788 608
rect 15814 602 15817 608
rect 16154 603 16183 606
rect 16154 602 16160 603
rect 15814 588 16160 602
rect 15814 582 15817 588
rect 16154 586 16160 588
rect 16177 586 16183 603
rect 16154 583 16183 586
rect 16199 582 16202 608
rect 16228 602 16231 608
rect 16292 603 16321 606
rect 16292 602 16298 603
rect 16228 588 16298 602
rect 16228 582 16231 588
rect 16292 586 16298 588
rect 16315 586 16321 603
rect 16292 583 16321 586
rect 16337 582 16340 608
rect 16366 602 16369 608
rect 16706 603 16735 606
rect 16706 602 16712 603
rect 16366 588 16712 602
rect 16366 582 16369 588
rect 16706 586 16712 588
rect 16729 586 16735 603
rect 16706 583 16735 586
rect 16751 582 16754 608
rect 16780 602 16783 608
rect 17120 603 17149 606
rect 17120 602 17126 603
rect 16780 588 17126 602
rect 16780 582 16783 588
rect 17120 586 17126 588
rect 17143 586 17149 603
rect 17120 583 17149 586
rect 17165 582 17168 608
rect 17194 602 17197 608
rect 17580 603 17609 606
rect 17580 602 17586 603
rect 17194 588 17586 602
rect 17194 582 17197 588
rect 17580 586 17586 588
rect 17603 586 17609 603
rect 17855 602 17858 608
rect 17835 588 17858 602
rect 17580 583 17609 586
rect 17855 582 17858 588
rect 17884 582 17887 608
rect 17901 582 17904 608
rect 17930 602 17933 608
rect 17994 603 18023 606
rect 17994 602 18000 603
rect 17930 588 18000 602
rect 17930 582 17933 588
rect 17994 586 18000 588
rect 18017 586 18023 603
rect 17994 583 18023 586
rect 18039 582 18042 608
rect 18068 602 18071 608
rect 18408 603 18437 606
rect 18408 602 18414 603
rect 18068 588 18414 602
rect 18068 582 18071 588
rect 18408 586 18414 588
rect 18431 586 18437 603
rect 18408 583 18437 586
rect 18453 582 18456 608
rect 18482 602 18485 608
rect 18868 603 18897 606
rect 18868 602 18874 603
rect 18482 588 18874 602
rect 18482 582 18485 588
rect 18868 586 18874 588
rect 18891 586 18897 603
rect 18868 583 18897 586
rect 18913 582 18916 608
rect 18942 602 18945 608
rect 19282 603 19311 606
rect 19282 602 19288 603
rect 18942 588 19288 602
rect 18942 582 18945 588
rect 19282 586 19288 588
rect 19305 586 19311 603
rect 19282 583 19311 586
rect 19327 582 19330 608
rect 19356 602 19359 608
rect 19696 603 19725 606
rect 19696 602 19702 603
rect 19356 588 19702 602
rect 19356 582 19359 588
rect 19696 586 19702 588
rect 19719 586 19725 603
rect 19833 602 19836 608
rect 19813 588 19836 602
rect 19696 583 19725 586
rect 19833 582 19836 588
rect 19862 582 19865 608
rect 19879 582 19882 608
rect 19908 602 19911 608
rect 20118 602 20132 622
rect 20478 620 20484 622
rect 20501 620 20507 637
rect 20754 637 20783 640
rect 20754 636 20760 637
rect 20478 617 20507 620
rect 20532 622 20760 636
rect 19908 588 20132 602
rect 19908 582 19911 588
rect 20247 582 20250 608
rect 20276 602 20279 608
rect 20532 602 20546 622
rect 20754 620 20760 622
rect 20777 620 20783 637
rect 20754 617 20783 620
rect 21259 616 21262 642
rect 21288 636 21291 642
rect 21766 637 21795 640
rect 21766 636 21772 637
rect 21288 622 21772 636
rect 21288 616 21291 622
rect 21766 620 21772 622
rect 21789 620 21795 637
rect 21766 617 21795 620
rect 21811 616 21814 642
rect 21840 636 21843 642
rect 22234 636 22248 656
rect 22594 654 22600 656
rect 22617 654 22623 671
rect 22594 651 22623 654
rect 22639 650 22642 676
rect 22668 670 22671 676
rect 23192 671 23221 674
rect 23192 670 23198 671
rect 22668 656 23198 670
rect 22668 650 22671 656
rect 23192 654 23198 656
rect 23215 654 23221 671
rect 23192 651 23221 654
rect 23237 650 23240 676
rect 23266 670 23269 676
rect 23882 671 23911 674
rect 23882 670 23888 671
rect 23266 656 23888 670
rect 23266 650 23269 656
rect 23882 654 23888 656
rect 23905 654 23911 671
rect 23982 670 23996 690
rect 24433 684 24436 710
rect 24462 704 24465 710
rect 24462 690 24916 704
rect 24462 684 24465 690
rect 24296 671 24325 674
rect 24296 670 24302 671
rect 23982 656 24302 670
rect 23882 651 23911 654
rect 24296 654 24302 656
rect 24319 654 24325 671
rect 24296 651 24325 654
rect 24341 650 24344 676
rect 24370 670 24373 676
rect 24848 671 24877 674
rect 24848 670 24854 671
rect 24370 656 24854 670
rect 24370 650 24373 656
rect 24848 654 24854 656
rect 24871 654 24877 671
rect 24902 670 24916 690
rect 24939 684 24942 710
rect 24968 704 24971 710
rect 24968 690 25284 704
rect 24968 684 24971 690
rect 25170 671 25199 674
rect 25170 670 25176 671
rect 24902 656 25176 670
rect 24848 651 24877 654
rect 25170 654 25176 656
rect 25193 654 25199 671
rect 25270 670 25284 690
rect 25399 684 25402 710
rect 25428 704 25431 710
rect 26136 705 26165 708
rect 26136 704 26142 705
rect 25428 690 26142 704
rect 25428 684 25431 690
rect 26136 688 26142 690
rect 26159 688 26165 705
rect 26136 685 26165 688
rect 25584 671 25613 674
rect 25584 670 25590 671
rect 25270 656 25590 670
rect 25170 651 25199 654
rect 25584 654 25590 656
rect 25607 654 25613 671
rect 25584 651 25613 654
rect 25813 650 25816 676
rect 25842 670 25845 676
rect 26458 671 26487 674
rect 26458 670 26464 671
rect 25842 656 26464 670
rect 25842 650 25845 656
rect 26458 654 26464 656
rect 26481 654 26487 671
rect 26458 651 26487 654
rect 26503 650 26506 676
rect 26532 670 26535 676
rect 27010 671 27039 674
rect 27010 670 27016 671
rect 26532 656 27016 670
rect 26532 650 26535 656
rect 27010 654 27016 656
rect 27033 654 27039 671
rect 27010 651 27039 654
rect 27331 650 27334 676
rect 27360 670 27363 676
rect 27884 671 27913 674
rect 27884 670 27890 671
rect 27360 656 27890 670
rect 27360 650 27363 656
rect 27884 654 27890 656
rect 27907 654 27913 671
rect 27884 651 27913 654
rect 21840 622 22248 636
rect 21840 616 21843 622
rect 22363 616 22366 642
rect 22392 636 22395 642
rect 22916 637 22945 640
rect 22916 636 22922 637
rect 22392 622 22922 636
rect 22392 616 22395 622
rect 22916 620 22922 622
rect 22939 620 22945 637
rect 23330 637 23359 640
rect 23330 636 23336 637
rect 22916 617 22945 620
rect 22970 622 23336 636
rect 20615 602 20618 608
rect 20276 588 20546 602
rect 20595 588 20618 602
rect 20276 582 20279 588
rect 20615 582 20618 588
rect 20644 582 20647 608
rect 20661 582 20664 608
rect 20690 602 20693 608
rect 21030 603 21059 606
rect 21030 602 21036 603
rect 20690 588 21036 602
rect 20690 582 20693 588
rect 21030 586 21036 588
rect 21053 586 21059 603
rect 21305 602 21308 608
rect 21285 588 21308 602
rect 21030 583 21059 586
rect 21305 582 21308 588
rect 21334 582 21337 608
rect 21397 582 21400 608
rect 21426 602 21429 608
rect 21582 603 21611 606
rect 21582 602 21588 603
rect 21426 588 21588 602
rect 21426 582 21429 588
rect 21582 586 21588 588
rect 21605 586 21611 603
rect 21903 602 21906 608
rect 21883 588 21906 602
rect 21582 583 21611 586
rect 21903 582 21906 588
rect 21932 582 21935 608
rect 22041 602 22044 608
rect 22021 588 22044 602
rect 22041 582 22044 588
rect 22070 582 22073 608
rect 22317 602 22320 608
rect 22297 588 22320 602
rect 22317 582 22320 588
rect 22346 582 22349 608
rect 22731 602 22734 608
rect 22711 588 22734 602
rect 22731 582 22734 588
rect 22760 582 22763 608
rect 22777 582 22780 608
rect 22806 602 22809 608
rect 22970 602 22984 622
rect 23330 620 23336 622
rect 23353 620 23359 637
rect 23606 637 23635 640
rect 23606 636 23612 637
rect 23330 617 23359 620
rect 23430 622 23612 636
rect 23053 602 23056 608
rect 22806 588 22984 602
rect 23033 588 23056 602
rect 22806 582 22809 588
rect 23053 582 23056 588
rect 23082 582 23085 608
rect 23099 582 23102 608
rect 23128 602 23131 608
rect 23430 602 23444 622
rect 23606 620 23612 622
rect 23629 620 23635 637
rect 23606 617 23635 620
rect 23651 616 23654 642
rect 23680 636 23683 642
rect 24158 637 24187 640
rect 24158 636 24164 637
rect 23680 622 24164 636
rect 23680 616 23683 622
rect 24158 620 24164 622
rect 24181 620 24187 637
rect 24158 617 24187 620
rect 24203 616 24206 642
rect 24232 636 24235 642
rect 24710 637 24739 640
rect 24710 636 24716 637
rect 24232 622 24716 636
rect 24232 616 24235 622
rect 24710 620 24716 622
rect 24733 620 24739 637
rect 24710 617 24739 620
rect 24755 616 24758 642
rect 24784 636 24787 642
rect 25308 637 25337 640
rect 25308 636 25314 637
rect 24784 622 25314 636
rect 24784 616 24787 622
rect 25308 620 25314 622
rect 25331 620 25337 637
rect 25308 617 25337 620
rect 25362 622 25560 636
rect 23128 588 23444 602
rect 23128 582 23131 588
rect 23467 582 23470 608
rect 23496 602 23499 608
rect 24020 603 24049 606
rect 24020 602 24026 603
rect 23496 588 24026 602
rect 23496 582 23499 588
rect 24020 586 24026 588
rect 24043 586 24049 603
rect 24020 583 24049 586
rect 24065 582 24068 608
rect 24094 602 24097 608
rect 24434 603 24463 606
rect 24434 602 24440 603
rect 24094 588 24440 602
rect 24094 582 24097 588
rect 24434 586 24440 588
rect 24457 586 24463 603
rect 24571 602 24574 608
rect 24551 588 24574 602
rect 24434 583 24463 586
rect 24571 582 24574 588
rect 24600 582 24603 608
rect 24985 602 24988 608
rect 24965 588 24988 602
rect 24985 582 24988 588
rect 25014 582 25017 608
rect 25031 582 25034 608
rect 25060 602 25063 608
rect 25362 602 25376 622
rect 25445 602 25448 608
rect 25060 588 25376 602
rect 25425 588 25448 602
rect 25060 582 25063 588
rect 25445 582 25448 588
rect 25474 582 25477 608
rect 25546 602 25560 622
rect 25675 616 25678 642
rect 25704 636 25707 642
rect 26274 637 26303 640
rect 26274 636 26280 637
rect 25704 622 26280 636
rect 25704 616 25707 622
rect 26274 620 26280 622
rect 26297 620 26303 637
rect 26274 617 26303 620
rect 26319 616 26322 642
rect 26348 636 26351 642
rect 26734 637 26763 640
rect 26734 636 26740 637
rect 26348 622 26740 636
rect 26348 616 26351 622
rect 26734 620 26740 622
rect 26757 620 26763 637
rect 27148 637 27177 640
rect 27148 636 27154 637
rect 26734 617 26763 620
rect 26788 622 27154 636
rect 25722 603 25751 606
rect 25722 602 25728 603
rect 25546 588 25728 602
rect 25722 586 25728 588
rect 25745 586 25751 603
rect 25859 602 25862 608
rect 25839 588 25862 602
rect 25722 583 25751 586
rect 25859 582 25862 588
rect 25888 582 25891 608
rect 25905 582 25908 608
rect 25934 602 25937 608
rect 25998 603 26027 606
rect 25998 602 26004 603
rect 25934 588 26004 602
rect 25934 582 25937 588
rect 25998 586 26004 588
rect 26021 586 26027 603
rect 25998 583 26027 586
rect 26181 582 26184 608
rect 26210 602 26213 608
rect 26596 603 26625 606
rect 26596 602 26602 603
rect 26210 588 26602 602
rect 26210 582 26213 588
rect 26596 586 26602 588
rect 26619 586 26625 603
rect 26596 583 26625 586
rect 26641 582 26644 608
rect 26670 602 26673 608
rect 26788 602 26802 622
rect 27148 620 27154 622
rect 27171 620 27177 637
rect 27424 637 27453 640
rect 27424 636 27430 637
rect 27148 617 27177 620
rect 27202 622 27430 636
rect 26871 602 26874 608
rect 26670 588 26802 602
rect 26851 588 26874 602
rect 26670 582 26673 588
rect 26871 582 26874 588
rect 26900 582 26903 608
rect 26917 582 26920 608
rect 26946 602 26949 608
rect 27202 602 27216 622
rect 27424 620 27430 622
rect 27447 620 27453 637
rect 27424 617 27453 620
rect 27469 616 27472 642
rect 27498 636 27501 642
rect 28022 637 28051 640
rect 28022 636 28028 637
rect 27498 622 28028 636
rect 27498 616 27501 622
rect 28022 620 28028 622
rect 28045 620 28051 637
rect 28022 617 28051 620
rect 27285 602 27288 608
rect 26946 588 27216 602
rect 27265 588 27288 602
rect 26946 582 26949 588
rect 27285 582 27288 588
rect 27314 582 27317 608
rect 27561 602 27564 608
rect 27541 588 27564 602
rect 27561 582 27564 588
rect 27590 582 27593 608
rect 27745 602 27748 608
rect 27725 588 27748 602
rect 27745 582 27748 588
rect 27774 582 27777 608
rect 28159 602 28162 608
rect 28139 588 28162 602
rect 28159 582 28162 588
rect 28188 582 28191 608
rect 644 557 34408 568
rect 644 531 6631 557
rect 6657 531 12631 557
rect 12657 531 18631 557
rect 18657 531 24631 557
rect 24657 531 30631 557
rect 30657 531 34408 557
rect 644 520 34408 531
rect 927 480 930 506
rect 956 500 959 506
rect 2077 500 2080 506
rect 956 486 2080 500
rect 956 480 959 486
rect 2077 480 2080 486
rect 2106 480 2109 506
rect 605 446 608 472
rect 634 466 637 472
rect 2859 466 2862 472
rect 634 452 2862 466
rect 634 446 637 452
rect 2859 446 2862 452
rect 2888 446 2891 472
rect 21121 446 21124 472
rect 21150 466 21153 472
rect 22041 466 22044 472
rect 21150 452 22044 466
rect 21150 446 21153 452
rect 22041 446 22044 452
rect 22070 446 22073 472
rect 26917 446 26920 472
rect 26946 466 26949 472
rect 27561 466 27564 472
rect 26946 452 27564 466
rect 26946 446 26949 452
rect 27561 446 27564 452
rect 27590 446 27593 472
rect 7 412 10 438
rect 36 432 39 438
rect 1387 432 1390 438
rect 36 418 1390 432
rect 36 412 39 418
rect 1387 412 1390 418
rect 1416 412 1419 438
rect 20983 412 20986 438
rect 21012 432 21015 438
rect 21903 432 21906 438
rect 21012 418 21906 432
rect 21012 412 21015 418
rect 21903 412 21906 418
rect 21932 412 21935 438
rect 26641 412 26644 438
rect 26670 432 26673 438
rect 27285 432 27288 438
rect 26670 418 27288 432
rect 26670 412 26673 418
rect 27285 412 27288 418
rect 27314 412 27317 438
rect 145 378 148 404
rect 174 398 177 404
rect 1663 398 1666 404
rect 174 384 1666 398
rect 174 378 177 384
rect 1663 378 1666 384
rect 1692 378 1695 404
rect 14635 378 14638 404
rect 14664 398 14667 404
rect 15417 398 15420 404
rect 14664 384 15420 398
rect 14664 378 14667 384
rect 15417 378 15420 384
rect 15446 378 15449 404
rect 17395 378 17398 404
rect 17424 398 17427 404
rect 17855 398 17858 404
rect 17424 384 17858 398
rect 17424 378 17427 384
rect 17855 378 17858 384
rect 17884 378 17887 404
rect 20569 378 20572 404
rect 20598 398 20601 404
rect 21305 398 21308 404
rect 20598 384 21308 398
rect 20598 378 20601 384
rect 21305 378 21308 384
rect 21334 378 21337 404
rect 22087 378 22090 404
rect 22116 398 22119 404
rect 23053 398 23056 404
rect 22116 384 23056 398
rect 22116 378 22119 384
rect 23053 378 23056 384
rect 23082 378 23085 404
rect 24295 378 24298 404
rect 24324 398 24327 404
rect 24985 398 24988 404
rect 24324 384 24988 398
rect 24324 378 24327 384
rect 24985 378 24988 384
rect 25014 378 25017 404
rect 25261 378 25264 404
rect 25290 398 25293 404
rect 25905 398 25908 404
rect 25290 384 25908 398
rect 25290 378 25293 384
rect 25905 378 25908 384
rect 25934 378 25937 404
rect 27193 378 27196 404
rect 27222 398 27225 404
rect 28159 398 28162 404
rect 27222 384 28162 398
rect 27222 378 27225 384
rect 28159 378 28162 384
rect 28188 378 28191 404
rect 1387 344 1390 370
rect 1416 364 1419 370
rect 2537 364 2540 370
rect 1416 350 2540 364
rect 1416 344 1419 350
rect 2537 344 2540 350
rect 2566 344 2569 370
rect 6217 344 6220 370
rect 6246 364 6249 370
rect 6447 364 6450 370
rect 6246 350 6450 364
rect 6246 344 6249 350
rect 6447 344 6450 350
rect 6476 344 6479 370
rect 7735 344 7738 370
rect 7764 364 7767 370
rect 8011 364 8014 370
rect 7764 350 8014 364
rect 7764 344 7767 350
rect 8011 344 8014 350
rect 8040 344 8043 370
rect 9391 344 9394 370
rect 9420 364 9423 370
rect 10127 364 10130 370
rect 9420 350 10130 364
rect 9420 344 9423 350
rect 10127 344 10130 350
rect 10156 344 10159 370
rect 12703 344 12706 370
rect 12732 364 12735 370
rect 13071 364 13074 370
rect 12732 350 13074 364
rect 12732 344 12735 350
rect 13071 344 13074 350
rect 13100 344 13103 370
rect 13531 344 13534 370
rect 13560 364 13563 370
rect 14313 364 14316 370
rect 13560 350 14316 364
rect 13560 344 13563 350
rect 14313 344 14316 350
rect 14342 344 14345 370
rect 15049 344 15052 370
rect 15078 364 15081 370
rect 15509 364 15512 370
rect 15078 350 15512 364
rect 15078 344 15081 350
rect 15509 344 15512 350
rect 15538 344 15541 370
rect 15739 344 15742 370
rect 15768 364 15771 370
rect 16199 364 16202 370
rect 15768 350 16202 364
rect 15768 344 15771 350
rect 16199 344 16202 350
rect 16228 344 16231 370
rect 17533 344 17536 370
rect 17562 364 17565 370
rect 17901 364 17904 370
rect 17562 350 17904 364
rect 17562 344 17565 350
rect 17901 344 17904 350
rect 17930 344 17933 370
rect 19327 344 19330 370
rect 19356 364 19359 370
rect 19833 364 19836 370
rect 19356 350 19836 364
rect 19356 344 19359 350
rect 19833 344 19836 350
rect 19862 344 19865 370
rect 20017 344 20020 370
rect 20046 364 20049 370
rect 20615 364 20618 370
rect 20046 350 20618 364
rect 20046 344 20049 350
rect 20615 344 20618 350
rect 20644 344 20647 370
rect 20845 344 20848 370
rect 20874 364 20877 370
rect 21397 364 21400 370
rect 20874 350 21400 364
rect 20874 344 20877 350
rect 21397 344 21400 350
rect 21426 344 21429 370
rect 21949 344 21952 370
rect 21978 364 21981 370
rect 22731 364 22734 370
rect 21978 350 22734 364
rect 21978 344 21981 350
rect 22731 344 22734 350
rect 22760 344 22763 370
rect 23881 344 23884 370
rect 23910 364 23913 370
rect 24571 364 24574 370
rect 23910 350 24574 364
rect 23910 344 23913 350
rect 24571 344 24574 350
rect 24600 344 24603 370
rect 25123 344 25126 370
rect 25152 364 25155 370
rect 25859 364 25862 370
rect 25152 350 25862 364
rect 25152 344 25155 350
rect 25859 344 25862 350
rect 25888 344 25891 370
rect 27055 344 27058 370
rect 27084 364 27087 370
rect 27745 364 27748 370
rect 27084 350 27748 364
rect 27084 344 27087 350
rect 27745 344 27748 350
rect 27774 344 27777 370
rect 881 310 884 336
rect 910 330 913 336
rect 2583 330 2586 336
rect 910 316 2586 330
rect 910 310 913 316
rect 2583 310 2586 316
rect 2612 310 2615 336
rect 21443 310 21446 336
rect 21472 330 21475 336
rect 22317 330 22320 336
rect 21472 316 22320 330
rect 21472 310 21475 316
rect 22317 310 22320 316
rect 22346 310 22349 336
rect 24755 276 24758 302
rect 24784 296 24787 302
rect 25445 296 25448 302
rect 24784 282 25448 296
rect 24784 276 24787 282
rect 25445 276 25448 282
rect 25474 276 25477 302
rect 26273 276 26276 302
rect 26302 296 26305 302
rect 26871 296 26874 302
rect 26302 282 26874 296
rect 26302 276 26305 282
rect 26871 276 26874 282
rect 26900 276 26903 302
<< via1 >>
rect 332 1704 358 1730
rect 3414 1704 3440 1730
rect 838 1670 864 1696
rect 2954 1670 2980 1696
rect 12430 1670 12456 1696
rect 12936 1670 12962 1696
rect 6631 1619 6657 1645
rect 12631 1619 12657 1645
rect 18631 1619 18657 1645
rect 24631 1619 24657 1645
rect 30631 1619 30657 1645
rect 700 1568 726 1594
rect 1666 1568 1692 1594
rect 1804 1568 1830 1594
rect 2034 1568 2060 1594
rect 2494 1568 2520 1594
rect 2632 1568 2658 1594
rect 2770 1568 2796 1594
rect 2908 1568 2934 1594
rect 3184 1568 3210 1594
rect 3322 1568 3348 1594
rect 3460 1568 3486 1594
rect 3690 1589 3716 1594
rect 3690 1572 3694 1589
rect 3694 1572 3711 1589
rect 3711 1572 3716 1589
rect 3690 1568 3716 1572
rect 3736 1568 3762 1594
rect 3874 1568 3900 1594
rect 4012 1568 4038 1594
rect 4150 1568 4176 1594
rect 4288 1568 4314 1594
rect 4426 1568 4452 1594
rect 4840 1589 4866 1594
rect 4840 1572 4844 1589
rect 4844 1572 4861 1589
rect 4861 1572 4866 1589
rect 4840 1568 4866 1572
rect 4886 1568 4912 1594
rect 5254 1568 5280 1594
rect 5530 1568 5556 1594
rect 5944 1568 5970 1594
rect 6220 1568 6246 1594
rect 6496 1568 6522 1594
rect 6726 1568 6752 1594
rect 6910 1589 6936 1594
rect 6910 1572 6914 1589
rect 6914 1572 6931 1589
rect 6931 1572 6936 1589
rect 6910 1568 6936 1572
rect 7048 1568 7074 1594
rect 7324 1568 7350 1594
rect 7646 1568 7672 1594
rect 8014 1568 8040 1594
rect 8474 1568 8500 1594
rect 8888 1568 8914 1594
rect 9302 1568 9328 1594
rect 9762 1568 9788 1594
rect 10222 1568 10248 1594
rect 10774 1568 10800 1594
rect 11326 1568 11352 1594
rect 11878 1568 11904 1594
rect 12568 1568 12594 1594
rect 13166 1568 13192 1594
rect 13810 1568 13836 1594
rect 14362 1568 14388 1594
rect 14914 1568 14940 1594
rect 15466 1568 15492 1594
rect 16018 1568 16044 1594
rect 16570 1568 16596 1594
rect 17030 1568 17056 1594
rect 17674 1568 17700 1594
rect 18364 1568 18390 1594
rect 18916 1568 18942 1594
rect 19468 1568 19494 1594
rect 20066 1568 20092 1594
rect 20618 1568 20644 1594
rect 2080 1534 2106 1560
rect 5116 1534 5142 1560
rect 148 1500 174 1526
rect 4564 1500 4590 1526
rect 8290 1534 8316 1560
rect 8612 1534 8638 1560
rect 9164 1534 9190 1560
rect 9578 1534 9604 1560
rect 10084 1534 10110 1560
rect 10636 1534 10662 1560
rect 11188 1534 11214 1560
rect 11740 1534 11766 1560
rect 12154 1534 12180 1560
rect 12982 1534 13008 1560
rect 13626 1534 13652 1560
rect 14500 1534 14526 1560
rect 15052 1534 15078 1560
rect 15880 1534 15906 1560
rect 16202 1534 16228 1560
rect 16754 1534 16780 1560
rect 17398 1534 17424 1560
rect 18226 1534 18252 1560
rect 18778 1534 18804 1560
rect 19330 1534 19356 1560
rect 19882 1534 19908 1560
rect 5530 1521 5556 1526
rect 5530 1504 5534 1521
rect 5534 1504 5551 1521
rect 5551 1504 5556 1521
rect 5530 1500 5556 1504
rect 5668 1500 5694 1526
rect 6220 1521 6246 1526
rect 6220 1504 6224 1521
rect 6224 1504 6241 1521
rect 6241 1504 6246 1521
rect 6220 1500 6246 1504
rect 6358 1500 6384 1526
rect 7186 1500 7212 1526
rect 7600 1500 7626 1526
rect 7784 1500 7810 1526
rect 8336 1500 8362 1526
rect 8750 1500 8776 1526
rect 9440 1500 9466 1526
rect 9946 1500 9972 1526
rect 10498 1500 10524 1526
rect 11050 1500 11076 1526
rect 11464 1500 11490 1526
rect 12016 1500 12042 1526
rect 12752 1500 12778 1526
rect 13304 1500 13330 1526
rect 13902 1500 13928 1526
rect 14638 1500 14664 1526
rect 15190 1500 15216 1526
rect 15926 1500 15952 1526
rect 16340 1500 16366 1526
rect 16892 1500 16918 1526
rect 17536 1500 17562 1526
rect 10 1466 36 1492
rect 2080 1487 2106 1492
rect 2080 1470 2084 1487
rect 2084 1470 2101 1487
rect 2101 1470 2106 1487
rect 2080 1466 2106 1470
rect 286 1432 312 1458
rect 4978 1466 5004 1492
rect 6956 1466 6982 1492
rect 7876 1466 7902 1492
rect 8980 1466 9006 1492
rect 9808 1466 9834 1492
rect 10360 1466 10386 1492
rect 11096 1466 11122 1492
rect 11786 1466 11812 1492
rect 12430 1466 12456 1492
rect 12936 1466 12962 1492
rect 12890 1432 12916 1458
rect 13442 1466 13468 1492
rect 14040 1466 14066 1492
rect 14086 1432 14112 1458
rect 14776 1466 14802 1492
rect 15328 1466 15354 1492
rect 16064 1466 16090 1492
rect 16616 1466 16642 1492
rect 17260 1466 17286 1492
rect 17306 1432 17332 1458
rect 17950 1466 17976 1492
rect 18502 1500 18528 1526
rect 19054 1500 19080 1526
rect 19606 1500 19632 1526
rect 20204 1500 20230 1526
rect 20848 1568 20874 1594
rect 21400 1568 21426 1594
rect 21768 1568 21794 1594
rect 22228 1568 22254 1594
rect 23746 1568 23772 1594
rect 24298 1568 24324 1594
rect 24436 1568 24462 1594
rect 24574 1568 24600 1594
rect 24712 1568 24738 1594
rect 24850 1568 24876 1594
rect 24988 1568 25014 1594
rect 25264 1568 25290 1594
rect 25540 1568 25566 1594
rect 25678 1568 25704 1594
rect 25954 1568 25980 1594
rect 26230 1568 26256 1594
rect 26368 1568 26394 1594
rect 26644 1568 26670 1594
rect 26920 1568 26946 1594
rect 27058 1568 27084 1594
rect 27334 1568 27360 1594
rect 27702 1568 27728 1594
rect 28024 1568 28050 1594
rect 28346 1568 28372 1594
rect 28760 1568 28786 1594
rect 29128 1568 29154 1594
rect 29542 1568 29568 1594
rect 29956 1568 29982 1594
rect 30370 1568 30396 1594
rect 30692 1568 30718 1594
rect 31060 1568 31086 1594
rect 31336 1568 31362 1594
rect 32164 1568 32190 1594
rect 32854 1568 32880 1594
rect 33268 1568 33294 1594
rect 33544 1589 33570 1594
rect 33544 1572 33548 1589
rect 33548 1572 33565 1589
rect 33565 1572 33570 1589
rect 33544 1568 33570 1572
rect 33728 1568 33754 1594
rect 33820 1589 33846 1594
rect 33820 1572 33824 1589
rect 33824 1572 33841 1589
rect 33841 1572 33846 1589
rect 33820 1568 33846 1572
rect 20986 1534 21012 1560
rect 21538 1534 21564 1560
rect 22366 1534 22392 1560
rect 25126 1534 25152 1560
rect 25816 1534 25842 1560
rect 26506 1534 26532 1560
rect 26966 1534 26992 1560
rect 27196 1534 27222 1560
rect 27472 1534 27498 1560
rect 28484 1534 28510 1560
rect 28990 1534 29016 1560
rect 29266 1534 29292 1560
rect 29680 1534 29706 1560
rect 30094 1534 30120 1560
rect 30508 1534 30534 1560
rect 31106 1534 31132 1560
rect 31474 1534 31500 1560
rect 32026 1534 32052 1560
rect 32624 1534 32650 1560
rect 21170 1500 21196 1526
rect 21814 1500 21840 1526
rect 22504 1500 22530 1526
rect 23884 1500 23910 1526
rect 25586 1500 25612 1526
rect 26276 1500 26302 1526
rect 27886 1500 27912 1526
rect 28300 1500 28326 1526
rect 28576 1500 28602 1526
rect 29036 1500 29062 1526
rect 29404 1500 29430 1526
rect 29818 1500 29844 1526
rect 30416 1500 30442 1526
rect 30784 1500 30810 1526
rect 31198 1500 31224 1526
rect 31796 1500 31822 1526
rect 32348 1500 32374 1526
rect 33958 1500 33984 1526
rect 17996 1432 18022 1458
rect 18686 1466 18712 1492
rect 19192 1466 19218 1492
rect 19744 1466 19770 1492
rect 20342 1466 20368 1492
rect 20434 1432 20460 1458
rect 21446 1466 21472 1492
rect 21952 1466 21978 1492
rect 27748 1466 27774 1492
rect 31750 1466 31776 1492
rect 31888 1432 31914 1458
rect 470 1398 496 1424
rect 2816 1398 2842 1424
rect 3631 1347 3657 1373
rect 9631 1347 9657 1373
rect 15631 1347 15657 1373
rect 21631 1347 21657 1373
rect 27631 1347 27657 1373
rect 33631 1347 33657 1373
rect 1482 1262 1508 1288
rect 976 1228 1002 1254
rect 1942 1228 1968 1254
rect 2218 1228 2244 1254
rect 3046 1228 3072 1254
rect 5806 1228 5832 1254
rect 14224 1228 14250 1254
rect 18088 1228 18114 1254
rect 20710 1228 20736 1254
rect 22090 1228 22116 1254
rect 22642 1249 22668 1254
rect 22642 1232 22646 1249
rect 22646 1232 22663 1249
rect 22663 1232 22668 1249
rect 22642 1228 22668 1232
rect 22780 1249 22806 1254
rect 22780 1232 22784 1249
rect 22784 1232 22801 1249
rect 22801 1232 22806 1249
rect 22918 1249 22944 1254
rect 22780 1228 22806 1232
rect 22918 1232 22922 1249
rect 22922 1232 22939 1249
rect 22939 1232 22944 1249
rect 22918 1228 22944 1232
rect 23056 1249 23082 1254
rect 23056 1232 23060 1249
rect 23060 1232 23077 1249
rect 23077 1232 23082 1249
rect 23056 1228 23082 1232
rect 23194 1249 23220 1254
rect 23194 1232 23198 1249
rect 23198 1232 23215 1249
rect 23215 1232 23220 1249
rect 23194 1228 23220 1232
rect 23332 1249 23358 1254
rect 23332 1232 23336 1249
rect 23336 1232 23353 1249
rect 23353 1232 23358 1249
rect 23332 1228 23358 1232
rect 23470 1249 23496 1254
rect 23470 1232 23474 1249
rect 23474 1232 23491 1249
rect 23491 1232 23496 1249
rect 23470 1228 23496 1232
rect 23608 1249 23634 1254
rect 23608 1232 23612 1249
rect 23612 1232 23629 1249
rect 23629 1232 23634 1249
rect 23608 1228 23634 1232
rect 24022 1249 24048 1254
rect 24022 1232 24026 1249
rect 24026 1232 24043 1249
rect 24043 1232 24048 1249
rect 24022 1228 24048 1232
rect 24160 1249 24186 1254
rect 24160 1232 24164 1249
rect 24164 1232 24181 1249
rect 24181 1232 24186 1249
rect 24160 1228 24186 1232
rect 32440 1228 32466 1254
rect 32716 1249 32742 1254
rect 32716 1232 32720 1249
rect 32720 1232 32737 1249
rect 32737 1232 32742 1249
rect 32716 1228 32742 1232
rect 32992 1249 33018 1254
rect 32992 1232 32996 1249
rect 32996 1232 33013 1249
rect 33013 1232 33018 1249
rect 32992 1228 33018 1232
rect 33130 1249 33156 1254
rect 33130 1232 33134 1249
rect 33134 1232 33151 1249
rect 33151 1232 33156 1249
rect 33130 1228 33156 1232
rect 33406 1228 33432 1254
rect 1252 1194 1278 1220
rect 1896 1194 1922 1220
rect 1114 1160 1140 1186
rect 1666 1160 1692 1186
rect 1850 1160 1876 1186
rect 424 1126 450 1152
rect 1390 1126 1416 1152
rect 1758 1126 1784 1152
rect 1804 1147 1830 1152
rect 1804 1130 1808 1147
rect 1808 1130 1825 1147
rect 1825 1130 1830 1147
rect 1988 1160 2014 1186
rect 2356 1194 2382 1220
rect 2908 1194 2934 1220
rect 1804 1126 1830 1130
rect 2862 1126 2888 1152
rect 6631 1075 6657 1101
rect 12631 1075 12657 1101
rect 18631 1075 18657 1101
rect 24631 1075 24657 1101
rect 30631 1075 30657 1101
rect 1482 1024 1508 1050
rect 1528 1024 1554 1050
rect 2126 1024 2152 1050
rect 2356 1024 2382 1050
rect 3414 1045 3440 1050
rect 3414 1028 3418 1045
rect 3418 1028 3435 1045
rect 3435 1028 3440 1045
rect 3414 1024 3440 1028
rect 1390 990 1416 1016
rect 2770 990 2796 1016
rect 562 956 588 982
rect 700 888 726 914
rect 1436 956 1462 982
rect 2678 956 2704 982
rect 22504 956 22530 982
rect 1528 943 1554 948
rect 1528 926 1532 943
rect 1532 926 1549 943
rect 1549 926 1554 943
rect 1528 922 1554 926
rect 1666 943 1692 948
rect 1666 926 1670 943
rect 1670 926 1687 943
rect 1687 926 1692 943
rect 1666 922 1692 926
rect 1758 922 1784 948
rect 1482 888 1508 914
rect 2586 922 2612 948
rect 2954 922 2980 948
rect 3460 922 3486 948
rect 4702 922 4728 948
rect 5806 922 5832 948
rect 6772 922 6798 948
rect 8060 922 8086 948
rect 9808 922 9834 948
rect 10774 922 10800 948
rect 12154 922 12180 948
rect 14224 922 14250 948
rect 15328 922 15354 948
rect 15880 922 15906 948
rect 21722 922 21748 948
rect 22228 922 22254 948
rect 25540 922 25566 948
rect 1942 854 1968 880
rect 3631 803 3657 829
rect 9631 803 9657 829
rect 15631 803 15657 829
rect 21631 803 21657 829
rect 27631 803 27657 829
rect 33631 803 33657 829
rect 1114 684 1140 710
rect 1206 650 1232 676
rect 1574 684 1600 710
rect 1804 684 1830 710
rect 13258 684 13284 710
rect 13948 684 13974 710
rect 1896 650 1922 676
rect 2494 650 2520 676
rect 2816 650 2842 676
rect 3322 650 3348 676
rect 3736 650 3762 676
rect 4840 650 4866 676
rect 5668 650 5694 676
rect 6496 650 6522 676
rect 6910 650 6936 676
rect 7876 650 7902 676
rect 8428 650 8454 676
rect 8842 650 8868 676
rect 9716 650 9742 676
rect 10084 650 10110 676
rect 10498 650 10524 676
rect 11188 650 11214 676
rect 11740 650 11766 676
rect 12430 650 12456 676
rect 12982 650 13008 676
rect 13672 650 13698 676
rect 19468 684 19494 710
rect 20710 684 20736 710
rect 14776 650 14802 676
rect 15466 650 15492 676
rect 16156 650 16182 676
rect 16616 650 16642 676
rect 17030 650 17056 676
rect 976 616 1002 642
rect 930 603 956 608
rect 930 586 934 603
rect 934 586 951 603
rect 951 586 956 603
rect 930 582 956 586
rect 1620 616 1646 642
rect 1758 616 1784 642
rect 2264 616 2290 642
rect 3092 616 3118 642
rect 3874 616 3900 642
rect 4150 616 4176 642
rect 4426 616 4452 642
rect 5116 616 5142 642
rect 5392 616 5418 642
rect 5944 616 5970 642
rect 6404 616 6430 642
rect 7048 616 7074 642
rect 7370 616 7396 642
rect 7646 616 7672 642
rect 1390 603 1416 608
rect 1390 586 1394 603
rect 1394 586 1411 603
rect 1411 586 1416 603
rect 1666 603 1692 608
rect 1390 582 1416 586
rect 1666 586 1670 603
rect 1670 586 1687 603
rect 1687 586 1692 603
rect 1666 582 1692 586
rect 1712 582 1738 608
rect 1850 582 1876 608
rect 2126 582 2152 608
rect 2540 582 2566 608
rect 3184 582 3210 608
rect 3690 582 3716 608
rect 4012 582 4038 608
rect 4288 582 4314 608
rect 4610 582 4636 608
rect 4978 582 5004 608
rect 5254 582 5280 608
rect 5530 582 5556 608
rect 6082 582 6108 608
rect 6450 582 6476 608
rect 6726 582 6752 608
rect 7186 582 7212 608
rect 7508 582 7534 608
rect 8290 616 8316 642
rect 8704 616 8730 642
rect 8014 603 8040 608
rect 8014 586 8018 603
rect 8018 586 8035 603
rect 8035 586 8040 603
rect 8014 582 8040 586
rect 8198 582 8224 608
rect 8566 582 8592 608
rect 8980 616 9006 642
rect 9532 616 9558 642
rect 9946 616 9972 642
rect 10360 616 10386 642
rect 10912 616 10938 642
rect 11326 616 11352 642
rect 9118 582 9144 608
rect 9486 582 9512 608
rect 10130 603 10156 608
rect 10130 586 10134 603
rect 10134 586 10151 603
rect 10151 586 10156 603
rect 10130 582 10156 586
rect 10314 582 10340 608
rect 10636 582 10662 608
rect 11050 582 11076 608
rect 11464 616 11490 642
rect 11878 616 11904 642
rect 12338 616 12364 642
rect 12844 616 12870 642
rect 13396 616 13422 642
rect 13810 616 13836 642
rect 11694 582 11720 608
rect 12016 582 12042 608
rect 12568 582 12594 608
rect 13074 603 13100 608
rect 13074 586 13078 603
rect 13078 586 13095 603
rect 13095 586 13100 603
rect 13074 582 13100 586
rect 13120 582 13146 608
rect 14086 616 14112 642
rect 14500 616 14526 642
rect 14960 616 14986 642
rect 14316 603 14342 608
rect 14316 586 14320 603
rect 14320 586 14337 603
rect 14337 586 14342 603
rect 14316 582 14342 586
rect 14362 582 14388 608
rect 15190 582 15216 608
rect 16018 616 16044 642
rect 16478 616 16504 642
rect 16892 616 16918 642
rect 17306 616 17332 642
rect 17812 650 17838 676
rect 18318 650 18344 676
rect 18778 650 18804 676
rect 19192 650 19218 676
rect 19744 650 19770 676
rect 20388 650 20414 676
rect 22918 684 22944 710
rect 23700 684 23726 710
rect 21538 650 21564 676
rect 17674 616 17700 642
rect 18180 616 18206 642
rect 18686 616 18712 642
rect 19054 616 19080 642
rect 19606 616 19632 642
rect 15420 582 15446 608
rect 15512 582 15538 608
rect 15788 582 15814 608
rect 16202 582 16228 608
rect 16340 582 16366 608
rect 16754 582 16780 608
rect 17168 582 17194 608
rect 17858 603 17884 608
rect 17858 586 17862 603
rect 17862 586 17879 603
rect 17879 586 17884 603
rect 17858 582 17884 586
rect 17904 582 17930 608
rect 18042 582 18068 608
rect 18456 582 18482 608
rect 18916 582 18942 608
rect 19330 582 19356 608
rect 19836 603 19862 608
rect 19836 586 19840 603
rect 19840 586 19857 603
rect 19857 586 19862 603
rect 19836 582 19862 586
rect 19882 582 19908 608
rect 20250 582 20276 608
rect 21262 616 21288 642
rect 21814 616 21840 642
rect 22642 650 22668 676
rect 23240 650 23266 676
rect 24436 684 24462 710
rect 24344 650 24370 676
rect 24942 684 24968 710
rect 25402 684 25428 710
rect 25816 650 25842 676
rect 26506 650 26532 676
rect 27334 650 27360 676
rect 22366 616 22392 642
rect 20618 603 20644 608
rect 20618 586 20622 603
rect 20622 586 20639 603
rect 20639 586 20644 603
rect 20618 582 20644 586
rect 20664 582 20690 608
rect 21308 603 21334 608
rect 21308 586 21312 603
rect 21312 586 21329 603
rect 21329 586 21334 603
rect 21308 582 21334 586
rect 21400 582 21426 608
rect 21906 603 21932 608
rect 21906 586 21910 603
rect 21910 586 21927 603
rect 21927 586 21932 603
rect 21906 582 21932 586
rect 22044 603 22070 608
rect 22044 586 22048 603
rect 22048 586 22065 603
rect 22065 586 22070 603
rect 22044 582 22070 586
rect 22320 603 22346 608
rect 22320 586 22324 603
rect 22324 586 22341 603
rect 22341 586 22346 603
rect 22320 582 22346 586
rect 22734 603 22760 608
rect 22734 586 22738 603
rect 22738 586 22755 603
rect 22755 586 22760 603
rect 22734 582 22760 586
rect 22780 582 22806 608
rect 23056 603 23082 608
rect 23056 586 23060 603
rect 23060 586 23077 603
rect 23077 586 23082 603
rect 23056 582 23082 586
rect 23102 582 23128 608
rect 23654 616 23680 642
rect 24206 616 24232 642
rect 24758 616 24784 642
rect 23470 582 23496 608
rect 24068 582 24094 608
rect 24574 603 24600 608
rect 24574 586 24578 603
rect 24578 586 24595 603
rect 24595 586 24600 603
rect 24574 582 24600 586
rect 24988 603 25014 608
rect 24988 586 24992 603
rect 24992 586 25009 603
rect 25009 586 25014 603
rect 24988 582 25014 586
rect 25034 582 25060 608
rect 25448 603 25474 608
rect 25448 586 25452 603
rect 25452 586 25469 603
rect 25469 586 25474 603
rect 25448 582 25474 586
rect 25678 616 25704 642
rect 26322 616 26348 642
rect 25862 603 25888 608
rect 25862 586 25866 603
rect 25866 586 25883 603
rect 25883 586 25888 603
rect 25862 582 25888 586
rect 25908 582 25934 608
rect 26184 582 26210 608
rect 26644 582 26670 608
rect 26874 603 26900 608
rect 26874 586 26878 603
rect 26878 586 26895 603
rect 26895 586 26900 603
rect 26874 582 26900 586
rect 26920 582 26946 608
rect 27472 616 27498 642
rect 27288 603 27314 608
rect 27288 586 27292 603
rect 27292 586 27309 603
rect 27309 586 27314 603
rect 27288 582 27314 586
rect 27564 603 27590 608
rect 27564 586 27568 603
rect 27568 586 27585 603
rect 27585 586 27590 603
rect 27564 582 27590 586
rect 27748 603 27774 608
rect 27748 586 27752 603
rect 27752 586 27769 603
rect 27769 586 27774 603
rect 27748 582 27774 586
rect 28162 603 28188 608
rect 28162 586 28166 603
rect 28166 586 28183 603
rect 28183 586 28188 603
rect 28162 582 28188 586
rect 6631 531 6657 557
rect 12631 531 12657 557
rect 18631 531 18657 557
rect 24631 531 24657 557
rect 30631 531 30657 557
rect 930 480 956 506
rect 2080 480 2106 506
rect 608 446 634 472
rect 2862 446 2888 472
rect 21124 446 21150 472
rect 22044 446 22070 472
rect 26920 446 26946 472
rect 27564 446 27590 472
rect 10 412 36 438
rect 1390 412 1416 438
rect 20986 412 21012 438
rect 21906 412 21932 438
rect 26644 412 26670 438
rect 27288 412 27314 438
rect 148 378 174 404
rect 1666 378 1692 404
rect 14638 378 14664 404
rect 15420 378 15446 404
rect 17398 378 17424 404
rect 17858 378 17884 404
rect 20572 378 20598 404
rect 21308 378 21334 404
rect 22090 378 22116 404
rect 23056 378 23082 404
rect 24298 378 24324 404
rect 24988 378 25014 404
rect 25264 378 25290 404
rect 25908 378 25934 404
rect 27196 378 27222 404
rect 28162 378 28188 404
rect 1390 344 1416 370
rect 2540 344 2566 370
rect 6220 344 6246 370
rect 6450 344 6476 370
rect 7738 344 7764 370
rect 8014 344 8040 370
rect 9394 344 9420 370
rect 10130 344 10156 370
rect 12706 344 12732 370
rect 13074 344 13100 370
rect 13534 344 13560 370
rect 14316 344 14342 370
rect 15052 344 15078 370
rect 15512 344 15538 370
rect 15742 344 15768 370
rect 16202 344 16228 370
rect 17536 344 17562 370
rect 17904 344 17930 370
rect 19330 344 19356 370
rect 19836 344 19862 370
rect 20020 344 20046 370
rect 20618 344 20644 370
rect 20848 344 20874 370
rect 21400 344 21426 370
rect 21952 344 21978 370
rect 22734 344 22760 370
rect 23884 344 23910 370
rect 24574 344 24600 370
rect 25126 344 25152 370
rect 25862 344 25888 370
rect 27058 344 27084 370
rect 27748 344 27774 370
rect 884 310 910 336
rect 2586 310 2612 336
rect 21446 310 21472 336
rect 22320 310 22346 336
rect 24758 276 24784 302
rect 25448 276 25474 302
rect 26276 276 26302 302
rect 26874 276 26900 302
<< metal2 >>
rect 9 1900 37 2200
rect 147 1900 175 2200
rect 285 1900 313 2200
rect 423 1900 451 2200
rect 561 1900 589 2200
rect 699 1900 727 2200
rect 837 1900 865 2200
rect 975 1900 1003 2200
rect 1113 1900 1141 2200
rect 1251 1900 1279 2200
rect 1389 1900 1417 2200
rect 1527 1900 1555 2200
rect 1665 1900 1693 2200
rect 1803 1900 1831 2200
rect 1941 1900 1969 2200
rect 2079 1900 2107 2200
rect 2217 1900 2245 2200
rect 2355 1900 2383 2200
rect 2493 1900 2521 2200
rect 2631 1900 2659 2200
rect 2769 1900 2797 2200
rect 2907 1900 2935 2200
rect 3045 1900 3073 2200
rect 3183 1900 3211 2200
rect 3321 1900 3349 2200
rect 3459 1900 3487 2200
rect 3597 1900 3625 2200
rect 3735 1900 3763 2200
rect 3873 1900 3901 2200
rect 4011 1900 4039 2200
rect 4149 1900 4177 2200
rect 4287 1900 4315 2200
rect 4425 1900 4453 2200
rect 4563 1900 4591 2200
rect 4701 1900 4729 2200
rect 4839 1900 4867 2200
rect 4977 1900 5005 2200
rect 5115 1900 5143 2200
rect 5253 1900 5281 2200
rect 5391 1900 5419 2200
rect 5529 1900 5557 2200
rect 5667 1900 5695 2200
rect 5805 1900 5833 2200
rect 5943 1900 5971 2200
rect 6081 1900 6109 2200
rect 6219 1900 6247 2200
rect 6357 1900 6385 2200
rect 6495 1900 6523 2200
rect 6633 1900 6661 2200
rect 6771 1900 6799 2200
rect 6909 1900 6937 2200
rect 7047 1900 7075 2200
rect 7185 1900 7213 2200
rect 7323 1900 7351 2200
rect 7461 1900 7489 2200
rect 7599 1900 7627 2200
rect 7737 1900 7765 2200
rect 7875 1900 7903 2200
rect 8013 1900 8041 2200
rect 8151 1900 8179 2200
rect 8289 1900 8317 2200
rect 8427 1900 8455 2200
rect 8565 1900 8593 2200
rect 8703 1900 8731 2200
rect 8841 1900 8869 2200
rect 8979 1900 9007 2200
rect 9117 1900 9145 2200
rect 9255 1900 9283 2200
rect 9393 1900 9421 2200
rect 9531 1900 9559 2200
rect 9669 1900 9697 2200
rect 9807 1900 9835 2200
rect 9945 1900 9973 2200
rect 10083 1900 10111 2200
rect 10221 1900 10249 2200
rect 10359 1900 10387 2200
rect 10497 1900 10525 2200
rect 10635 1900 10663 2200
rect 10773 1900 10801 2200
rect 10911 1900 10939 2200
rect 11049 1900 11077 2200
rect 11187 1900 11215 2200
rect 11325 1900 11353 2200
rect 11463 1900 11491 2200
rect 11601 1900 11629 2200
rect 11739 1900 11767 2200
rect 11877 1900 11905 2200
rect 12015 1900 12043 2200
rect 12153 1900 12181 2200
rect 12291 1900 12319 2200
rect 12429 1900 12457 2200
rect 12567 1900 12595 2200
rect 12705 1900 12733 2200
rect 12843 1900 12871 2200
rect 12981 1900 13009 2200
rect 13119 1900 13147 2200
rect 13257 1900 13285 2200
rect 13395 1900 13423 2200
rect 13533 1900 13561 2200
rect 13671 1900 13699 2200
rect 13809 1900 13837 2200
rect 13947 1900 13975 2200
rect 14085 1900 14113 2200
rect 14223 1900 14251 2200
rect 14361 1900 14389 2200
rect 14499 1900 14527 2200
rect 14637 1900 14665 2200
rect 14775 1900 14803 2200
rect 14913 1900 14941 2200
rect 15051 1900 15079 2200
rect 15189 1900 15217 2200
rect 15327 1900 15355 2200
rect 15465 1900 15493 2200
rect 15603 1900 15631 2200
rect 15741 1900 15769 2200
rect 15879 1900 15907 2200
rect 16017 1900 16045 2200
rect 16155 1900 16183 2200
rect 16293 1900 16321 2200
rect 16431 1900 16459 2200
rect 16569 1900 16597 2200
rect 16707 1900 16735 2200
rect 16845 1900 16873 2200
rect 16983 1900 17011 2200
rect 17121 1900 17149 2200
rect 17259 1900 17287 2200
rect 17397 1900 17425 2200
rect 17535 1900 17563 2200
rect 17673 1900 17701 2200
rect 17811 1900 17839 2200
rect 17949 1900 17977 2200
rect 18087 1900 18115 2200
rect 18225 1900 18253 2200
rect 18363 1900 18391 2200
rect 18501 1900 18529 2200
rect 18639 1900 18667 2200
rect 18777 1900 18805 2200
rect 18915 1900 18943 2200
rect 19053 1900 19081 2200
rect 19191 1900 19219 2200
rect 19329 1900 19357 2200
rect 19467 1900 19495 2200
rect 19605 1900 19633 2200
rect 19743 1900 19771 2200
rect 19881 1900 19909 2200
rect 20019 1900 20047 2200
rect 20157 1900 20185 2200
rect 20295 1900 20323 2200
rect 20433 1900 20461 2200
rect 20571 1900 20599 2200
rect 20709 1900 20737 2200
rect 20847 1900 20875 2200
rect 20985 1900 21013 2200
rect 21123 1900 21151 2200
rect 21261 1900 21289 2200
rect 21399 1900 21427 2200
rect 21537 1900 21565 2200
rect 21675 1900 21703 2200
rect 21813 1900 21841 2200
rect 21951 1900 21979 2200
rect 22089 1900 22117 2200
rect 22227 1900 22255 2200
rect 22365 1900 22393 2200
rect 22503 1900 22531 2200
rect 22641 1900 22669 2200
rect 22779 1900 22807 2200
rect 22917 1900 22945 2200
rect 23055 1900 23083 2200
rect 23193 1900 23221 2200
rect 23331 1900 23359 2200
rect 23469 1900 23497 2200
rect 23607 1900 23635 2200
rect 23745 1900 23773 2200
rect 23883 1900 23911 2200
rect 24021 1900 24049 2200
rect 24159 1900 24187 2200
rect 24297 1900 24325 2200
rect 24435 1900 24463 2200
rect 24573 1900 24601 2200
rect 24711 1900 24739 2200
rect 24849 1900 24877 2200
rect 24987 1900 25015 2200
rect 25125 1900 25153 2200
rect 25263 1900 25291 2200
rect 25401 1900 25429 2200
rect 25539 1900 25567 2200
rect 25677 1900 25705 2200
rect 25815 1900 25843 2200
rect 25953 1900 25981 2200
rect 26091 1900 26119 2200
rect 26229 1900 26257 2200
rect 26367 1900 26395 2200
rect 26505 1900 26533 2200
rect 26643 1900 26671 2200
rect 26781 1900 26809 2200
rect 26919 1900 26947 2200
rect 27057 1900 27085 2200
rect 27195 1900 27223 2200
rect 27333 1900 27361 2200
rect 27471 1900 27499 2200
rect 27609 1900 27637 2200
rect 27747 1900 27775 2200
rect 27885 1900 27913 2200
rect 28023 1900 28051 2200
rect 28161 1900 28189 2200
rect 28299 1900 28327 2200
rect 28437 1900 28465 2200
rect 28575 1900 28603 2200
rect 28713 1900 28741 2200
rect 28851 1900 28879 2200
rect 28989 1900 29017 2200
rect 29127 1900 29155 2200
rect 29265 1900 29293 2200
rect 29403 1900 29431 2200
rect 29541 1900 29569 2200
rect 29679 1900 29707 2200
rect 29817 1900 29845 2200
rect 29955 1900 29983 2200
rect 30093 1900 30121 2200
rect 30231 1900 30259 2200
rect 30369 1900 30397 2200
rect 30507 1900 30535 2200
rect 30645 1900 30673 2200
rect 30783 1900 30811 2200
rect 30921 1900 30949 2200
rect 31059 1900 31087 2200
rect 31197 1900 31225 2200
rect 31335 1900 31363 2200
rect 31473 1900 31501 2200
rect 31611 1900 31639 2200
rect 31749 1900 31777 2200
rect 31887 1900 31915 2200
rect 32025 1900 32053 2200
rect 32163 1900 32191 2200
rect 32301 1900 32329 2200
rect 32439 1900 32467 2200
rect 32577 1900 32605 2200
rect 32715 1900 32743 2200
rect 32853 1900 32881 2200
rect 32991 1900 33019 2200
rect 33129 1900 33157 2200
rect 33267 1900 33295 2200
rect 33405 1900 33433 2200
rect 33543 1900 33571 2200
rect 33681 1900 33709 2200
rect 33819 1900 33847 2200
rect 33957 1900 33985 2200
rect 16 1495 30 1900
rect 154 1529 168 1900
rect 148 1526 174 1529
rect 148 1497 174 1500
rect 10 1492 36 1495
rect 10 1463 36 1466
rect 292 1461 306 1900
rect 332 1730 358 1733
rect 332 1701 358 1704
rect 286 1458 312 1461
rect 286 1429 312 1432
rect 338 517 352 1701
rect 430 1155 444 1900
rect 470 1424 496 1427
rect 470 1395 496 1398
rect 424 1152 450 1155
rect 424 1123 450 1126
rect 292 503 352 517
rect 10 438 36 441
rect 10 409 36 412
rect 16 300 30 409
rect 148 404 174 407
rect 148 375 174 378
rect 154 300 168 375
rect 292 300 306 503
rect 476 313 490 1395
rect 568 1061 582 1900
rect 706 1597 720 1900
rect 844 1741 858 1900
rect 844 1727 904 1741
rect 838 1696 864 1699
rect 838 1667 864 1670
rect 700 1594 726 1597
rect 700 1565 726 1568
rect 568 1047 628 1061
rect 562 982 588 985
rect 562 953 588 956
rect 430 300 490 313
rect 568 300 582 953
rect 614 475 628 1047
rect 700 914 726 917
rect 700 885 726 888
rect 608 472 634 475
rect 608 443 634 446
rect 706 300 720 885
rect 844 300 858 1667
rect 890 339 904 1727
rect 982 1257 996 1900
rect 976 1254 1002 1257
rect 976 1225 1002 1228
rect 1120 1189 1134 1900
rect 1258 1223 1272 1900
rect 1252 1220 1278 1223
rect 1252 1191 1278 1194
rect 1114 1186 1140 1189
rect 1114 1157 1140 1160
rect 1396 1155 1410 1900
rect 1481 1884 1509 1888
rect 1481 1851 1509 1856
rect 1488 1291 1502 1851
rect 1482 1288 1508 1291
rect 1482 1259 1508 1262
rect 1390 1152 1416 1155
rect 1390 1123 1416 1126
rect 1534 1053 1548 1900
rect 1672 1597 1686 1900
rect 1810 1597 1824 1900
rect 1849 1680 1877 1684
rect 1849 1647 1877 1652
rect 1666 1594 1692 1597
rect 1666 1565 1692 1568
rect 1804 1594 1830 1597
rect 1804 1565 1830 1568
rect 1856 1189 1870 1647
rect 1895 1544 1923 1548
rect 1895 1511 1923 1516
rect 1902 1223 1916 1511
rect 1948 1257 1962 1900
rect 2033 1884 2061 1888
rect 2033 1851 2061 1856
rect 1987 1816 2015 1820
rect 1987 1783 2015 1788
rect 1942 1254 1968 1257
rect 1942 1225 1968 1228
rect 1896 1220 1922 1223
rect 1896 1191 1922 1194
rect 1994 1189 2008 1783
rect 2040 1597 2054 1851
rect 2034 1594 2060 1597
rect 2034 1565 2060 1568
rect 2086 1563 2100 1900
rect 2080 1560 2106 1563
rect 2080 1531 2106 1534
rect 2080 1492 2106 1495
rect 2080 1463 2106 1466
rect 2033 1272 2061 1276
rect 2086 1265 2100 1463
rect 2125 1408 2153 1412
rect 2125 1375 2153 1380
rect 2061 1251 2100 1265
rect 2033 1239 2061 1244
rect 1666 1186 1692 1189
rect 1666 1157 1692 1160
rect 1850 1186 1876 1189
rect 1850 1157 1876 1160
rect 1988 1186 2014 1189
rect 1988 1157 2014 1160
rect 1482 1050 1508 1053
rect 1482 1021 1508 1024
rect 1528 1050 1554 1053
rect 1528 1021 1554 1024
rect 1390 1016 1416 1019
rect 1389 1000 1390 1004
rect 1416 1000 1417 1004
rect 1488 993 1502 1021
rect 1389 967 1417 972
rect 1436 982 1462 985
rect 1488 979 1594 993
rect 1436 953 1462 956
rect 1442 868 1456 953
rect 1528 948 1554 951
rect 1528 919 1554 922
rect 1482 914 1508 917
rect 1482 885 1508 888
rect 1435 864 1463 868
rect 1435 831 1463 836
rect 1488 732 1502 885
rect 1481 728 1509 732
rect 1114 710 1140 713
rect 1481 695 1509 700
rect 1114 681 1140 684
rect 976 642 1002 645
rect 976 613 1002 616
rect 930 608 956 611
rect 930 579 956 582
rect 936 509 950 579
rect 930 506 956 509
rect 930 477 956 480
rect 884 336 910 339
rect 884 307 910 310
rect 982 300 996 613
rect 1120 300 1134 681
rect 1206 676 1232 679
rect 1206 647 1232 650
rect 1212 313 1226 647
rect 1390 608 1416 611
rect 1390 579 1416 582
rect 1396 441 1410 579
rect 1390 438 1416 441
rect 1390 409 1416 412
rect 1390 370 1416 373
rect 1390 341 1416 344
rect 1212 300 1272 313
rect 1396 300 1410 341
rect 1534 300 1548 919
rect 1580 713 1594 979
rect 1672 951 1686 1157
rect 1758 1152 1784 1155
rect 1758 1123 1784 1126
rect 1804 1152 1830 1155
rect 1804 1123 1830 1126
rect 1764 951 1778 1123
rect 1810 1072 1824 1123
rect 1803 1068 1831 1072
rect 2132 1053 2146 1375
rect 2224 1257 2238 1900
rect 2218 1254 2244 1257
rect 2218 1225 2244 1228
rect 2362 1223 2376 1900
rect 2500 1597 2514 1900
rect 2638 1597 2652 1900
rect 2776 1597 2790 1900
rect 2914 1597 2928 1900
rect 2954 1696 2980 1699
rect 2954 1667 2980 1670
rect 2494 1594 2520 1597
rect 2494 1565 2520 1568
rect 2632 1594 2658 1597
rect 2632 1565 2658 1568
rect 2770 1594 2796 1597
rect 2770 1565 2796 1568
rect 2908 1594 2934 1597
rect 2908 1565 2934 1568
rect 2816 1424 2842 1427
rect 2816 1395 2842 1398
rect 2356 1220 2382 1223
rect 2356 1191 2382 1194
rect 1803 1035 1831 1040
rect 2126 1050 2152 1053
rect 2126 1021 2152 1024
rect 2356 1050 2382 1053
rect 2356 1021 2382 1024
rect 1666 948 1692 951
rect 1666 919 1692 922
rect 1758 948 1784 951
rect 1758 919 1784 922
rect 1942 880 1968 883
rect 1942 851 1968 854
rect 1574 710 1600 713
rect 1574 681 1600 684
rect 1804 710 1830 713
rect 1804 681 1830 684
rect 1620 642 1646 645
rect 1620 613 1646 616
rect 1758 642 1784 645
rect 1758 613 1784 616
rect 1626 313 1640 613
rect 1666 608 1692 611
rect 1666 579 1692 582
rect 1712 608 1738 611
rect 1712 579 1738 582
rect 1672 407 1686 579
rect 1666 404 1692 407
rect 1666 375 1692 378
rect 1718 324 1732 579
rect 1764 460 1778 613
rect 1757 456 1785 460
rect 1757 423 1785 428
rect 1711 320 1739 324
rect 1626 300 1686 313
rect 9 0 37 300
rect 147 0 175 300
rect 285 0 313 300
rect 423 299 490 300
rect 423 0 451 299
rect 561 0 589 300
rect 699 0 727 300
rect 837 0 865 300
rect 975 0 1003 300
rect 1113 0 1141 300
rect 1212 299 1279 300
rect 1251 0 1279 299
rect 1389 0 1417 300
rect 1527 0 1555 300
rect 1626 299 1693 300
rect 1665 0 1693 299
rect 1810 300 1824 681
rect 1896 676 1922 679
rect 1896 647 1922 650
rect 1850 608 1876 611
rect 1850 579 1876 582
rect 1856 528 1870 579
rect 1849 524 1877 528
rect 1849 491 1877 496
rect 1902 324 1916 647
rect 1895 320 1923 324
rect 1711 287 1739 292
rect 1803 0 1831 300
rect 1948 300 1962 851
rect 2264 642 2290 645
rect 2264 613 2290 616
rect 2126 608 2152 611
rect 2040 582 2126 585
rect 2040 579 2152 582
rect 2040 571 2146 579
rect 2040 324 2054 571
rect 2080 506 2106 509
rect 2080 477 2106 480
rect 2033 320 2061 324
rect 1895 287 1923 292
rect 1941 0 1969 300
rect 2086 300 2100 477
rect 2270 313 2284 613
rect 2224 300 2284 313
rect 2362 300 2376 1021
rect 2770 1016 2796 1019
rect 2770 987 2796 990
rect 2678 982 2704 985
rect 2678 953 2704 956
rect 2586 948 2612 951
rect 2586 919 2612 922
rect 2494 676 2520 679
rect 2494 647 2520 650
rect 2500 300 2514 647
rect 2540 608 2566 611
rect 2540 579 2566 582
rect 2546 373 2560 579
rect 2540 370 2566 373
rect 2540 341 2566 344
rect 2592 339 2606 919
rect 2684 517 2698 953
rect 2638 503 2698 517
rect 2586 336 2612 339
rect 2586 307 2612 310
rect 2638 300 2652 503
rect 2776 300 2790 987
rect 2822 679 2836 1395
rect 2908 1220 2934 1223
rect 2908 1191 2934 1194
rect 2862 1152 2888 1155
rect 2862 1123 2888 1126
rect 2816 676 2842 679
rect 2816 647 2842 650
rect 2868 475 2882 1123
rect 2862 472 2888 475
rect 2862 443 2888 446
rect 2914 300 2928 1191
rect 2960 951 2974 1667
rect 3052 1257 3066 1900
rect 3190 1597 3204 1900
rect 3328 1597 3342 1900
rect 3414 1730 3440 1733
rect 3414 1701 3440 1704
rect 3184 1594 3210 1597
rect 3184 1565 3210 1568
rect 3322 1594 3348 1597
rect 3322 1565 3348 1568
rect 3046 1254 3072 1257
rect 3046 1225 3072 1228
rect 3420 1053 3434 1701
rect 3466 1597 3480 1900
rect 3604 1724 3618 1900
rect 3604 1710 3710 1724
rect 3460 1594 3486 1597
rect 3460 1565 3486 1568
rect 3619 1373 3669 1656
rect 3696 1597 3710 1710
rect 3742 1597 3756 1900
rect 3880 1597 3894 1900
rect 4018 1597 4032 1900
rect 4156 1597 4170 1900
rect 4294 1597 4308 1900
rect 4432 1597 4446 1900
rect 3690 1594 3716 1597
rect 3690 1565 3716 1568
rect 3736 1594 3762 1597
rect 3736 1565 3762 1568
rect 3874 1594 3900 1597
rect 3874 1565 3900 1568
rect 4012 1594 4038 1597
rect 4012 1565 4038 1568
rect 4150 1594 4176 1597
rect 4150 1565 4176 1568
rect 4288 1594 4314 1597
rect 4288 1565 4314 1568
rect 4426 1594 4452 1597
rect 4426 1565 4452 1568
rect 4570 1529 4584 1900
rect 4708 1588 4722 1900
rect 4846 1673 4860 1900
rect 4846 1659 4906 1673
rect 4892 1597 4906 1659
rect 4840 1594 4866 1597
rect 4708 1574 4840 1588
rect 4840 1565 4866 1568
rect 4886 1594 4912 1597
rect 4886 1565 4912 1568
rect 4564 1526 4590 1529
rect 4564 1497 4590 1500
rect 4984 1495 4998 1900
rect 5122 1563 5136 1900
rect 5260 1597 5274 1900
rect 5254 1594 5280 1597
rect 5398 1588 5412 1900
rect 5536 1597 5550 1900
rect 5530 1594 5556 1597
rect 5398 1574 5504 1588
rect 5254 1565 5280 1568
rect 5116 1560 5142 1563
rect 5116 1531 5142 1534
rect 5490 1520 5504 1574
rect 5530 1565 5556 1568
rect 5674 1529 5688 1900
rect 5530 1526 5556 1529
rect 5490 1506 5530 1520
rect 5530 1497 5556 1500
rect 5668 1526 5694 1529
rect 5668 1497 5694 1500
rect 4978 1492 5004 1495
rect 4978 1463 5004 1466
rect 3619 1347 3631 1373
rect 3657 1347 3669 1373
rect 3414 1050 3440 1053
rect 3414 1021 3440 1024
rect 2954 948 2980 951
rect 2954 919 2980 922
rect 3460 948 3486 951
rect 3460 919 3486 922
rect 3322 676 3348 679
rect 3322 647 3348 650
rect 3092 642 3118 645
rect 3092 613 3118 616
rect 3098 313 3112 613
rect 3184 608 3210 611
rect 3184 579 3210 582
rect 3052 300 3112 313
rect 3190 300 3204 579
rect 3328 300 3342 647
rect 3466 300 3480 919
rect 3619 829 3669 1347
rect 5812 1257 5826 1900
rect 5950 1597 5964 1900
rect 5944 1594 5970 1597
rect 5944 1565 5970 1568
rect 6088 1520 6102 1900
rect 6226 1597 6240 1900
rect 6220 1594 6246 1597
rect 6220 1565 6246 1568
rect 6364 1529 6378 1900
rect 6502 1597 6516 1900
rect 6640 1724 6654 1900
rect 6640 1710 6746 1724
rect 6619 1645 6669 1656
rect 6619 1619 6631 1645
rect 6657 1619 6669 1645
rect 6496 1594 6522 1597
rect 6496 1565 6522 1568
rect 6220 1526 6246 1529
rect 6088 1506 6220 1520
rect 6220 1497 6246 1500
rect 6358 1526 6384 1529
rect 6358 1497 6384 1500
rect 5806 1254 5832 1257
rect 5806 1225 5832 1228
rect 6619 1174 6669 1619
rect 6732 1597 6746 1710
rect 6726 1594 6752 1597
rect 6778 1588 6792 1900
rect 6916 1673 6930 1900
rect 6916 1659 6976 1673
rect 6910 1594 6936 1597
rect 6778 1574 6910 1588
rect 6726 1565 6752 1568
rect 6910 1565 6936 1568
rect 6962 1495 6976 1659
rect 7054 1597 7068 1900
rect 7048 1594 7074 1597
rect 7048 1565 7074 1568
rect 7192 1529 7206 1900
rect 7330 1597 7344 1900
rect 7324 1594 7350 1597
rect 7324 1565 7350 1568
rect 7468 1537 7482 1900
rect 7606 1588 7620 1900
rect 7646 1594 7672 1597
rect 7606 1574 7646 1588
rect 7646 1565 7672 1568
rect 7468 1529 7620 1537
rect 7186 1526 7212 1529
rect 7468 1526 7626 1529
rect 7468 1523 7600 1526
rect 7186 1497 7212 1500
rect 7744 1520 7758 1900
rect 7784 1526 7810 1529
rect 7744 1506 7784 1520
rect 7600 1497 7626 1500
rect 7784 1497 7810 1500
rect 7882 1495 7896 1900
rect 8020 1597 8034 1900
rect 8014 1594 8040 1597
rect 8014 1565 8040 1568
rect 8158 1554 8172 1900
rect 8296 1605 8310 1900
rect 8296 1591 8356 1605
rect 8290 1560 8316 1563
rect 8158 1540 8290 1554
rect 8290 1531 8316 1534
rect 8342 1529 8356 1591
rect 8434 1588 8448 1900
rect 8474 1594 8500 1597
rect 8434 1574 8474 1588
rect 8474 1565 8500 1568
rect 8572 1554 8586 1900
rect 8612 1560 8638 1563
rect 8572 1540 8612 1554
rect 8612 1531 8638 1534
rect 8336 1526 8362 1529
rect 8710 1520 8724 1900
rect 8848 1588 8862 1900
rect 8888 1594 8914 1597
rect 8848 1574 8888 1588
rect 8888 1565 8914 1568
rect 8750 1526 8776 1529
rect 8710 1506 8750 1520
rect 8336 1497 8362 1500
rect 8750 1497 8776 1500
rect 8986 1495 9000 1900
rect 9124 1554 9138 1900
rect 9262 1588 9276 1900
rect 9302 1594 9328 1597
rect 9262 1574 9302 1588
rect 9302 1565 9328 1568
rect 9164 1560 9190 1563
rect 9124 1540 9164 1554
rect 9164 1531 9190 1534
rect 9400 1537 9414 1900
rect 9538 1554 9552 1900
rect 9676 1741 9690 1900
rect 9676 1727 9782 1741
rect 9578 1560 9604 1563
rect 9538 1540 9578 1554
rect 9400 1529 9460 1537
rect 9578 1531 9604 1534
rect 9400 1526 9466 1529
rect 9400 1523 9440 1526
rect 9440 1497 9466 1500
rect 6956 1492 6982 1495
rect 6956 1463 6982 1466
rect 7876 1492 7902 1495
rect 7876 1463 7902 1466
rect 8980 1492 9006 1495
rect 8980 1463 9006 1466
rect 6619 1146 6630 1174
rect 6658 1146 6669 1174
rect 6619 1101 6669 1146
rect 6619 1075 6631 1101
rect 6657 1075 6669 1101
rect 4702 948 4728 951
rect 4702 919 4728 922
rect 5806 948 5832 951
rect 5806 919 5832 922
rect 3619 803 3631 829
rect 3657 803 3669 829
rect 3619 634 3669 803
rect 3736 676 3762 679
rect 3736 647 3762 650
rect 3619 606 3630 634
rect 3658 606 3669 634
rect 3619 520 3669 606
rect 3690 608 3716 611
rect 3690 579 3716 582
rect 3696 313 3710 579
rect 3604 300 3710 313
rect 3742 300 3756 647
rect 3874 642 3900 645
rect 3874 613 3900 616
rect 4150 642 4176 645
rect 4150 613 4176 616
rect 4426 642 4452 645
rect 4426 613 4452 616
rect 3880 300 3894 613
rect 4012 608 4038 611
rect 4012 579 4038 582
rect 4018 300 4032 579
rect 4156 300 4170 613
rect 4288 608 4314 611
rect 4288 579 4314 582
rect 4294 300 4308 579
rect 4432 300 4446 613
rect 4610 608 4636 611
rect 4610 579 4636 582
rect 4616 313 4630 579
rect 4570 300 4630 313
rect 4708 300 4722 919
rect 4840 676 4866 679
rect 4840 647 4866 650
rect 5668 676 5694 679
rect 5668 647 5694 650
rect 4846 300 4860 647
rect 5116 642 5142 645
rect 5116 613 5142 616
rect 5392 642 5418 645
rect 5392 613 5418 616
rect 4978 608 5004 611
rect 4978 579 5004 582
rect 4984 300 4998 579
rect 5122 300 5136 613
rect 5254 608 5280 611
rect 5254 579 5280 582
rect 5260 300 5274 579
rect 5398 300 5412 613
rect 5530 608 5556 611
rect 5530 579 5556 582
rect 5536 300 5550 579
rect 5674 300 5688 647
rect 5812 300 5826 919
rect 6496 676 6522 679
rect 6496 647 6522 650
rect 5944 642 5970 645
rect 6404 642 6430 645
rect 5944 613 5970 616
rect 6364 622 6404 636
rect 5950 300 5964 613
rect 6082 608 6108 611
rect 6082 579 6108 582
rect 6088 300 6102 579
rect 6220 370 6246 373
rect 6220 341 6246 344
rect 6226 300 6240 341
rect 6364 300 6378 622
rect 6404 613 6430 616
rect 6450 608 6476 611
rect 6450 579 6476 582
rect 6456 373 6470 579
rect 6450 370 6476 373
rect 6450 341 6476 344
rect 6502 300 6516 647
rect 6619 557 6669 1075
rect 9619 1373 9669 1656
rect 9768 1597 9782 1727
rect 9762 1594 9788 1597
rect 9762 1565 9788 1568
rect 9814 1495 9828 1900
rect 9952 1529 9966 1900
rect 10090 1563 10104 1900
rect 10228 1597 10242 1900
rect 10222 1594 10248 1597
rect 10222 1565 10248 1568
rect 10084 1560 10110 1563
rect 10084 1531 10110 1534
rect 9946 1526 9972 1529
rect 9946 1497 9972 1500
rect 10366 1495 10380 1900
rect 10504 1529 10518 1900
rect 10642 1563 10656 1900
rect 10780 1597 10794 1900
rect 10774 1594 10800 1597
rect 10774 1565 10800 1568
rect 10636 1560 10662 1563
rect 10636 1531 10662 1534
rect 10918 1537 10932 1900
rect 11056 1588 11070 1900
rect 11056 1574 11116 1588
rect 10918 1529 11070 1537
rect 10498 1526 10524 1529
rect 10918 1526 11076 1529
rect 10918 1523 11050 1526
rect 10498 1497 10524 1500
rect 11050 1497 11076 1500
rect 11102 1495 11116 1574
rect 11194 1563 11208 1900
rect 11332 1597 11346 1900
rect 11326 1594 11352 1597
rect 11326 1565 11352 1568
rect 11188 1560 11214 1563
rect 11188 1531 11214 1534
rect 11470 1529 11484 1900
rect 11608 1588 11622 1900
rect 11746 1605 11760 1900
rect 11746 1591 11806 1605
rect 11884 1597 11898 1900
rect 11608 1574 11714 1588
rect 11700 1554 11714 1574
rect 11740 1560 11766 1563
rect 11700 1540 11740 1554
rect 11740 1531 11766 1534
rect 11464 1526 11490 1529
rect 11464 1497 11490 1500
rect 11792 1495 11806 1591
rect 11878 1594 11904 1597
rect 11878 1565 11904 1568
rect 12022 1529 12036 1900
rect 12160 1563 12174 1900
rect 12154 1560 12180 1563
rect 12154 1531 12180 1534
rect 12298 1537 12312 1900
rect 12436 1699 12450 1900
rect 12430 1696 12456 1699
rect 12430 1667 12456 1670
rect 12574 1597 12588 1900
rect 12619 1645 12669 1656
rect 12619 1619 12631 1645
rect 12657 1619 12669 1645
rect 12568 1594 12594 1597
rect 12568 1565 12594 1568
rect 12016 1526 12042 1529
rect 12298 1523 12450 1537
rect 12016 1497 12042 1500
rect 12436 1495 12450 1523
rect 9808 1492 9834 1495
rect 9808 1463 9834 1466
rect 10360 1492 10386 1495
rect 10360 1463 10386 1466
rect 11096 1492 11122 1495
rect 11096 1463 11122 1466
rect 11786 1492 11812 1495
rect 11786 1463 11812 1466
rect 12430 1492 12456 1495
rect 12430 1463 12456 1466
rect 9619 1347 9631 1373
rect 9657 1347 9669 1373
rect 6772 948 6798 951
rect 6772 919 6798 922
rect 8060 948 8086 951
rect 8060 919 8086 922
rect 6726 608 6752 611
rect 6726 579 6752 582
rect 6619 531 6631 557
rect 6657 531 6669 557
rect 6619 520 6669 531
rect 6732 313 6746 579
rect 6640 300 6746 313
rect 6778 300 6792 919
rect 6910 676 6936 679
rect 6910 647 6936 650
rect 7876 676 7902 679
rect 7876 647 7902 650
rect 6916 300 6930 647
rect 7048 642 7074 645
rect 7370 642 7396 645
rect 7048 613 7074 616
rect 7330 622 7370 636
rect 7054 300 7068 613
rect 7186 608 7212 611
rect 7186 579 7212 582
rect 7192 300 7206 579
rect 7330 300 7344 622
rect 7646 642 7672 645
rect 7370 613 7396 616
rect 7606 622 7646 636
rect 7508 608 7534 611
rect 7508 579 7534 582
rect 7514 313 7528 579
rect 7468 300 7528 313
rect 7606 300 7620 622
rect 7646 613 7672 616
rect 7738 370 7764 373
rect 7738 341 7764 344
rect 7744 300 7758 341
rect 7882 300 7896 647
rect 8014 608 8040 611
rect 8014 579 8040 582
rect 8020 373 8034 579
rect 8014 370 8040 373
rect 8014 341 8040 344
rect 8066 313 8080 919
rect 9619 829 9669 1347
rect 12619 1174 12669 1619
rect 12712 1520 12726 1900
rect 12752 1526 12778 1529
rect 12712 1506 12752 1520
rect 12752 1497 12778 1500
rect 12850 1469 12864 1900
rect 12936 1696 12962 1699
rect 12936 1667 12962 1670
rect 12942 1495 12956 1667
rect 12988 1563 13002 1900
rect 13126 1605 13140 1900
rect 13126 1597 13186 1605
rect 13126 1594 13192 1597
rect 13126 1591 13166 1594
rect 13166 1565 13192 1568
rect 12982 1560 13008 1563
rect 12982 1531 13008 1534
rect 13264 1537 13278 1900
rect 13264 1529 13324 1537
rect 13264 1526 13330 1529
rect 13264 1523 13304 1526
rect 13304 1497 13330 1500
rect 12936 1492 12962 1495
rect 12850 1461 12910 1469
rect 13402 1486 13416 1900
rect 13540 1605 13554 1900
rect 13678 1605 13692 1900
rect 13816 1673 13830 1900
rect 13816 1659 13922 1673
rect 13540 1591 13646 1605
rect 13678 1597 13830 1605
rect 13678 1594 13836 1597
rect 13678 1591 13810 1594
rect 13632 1563 13646 1591
rect 13810 1565 13836 1568
rect 13626 1560 13652 1563
rect 13626 1531 13652 1534
rect 13908 1529 13922 1659
rect 13902 1526 13928 1529
rect 13902 1497 13928 1500
rect 13442 1492 13468 1495
rect 13402 1472 13442 1486
rect 12936 1463 12962 1466
rect 13954 1486 13968 1900
rect 14040 1492 14066 1495
rect 13954 1472 14040 1486
rect 13442 1463 13468 1466
rect 14040 1463 14066 1466
rect 14092 1461 14106 1900
rect 12850 1458 12916 1461
rect 12850 1455 12890 1458
rect 12890 1429 12916 1432
rect 14086 1458 14112 1461
rect 14086 1429 14112 1432
rect 14230 1257 14244 1900
rect 14368 1597 14382 1900
rect 14362 1594 14388 1597
rect 14362 1565 14388 1568
rect 14506 1563 14520 1900
rect 14500 1560 14526 1563
rect 14500 1531 14526 1534
rect 14644 1529 14658 1900
rect 14638 1526 14664 1529
rect 14638 1497 14664 1500
rect 14782 1495 14796 1900
rect 14920 1597 14934 1900
rect 14914 1594 14940 1597
rect 14914 1565 14940 1568
rect 15058 1563 15072 1900
rect 15052 1560 15078 1563
rect 15052 1531 15078 1534
rect 15196 1529 15210 1900
rect 15190 1526 15216 1529
rect 15190 1497 15216 1500
rect 15334 1495 15348 1900
rect 15472 1597 15486 1900
rect 15610 1690 15624 1900
rect 15748 1741 15762 1900
rect 15886 1809 15900 1900
rect 16024 1877 16038 1900
rect 16024 1863 16084 1877
rect 15886 1795 16038 1809
rect 15748 1727 15946 1741
rect 15610 1676 15900 1690
rect 15466 1594 15492 1597
rect 15466 1565 15492 1568
rect 14776 1492 14802 1495
rect 14776 1463 14802 1466
rect 15328 1492 15354 1495
rect 15328 1463 15354 1466
rect 15619 1373 15669 1656
rect 15886 1563 15900 1676
rect 15880 1560 15906 1563
rect 15880 1531 15906 1534
rect 15932 1529 15946 1727
rect 16024 1597 16038 1795
rect 16018 1594 16044 1597
rect 16018 1565 16044 1568
rect 15926 1526 15952 1529
rect 15926 1497 15952 1500
rect 16070 1495 16084 1863
rect 16162 1554 16176 1900
rect 16202 1560 16228 1563
rect 16162 1540 16202 1554
rect 16202 1531 16228 1534
rect 16300 1537 16314 1900
rect 16438 1673 16452 1900
rect 16576 1741 16590 1900
rect 16576 1727 16636 1741
rect 16438 1659 16590 1673
rect 16576 1597 16590 1659
rect 16570 1594 16596 1597
rect 16570 1565 16596 1568
rect 16300 1529 16360 1537
rect 16300 1526 16366 1529
rect 16300 1523 16340 1526
rect 16340 1497 16366 1500
rect 16622 1495 16636 1727
rect 16714 1554 16728 1900
rect 16754 1560 16780 1563
rect 16714 1540 16754 1554
rect 16754 1531 16780 1534
rect 16852 1537 16866 1900
rect 16990 1605 17004 1900
rect 16990 1597 17050 1605
rect 16990 1594 17056 1597
rect 16990 1591 17030 1594
rect 17030 1565 17056 1568
rect 16852 1529 16912 1537
rect 16852 1526 16918 1529
rect 16852 1523 16892 1526
rect 16892 1497 16918 1500
rect 16064 1492 16090 1495
rect 16064 1463 16090 1466
rect 16616 1492 16642 1495
rect 17128 1486 17142 1900
rect 17266 1537 17280 1900
rect 17404 1563 17418 1900
rect 17398 1560 17424 1563
rect 17266 1523 17326 1537
rect 17398 1531 17424 1534
rect 17542 1529 17556 1900
rect 17680 1597 17694 1900
rect 17674 1594 17700 1597
rect 17674 1565 17700 1568
rect 17260 1492 17286 1495
rect 17128 1472 17260 1486
rect 16616 1463 16642 1466
rect 17260 1463 17286 1466
rect 17312 1461 17326 1523
rect 17536 1526 17562 1529
rect 17536 1497 17562 1500
rect 17818 1486 17832 1900
rect 17956 1537 17970 1900
rect 17956 1523 18016 1537
rect 17950 1492 17976 1495
rect 17818 1472 17950 1486
rect 17950 1463 17976 1466
rect 18002 1461 18016 1523
rect 17306 1458 17332 1461
rect 17306 1429 17332 1432
rect 17996 1458 18022 1461
rect 17996 1429 18022 1432
rect 15619 1347 15631 1373
rect 15657 1347 15669 1373
rect 14224 1254 14250 1257
rect 14224 1225 14250 1228
rect 12619 1146 12630 1174
rect 12658 1146 12669 1174
rect 12619 1101 12669 1146
rect 12619 1075 12631 1101
rect 12657 1075 12669 1101
rect 9808 948 9834 951
rect 9808 919 9834 922
rect 10774 948 10800 951
rect 10774 919 10800 922
rect 12154 948 12180 951
rect 12154 919 12180 922
rect 9619 803 9631 829
rect 9657 803 9669 829
rect 8428 676 8454 679
rect 8428 647 8454 650
rect 8842 676 8868 679
rect 8842 647 8868 650
rect 8290 642 8316 645
rect 8290 613 8316 616
rect 8198 608 8224 611
rect 8198 579 8224 582
rect 8204 313 8218 579
rect 8020 300 8080 313
rect 8158 300 8218 313
rect 8296 300 8310 613
rect 8434 300 8448 647
rect 8704 642 8730 645
rect 8704 613 8730 616
rect 8566 608 8592 611
rect 8566 579 8592 582
rect 8572 300 8586 579
rect 8710 300 8724 613
rect 8848 300 8862 647
rect 8980 642 9006 645
rect 8980 613 9006 616
rect 9532 642 9558 645
rect 9532 613 9558 616
rect 9619 634 9669 803
rect 9716 676 9742 679
rect 9716 647 9742 650
rect 8986 300 9000 613
rect 9118 608 9144 611
rect 9486 608 9512 611
rect 9118 579 9144 582
rect 9262 588 9486 602
rect 9124 300 9138 579
rect 9262 300 9276 588
rect 9486 579 9512 582
rect 9394 370 9420 373
rect 9394 341 9420 344
rect 9400 300 9414 341
rect 9538 300 9552 613
rect 9619 606 9630 634
rect 9658 606 9669 634
rect 9619 520 9669 606
rect 9722 313 9736 647
rect 9676 300 9736 313
rect 9814 300 9828 919
rect 10084 676 10110 679
rect 10084 647 10110 650
rect 10498 676 10524 679
rect 10498 647 10524 650
rect 9946 642 9972 645
rect 9946 613 9972 616
rect 9952 300 9966 613
rect 10090 300 10104 647
rect 10360 642 10386 645
rect 10360 613 10386 616
rect 10130 608 10156 611
rect 10314 608 10340 611
rect 10130 579 10156 582
rect 10228 588 10314 602
rect 10136 373 10150 579
rect 10130 370 10156 373
rect 10130 341 10156 344
rect 10228 300 10242 588
rect 10314 579 10340 582
rect 10366 300 10380 613
rect 10504 300 10518 647
rect 10636 608 10662 611
rect 10636 579 10662 582
rect 10642 300 10656 579
rect 10780 300 10794 919
rect 11188 676 11214 679
rect 11188 647 11214 650
rect 11740 676 11766 679
rect 11740 647 11766 650
rect 10912 642 10938 645
rect 10912 613 10938 616
rect 10918 300 10932 613
rect 11050 608 11076 611
rect 11050 579 11076 582
rect 11056 300 11070 579
rect 11194 300 11208 647
rect 11326 642 11352 645
rect 11326 613 11352 616
rect 11464 642 11490 645
rect 11464 613 11490 616
rect 11332 300 11346 613
rect 11470 300 11484 613
rect 11694 608 11720 611
rect 11608 588 11694 602
rect 11608 300 11622 588
rect 11694 579 11720 582
rect 11746 300 11760 647
rect 11878 642 11904 645
rect 11878 613 11904 616
rect 11884 300 11898 613
rect 12016 608 12042 611
rect 12016 579 12042 582
rect 12022 300 12036 579
rect 12160 300 12174 919
rect 12430 676 12456 679
rect 12430 647 12456 650
rect 12338 642 12364 645
rect 12338 613 12364 616
rect 12344 313 12358 613
rect 12298 300 12358 313
rect 12436 300 12450 647
rect 12568 608 12594 611
rect 12568 579 12594 582
rect 12574 300 12588 579
rect 12619 557 12669 1075
rect 14224 948 14250 951
rect 14224 919 14250 922
rect 15328 948 15354 951
rect 15328 919 15354 922
rect 13258 710 13284 713
rect 13258 681 13284 684
rect 13948 710 13974 713
rect 13948 681 13974 684
rect 12982 676 13008 679
rect 12982 647 13008 650
rect 12844 642 12870 645
rect 12844 613 12870 616
rect 12619 531 12631 557
rect 12657 531 12669 557
rect 12619 520 12669 531
rect 12706 370 12732 373
rect 12706 341 12732 344
rect 12712 300 12726 341
rect 12850 300 12864 613
rect 12988 300 13002 647
rect 13074 608 13100 611
rect 13074 579 13100 582
rect 13120 608 13146 611
rect 13120 579 13146 582
rect 13080 373 13094 579
rect 13074 370 13100 373
rect 13074 341 13100 344
rect 13126 300 13140 579
rect 13264 300 13278 681
rect 13672 676 13698 679
rect 13672 647 13698 650
rect 13396 642 13422 645
rect 13396 613 13422 616
rect 13402 300 13416 613
rect 13534 370 13560 373
rect 13534 341 13560 344
rect 13540 300 13554 341
rect 13678 300 13692 647
rect 13810 642 13836 645
rect 13810 613 13836 616
rect 13816 300 13830 613
rect 13954 300 13968 681
rect 14086 642 14112 645
rect 14086 613 14112 616
rect 14092 300 14106 613
rect 14230 300 14244 919
rect 14776 676 14802 679
rect 14776 647 14802 650
rect 14500 642 14526 645
rect 14500 613 14526 616
rect 14316 608 14342 611
rect 14316 579 14342 582
rect 14362 608 14388 611
rect 14362 579 14388 582
rect 14322 373 14336 579
rect 14316 370 14342 373
rect 14316 341 14342 344
rect 14368 300 14382 579
rect 14506 300 14520 613
rect 14638 404 14664 407
rect 14638 375 14664 378
rect 14644 300 14658 375
rect 14782 300 14796 647
rect 14960 642 14986 645
rect 14920 622 14960 636
rect 14920 300 14934 622
rect 14960 613 14986 616
rect 15190 608 15216 611
rect 15190 579 15216 582
rect 15052 370 15078 373
rect 15052 341 15078 344
rect 15058 300 15072 341
rect 15196 300 15210 579
rect 15334 300 15348 919
rect 15619 829 15669 1347
rect 18094 1257 18108 1900
rect 18232 1563 18246 1900
rect 18370 1597 18384 1900
rect 18364 1594 18390 1597
rect 18364 1565 18390 1568
rect 18226 1560 18252 1563
rect 18226 1531 18252 1534
rect 18508 1529 18522 1900
rect 18646 1741 18660 1900
rect 18646 1727 18706 1741
rect 18619 1645 18669 1656
rect 18619 1619 18631 1645
rect 18657 1619 18669 1645
rect 18502 1526 18528 1529
rect 18502 1497 18528 1500
rect 18088 1254 18114 1257
rect 18088 1225 18114 1228
rect 18619 1174 18669 1619
rect 18692 1495 18706 1727
rect 18784 1563 18798 1900
rect 18922 1597 18936 1900
rect 18916 1594 18942 1597
rect 18916 1565 18942 1568
rect 18778 1560 18804 1563
rect 18778 1531 18804 1534
rect 19060 1529 19074 1900
rect 19054 1526 19080 1529
rect 19054 1497 19080 1500
rect 19198 1495 19212 1900
rect 19336 1563 19350 1900
rect 19474 1597 19488 1900
rect 19468 1594 19494 1597
rect 19468 1565 19494 1568
rect 19330 1560 19356 1563
rect 19330 1531 19356 1534
rect 19612 1529 19626 1900
rect 19606 1526 19632 1529
rect 19606 1497 19632 1500
rect 19750 1495 19764 1900
rect 19888 1563 19902 1900
rect 20026 1588 20040 1900
rect 20066 1594 20092 1597
rect 20026 1574 20066 1588
rect 20066 1565 20092 1568
rect 19882 1560 19908 1563
rect 19882 1531 19908 1534
rect 20164 1537 20178 1900
rect 20164 1529 20224 1537
rect 20164 1526 20230 1529
rect 20164 1523 20204 1526
rect 20204 1497 20230 1500
rect 18686 1492 18712 1495
rect 18686 1463 18712 1466
rect 19192 1492 19218 1495
rect 19192 1463 19218 1466
rect 19744 1492 19770 1495
rect 20302 1486 20316 1900
rect 20342 1492 20368 1495
rect 20302 1472 20342 1486
rect 19744 1463 19770 1466
rect 20342 1463 20368 1466
rect 20440 1461 20454 1900
rect 20578 1588 20592 1900
rect 20618 1594 20644 1597
rect 20578 1574 20618 1588
rect 20618 1565 20644 1568
rect 20434 1458 20460 1461
rect 20434 1429 20460 1432
rect 20716 1257 20730 1900
rect 20854 1597 20868 1900
rect 20848 1594 20874 1597
rect 20848 1565 20874 1568
rect 20992 1563 21006 1900
rect 20986 1560 21012 1563
rect 20986 1531 21012 1534
rect 21130 1537 21144 1900
rect 21268 1588 21282 1900
rect 21406 1673 21420 1900
rect 21406 1659 21466 1673
rect 21400 1594 21426 1597
rect 21268 1574 21400 1588
rect 21400 1565 21426 1568
rect 21130 1529 21190 1537
rect 21130 1526 21196 1529
rect 21130 1523 21170 1526
rect 21170 1497 21196 1500
rect 21452 1495 21466 1659
rect 21544 1563 21558 1900
rect 21682 1741 21696 1900
rect 21682 1727 21788 1741
rect 21538 1560 21564 1563
rect 21538 1531 21564 1534
rect 21446 1492 21472 1495
rect 21446 1463 21472 1466
rect 21619 1373 21669 1656
rect 21774 1597 21788 1727
rect 21768 1594 21794 1597
rect 21768 1565 21794 1568
rect 21820 1529 21834 1900
rect 21814 1526 21840 1529
rect 21814 1497 21840 1500
rect 21958 1495 21972 1900
rect 21952 1492 21978 1495
rect 21952 1463 21978 1466
rect 21619 1347 21631 1373
rect 21657 1347 21669 1373
rect 20710 1254 20736 1257
rect 20710 1225 20736 1228
rect 18619 1146 18630 1174
rect 18658 1146 18669 1174
rect 18619 1101 18669 1146
rect 18619 1075 18631 1101
rect 18657 1075 18669 1101
rect 15880 948 15906 951
rect 15880 919 15906 922
rect 15619 803 15631 829
rect 15657 803 15669 829
rect 15466 676 15492 679
rect 15466 647 15492 650
rect 15420 608 15446 611
rect 15420 579 15446 582
rect 15426 407 15440 579
rect 15420 404 15446 407
rect 15420 375 15446 378
rect 15472 300 15486 647
rect 15619 634 15669 803
rect 15512 608 15538 611
rect 15512 579 15538 582
rect 15619 606 15630 634
rect 15658 606 15669 634
rect 15518 373 15532 579
rect 15619 520 15669 606
rect 15788 608 15814 611
rect 15702 588 15788 602
rect 15512 370 15538 373
rect 15512 341 15538 344
rect 15702 313 15716 588
rect 15788 579 15814 582
rect 15742 370 15768 373
rect 15742 341 15768 344
rect 15610 300 15716 313
rect 15748 300 15762 341
rect 15886 300 15900 919
rect 16156 676 16182 679
rect 16616 676 16642 679
rect 16156 647 16182 650
rect 16576 656 16616 670
rect 16018 642 16044 645
rect 16018 613 16044 616
rect 16024 300 16038 613
rect 16162 300 16176 647
rect 16478 642 16504 645
rect 16438 622 16478 636
rect 16202 608 16228 611
rect 16340 608 16366 611
rect 16202 579 16228 582
rect 16300 588 16340 602
rect 16208 373 16222 579
rect 16202 370 16228 373
rect 16202 341 16228 344
rect 16300 300 16314 588
rect 16340 579 16366 582
rect 16438 300 16452 622
rect 16478 613 16504 616
rect 16576 300 16590 656
rect 17030 676 17056 679
rect 16616 647 16642 650
rect 16990 656 17030 670
rect 16892 642 16918 645
rect 16852 622 16892 636
rect 16754 608 16780 611
rect 16714 588 16754 602
rect 16714 300 16728 588
rect 16754 579 16780 582
rect 16852 300 16866 622
rect 16892 613 16918 616
rect 16990 300 17004 656
rect 17030 647 17056 650
rect 17812 676 17838 679
rect 18318 676 18344 679
rect 17812 647 17838 650
rect 18232 656 18318 670
rect 17306 642 17332 645
rect 17266 622 17306 636
rect 17168 608 17194 611
rect 17128 588 17168 602
rect 17128 300 17142 588
rect 17168 579 17194 582
rect 17266 300 17280 622
rect 17306 613 17332 616
rect 17674 642 17700 645
rect 17674 613 17700 616
rect 17398 404 17424 407
rect 17398 375 17424 378
rect 17404 300 17418 375
rect 17536 370 17562 373
rect 17536 341 17562 344
rect 17542 300 17556 341
rect 17680 300 17694 613
rect 17818 300 17832 647
rect 18180 642 18206 645
rect 18094 622 18180 636
rect 17858 608 17884 611
rect 17858 579 17884 582
rect 17904 608 17930 611
rect 18042 608 18068 611
rect 17904 579 17930 582
rect 17956 588 18042 602
rect 17864 407 17878 579
rect 17858 404 17884 407
rect 17858 375 17884 378
rect 17910 373 17924 579
rect 17904 370 17930 373
rect 17904 341 17930 344
rect 17956 300 17970 588
rect 18042 579 18068 582
rect 18094 300 18108 622
rect 18180 613 18206 616
rect 18232 300 18246 656
rect 18318 647 18344 650
rect 18456 608 18482 611
rect 18370 588 18456 602
rect 18370 300 18384 588
rect 18456 579 18482 582
rect 18619 557 18669 1075
rect 21619 829 21669 1347
rect 22096 1257 22110 1900
rect 22234 1597 22248 1900
rect 22228 1594 22254 1597
rect 22228 1565 22254 1568
rect 22372 1563 22386 1900
rect 22366 1560 22392 1563
rect 22366 1531 22392 1534
rect 22510 1529 22524 1900
rect 22504 1526 22530 1529
rect 22504 1497 22530 1500
rect 22648 1257 22662 1900
rect 22786 1257 22800 1900
rect 22924 1257 22938 1900
rect 23062 1257 23076 1900
rect 23200 1257 23214 1900
rect 23338 1257 23352 1900
rect 23476 1257 23490 1900
rect 23614 1257 23628 1900
rect 23752 1597 23766 1900
rect 23746 1594 23772 1597
rect 23746 1565 23772 1568
rect 23890 1529 23904 1900
rect 23884 1526 23910 1529
rect 23884 1497 23910 1500
rect 24028 1257 24042 1900
rect 24166 1257 24180 1900
rect 24304 1597 24318 1900
rect 24442 1597 24456 1900
rect 24580 1597 24594 1900
rect 24619 1645 24669 1656
rect 24619 1619 24631 1645
rect 24657 1619 24669 1645
rect 24298 1594 24324 1597
rect 24298 1565 24324 1568
rect 24436 1594 24462 1597
rect 24436 1565 24462 1568
rect 24574 1594 24600 1597
rect 24574 1565 24600 1568
rect 22090 1254 22116 1257
rect 22090 1225 22116 1228
rect 22642 1254 22668 1257
rect 22642 1225 22668 1228
rect 22780 1254 22806 1257
rect 22780 1225 22806 1228
rect 22918 1254 22944 1257
rect 22918 1225 22944 1228
rect 23056 1254 23082 1257
rect 23056 1225 23082 1228
rect 23194 1254 23220 1257
rect 23194 1225 23220 1228
rect 23332 1254 23358 1257
rect 23332 1225 23358 1228
rect 23470 1254 23496 1257
rect 23470 1225 23496 1228
rect 23608 1254 23634 1257
rect 23608 1225 23634 1228
rect 24022 1254 24048 1257
rect 24022 1225 24048 1228
rect 24160 1254 24186 1257
rect 24160 1225 24186 1228
rect 24619 1174 24669 1619
rect 24718 1597 24732 1900
rect 24856 1597 24870 1900
rect 24994 1597 25008 1900
rect 24712 1594 24738 1597
rect 24712 1565 24738 1568
rect 24850 1594 24876 1597
rect 24850 1565 24876 1568
rect 24988 1594 25014 1597
rect 24988 1565 25014 1568
rect 25132 1563 25146 1900
rect 25270 1597 25284 1900
rect 25264 1594 25290 1597
rect 25408 1588 25422 1900
rect 25546 1673 25560 1900
rect 25546 1659 25606 1673
rect 25540 1594 25566 1597
rect 25408 1574 25540 1588
rect 25264 1565 25290 1568
rect 25540 1565 25566 1568
rect 25126 1560 25152 1563
rect 25126 1531 25152 1534
rect 25592 1529 25606 1659
rect 25684 1597 25698 1900
rect 25678 1594 25704 1597
rect 25678 1565 25704 1568
rect 25822 1563 25836 1900
rect 25960 1597 25974 1900
rect 25954 1594 25980 1597
rect 26098 1588 26112 1900
rect 26236 1673 26250 1900
rect 26236 1659 26296 1673
rect 26230 1594 26256 1597
rect 26098 1574 26230 1588
rect 25954 1565 25980 1568
rect 26230 1565 26256 1568
rect 25816 1560 25842 1563
rect 25816 1531 25842 1534
rect 26282 1529 26296 1659
rect 26374 1597 26388 1900
rect 26368 1594 26394 1597
rect 26368 1565 26394 1568
rect 26512 1563 26526 1900
rect 26650 1597 26664 1900
rect 26644 1594 26670 1597
rect 26788 1588 26802 1900
rect 26926 1673 26940 1900
rect 26926 1659 26986 1673
rect 26920 1594 26946 1597
rect 26788 1574 26920 1588
rect 26644 1565 26670 1568
rect 26920 1565 26946 1568
rect 26972 1563 26986 1659
rect 27064 1597 27078 1900
rect 27058 1594 27084 1597
rect 27058 1565 27084 1568
rect 27202 1563 27216 1900
rect 27340 1597 27354 1900
rect 27334 1594 27360 1597
rect 27334 1565 27360 1568
rect 27478 1563 27492 1900
rect 27616 1741 27630 1900
rect 27616 1727 27722 1741
rect 26506 1560 26532 1563
rect 26506 1531 26532 1534
rect 26966 1560 26992 1563
rect 26966 1531 26992 1534
rect 27196 1560 27222 1563
rect 27196 1531 27222 1534
rect 27472 1560 27498 1563
rect 27472 1531 27498 1534
rect 25586 1526 25612 1529
rect 25586 1497 25612 1500
rect 26276 1526 26302 1529
rect 26276 1497 26302 1500
rect 24619 1146 24630 1174
rect 24658 1146 24669 1174
rect 24619 1101 24669 1146
rect 24619 1075 24631 1101
rect 24657 1075 24669 1101
rect 22504 982 22530 985
rect 22504 953 22530 956
rect 21722 948 21748 951
rect 21722 919 21748 922
rect 22228 948 22254 951
rect 22228 919 22254 922
rect 21619 803 21631 829
rect 21657 803 21669 829
rect 19468 710 19494 713
rect 19468 681 19494 684
rect 20710 710 20736 713
rect 20710 681 20736 684
rect 18778 676 18804 679
rect 18738 656 18778 670
rect 18686 642 18712 645
rect 18686 613 18712 616
rect 18619 531 18631 557
rect 18657 531 18669 557
rect 18619 520 18669 531
rect 18692 381 18706 613
rect 18508 367 18706 381
rect 18508 300 18522 367
rect 18738 313 18752 656
rect 19192 676 19218 679
rect 18778 647 18804 650
rect 19106 656 19192 670
rect 19054 642 19080 645
rect 18968 622 19054 636
rect 18916 608 18942 611
rect 18646 300 18752 313
rect 18784 588 18916 602
rect 18784 300 18798 588
rect 18916 579 18942 582
rect 18968 313 18982 622
rect 19054 613 19080 616
rect 19106 313 19120 656
rect 19192 647 19218 650
rect 19330 608 19356 611
rect 18922 300 18982 313
rect 19060 300 19120 313
rect 19198 588 19330 602
rect 19198 300 19212 588
rect 19330 579 19356 582
rect 19330 370 19356 373
rect 19330 341 19356 344
rect 19336 300 19350 341
rect 19474 300 19488 681
rect 19744 676 19770 679
rect 20388 676 20414 679
rect 19744 647 19770 650
rect 20302 656 20388 670
rect 19606 642 19632 645
rect 19606 613 19632 616
rect 19612 300 19626 613
rect 19750 300 19764 647
rect 19836 608 19862 611
rect 19836 579 19862 582
rect 19882 608 19908 611
rect 20250 608 20276 611
rect 19882 579 19908 582
rect 20164 588 20250 602
rect 19842 373 19856 579
rect 19836 370 19862 373
rect 19836 341 19862 344
rect 19888 300 19902 579
rect 20020 370 20046 373
rect 20020 341 20046 344
rect 20026 300 20040 341
rect 20164 300 20178 588
rect 20250 579 20276 582
rect 20302 300 20316 656
rect 20388 647 20414 650
rect 20440 639 20684 653
rect 20440 300 20454 639
rect 20670 611 20684 639
rect 20618 608 20644 611
rect 20618 579 20644 582
rect 20664 608 20690 611
rect 20664 579 20690 582
rect 20572 404 20598 407
rect 20572 375 20598 378
rect 20578 300 20592 375
rect 20624 373 20638 579
rect 20618 370 20644 373
rect 20618 341 20644 344
rect 20716 300 20730 681
rect 21538 676 21564 679
rect 21538 647 21564 650
rect 21262 642 21288 645
rect 21262 613 21288 616
rect 21124 472 21150 475
rect 21124 443 21150 446
rect 20986 438 21012 441
rect 20986 409 21012 412
rect 20848 370 20874 373
rect 20848 341 20874 344
rect 20854 300 20868 341
rect 20992 300 21006 409
rect 21130 300 21144 443
rect 21268 300 21282 613
rect 21308 608 21334 611
rect 21308 579 21334 582
rect 21400 608 21426 611
rect 21400 579 21426 582
rect 21314 407 21328 579
rect 21308 404 21334 407
rect 21308 375 21334 378
rect 21406 373 21420 579
rect 21400 370 21426 373
rect 21400 341 21426 344
rect 21446 336 21472 339
rect 21406 310 21446 313
rect 21406 307 21472 310
rect 21406 300 21466 307
rect 21544 300 21558 647
rect 21619 634 21669 803
rect 21619 606 21630 634
rect 21658 606 21669 634
rect 21619 520 21669 606
rect 21728 449 21742 919
rect 21814 642 21840 645
rect 21814 613 21840 616
rect 21682 435 21742 449
rect 21682 300 21696 435
rect 21820 300 21834 613
rect 21906 608 21932 611
rect 21906 579 21932 582
rect 22044 608 22070 611
rect 22044 579 22070 582
rect 21912 441 21926 579
rect 22050 475 22064 579
rect 22044 472 22070 475
rect 22044 443 22070 446
rect 21906 438 21932 441
rect 21906 409 21932 412
rect 22090 404 22116 407
rect 22090 375 22116 378
rect 21952 370 21978 373
rect 21952 341 21978 344
rect 21958 300 21972 341
rect 22096 300 22110 375
rect 22234 300 22248 919
rect 22366 642 22392 645
rect 22366 613 22392 616
rect 22320 608 22346 611
rect 22320 579 22346 582
rect 22326 339 22340 579
rect 22320 336 22346 339
rect 22320 307 22346 310
rect 22372 300 22386 613
rect 22510 300 22524 953
rect 22918 710 22944 713
rect 22918 681 22944 684
rect 23700 710 23726 713
rect 23700 681 23726 684
rect 24436 710 24462 713
rect 24436 681 24462 684
rect 22642 676 22668 679
rect 22642 647 22668 650
rect 22648 300 22662 647
rect 22734 608 22760 611
rect 22734 579 22760 582
rect 22780 608 22806 611
rect 22780 579 22806 582
rect 22740 373 22754 579
rect 22734 370 22760 373
rect 22734 341 22760 344
rect 22786 300 22800 579
rect 22924 300 22938 681
rect 23240 676 23266 679
rect 23200 656 23240 670
rect 23056 608 23082 611
rect 23056 579 23082 582
rect 23102 608 23128 611
rect 23102 579 23128 582
rect 23062 407 23076 579
rect 23056 404 23082 407
rect 23056 375 23082 378
rect 23108 313 23122 579
rect 23062 300 23122 313
rect 23200 300 23214 656
rect 23240 647 23266 650
rect 23654 642 23680 645
rect 23654 613 23680 616
rect 23470 608 23496 611
rect 23338 588 23470 602
rect 23338 300 23352 588
rect 23470 579 23496 582
rect 23660 364 23674 613
rect 23476 350 23674 364
rect 23476 300 23490 350
rect 23706 313 23720 681
rect 24344 676 24370 679
rect 24258 656 24344 670
rect 24206 642 24232 645
rect 24206 613 24232 616
rect 24068 608 24094 611
rect 23614 300 23720 313
rect 23752 588 24068 602
rect 23752 300 23766 588
rect 24068 579 24094 582
rect 23884 370 23910 373
rect 24212 364 24226 613
rect 23884 341 23910 344
rect 24028 350 24226 364
rect 23890 300 23904 341
rect 24028 300 24042 350
rect 24258 313 24272 656
rect 24344 647 24370 650
rect 24298 404 24324 407
rect 24298 375 24324 378
rect 24166 300 24272 313
rect 24304 300 24318 375
rect 24442 300 24456 681
rect 24574 608 24600 611
rect 24574 579 24600 582
rect 24580 373 24594 579
rect 24619 557 24669 1075
rect 27619 1373 27669 1656
rect 27708 1597 27722 1727
rect 27702 1594 27728 1597
rect 27702 1565 27728 1568
rect 27754 1495 27768 1900
rect 27892 1529 27906 1900
rect 28030 1597 28044 1900
rect 28024 1594 28050 1597
rect 28024 1565 28050 1568
rect 28168 1537 28182 1900
rect 28306 1605 28320 1900
rect 28306 1597 28366 1605
rect 28306 1594 28372 1597
rect 28306 1591 28346 1594
rect 28346 1565 28372 1568
rect 28444 1554 28458 1900
rect 28484 1560 28510 1563
rect 28444 1540 28484 1554
rect 28168 1529 28320 1537
rect 28484 1531 28510 1534
rect 28582 1529 28596 1900
rect 28720 1605 28734 1900
rect 28858 1605 28872 1900
rect 28996 1673 29010 1900
rect 28996 1659 29056 1673
rect 28720 1597 28780 1605
rect 28720 1594 28786 1597
rect 28720 1591 28760 1594
rect 28858 1591 29010 1605
rect 28760 1565 28786 1568
rect 28996 1563 29010 1591
rect 28990 1560 29016 1563
rect 28990 1531 29016 1534
rect 29042 1529 29056 1659
rect 29134 1597 29148 1900
rect 29128 1594 29154 1597
rect 29128 1565 29154 1568
rect 29272 1563 29286 1900
rect 29266 1560 29292 1563
rect 29266 1531 29292 1534
rect 29410 1529 29424 1900
rect 29548 1597 29562 1900
rect 29542 1594 29568 1597
rect 29542 1565 29568 1568
rect 29686 1563 29700 1900
rect 29680 1560 29706 1563
rect 29680 1531 29706 1534
rect 29824 1529 29838 1900
rect 29962 1597 29976 1900
rect 29956 1594 29982 1597
rect 29956 1565 29982 1568
rect 30100 1563 30114 1900
rect 30238 1605 30252 1900
rect 30376 1673 30390 1900
rect 30376 1659 30436 1673
rect 30238 1597 30390 1605
rect 30238 1594 30396 1597
rect 30238 1591 30370 1594
rect 30370 1565 30396 1568
rect 30094 1560 30120 1563
rect 30094 1531 30120 1534
rect 30422 1529 30436 1659
rect 30514 1563 30528 1900
rect 30652 1741 30666 1900
rect 30652 1727 30712 1741
rect 30619 1645 30669 1656
rect 30619 1619 30631 1645
rect 30657 1619 30669 1645
rect 30508 1560 30534 1563
rect 30508 1531 30534 1534
rect 27886 1526 27912 1529
rect 28168 1526 28326 1529
rect 28168 1523 28300 1526
rect 27886 1497 27912 1500
rect 28300 1497 28326 1500
rect 28576 1526 28602 1529
rect 28576 1497 28602 1500
rect 29036 1526 29062 1529
rect 29036 1497 29062 1500
rect 29404 1526 29430 1529
rect 29404 1497 29430 1500
rect 29818 1526 29844 1529
rect 29818 1497 29844 1500
rect 30416 1526 30442 1529
rect 30416 1497 30442 1500
rect 27748 1492 27774 1495
rect 27748 1463 27774 1466
rect 27619 1347 27631 1373
rect 27657 1347 27669 1373
rect 25540 948 25566 951
rect 25540 919 25566 922
rect 24942 710 24968 713
rect 24942 681 24968 684
rect 25402 710 25428 713
rect 25402 681 25428 684
rect 24758 642 24784 645
rect 24758 613 24784 616
rect 24619 531 24631 557
rect 24657 531 24669 557
rect 24619 520 24669 531
rect 24574 370 24600 373
rect 24764 364 24778 613
rect 24574 341 24600 344
rect 24626 350 24778 364
rect 24626 313 24640 350
rect 24948 313 24962 681
rect 24988 608 25014 611
rect 24988 579 25014 582
rect 25034 608 25060 611
rect 25034 579 25060 582
rect 24994 407 25008 579
rect 24988 404 25014 407
rect 24988 375 25014 378
rect 25040 313 25054 579
rect 25264 404 25290 407
rect 25264 375 25290 378
rect 25126 370 25152 373
rect 25126 341 25152 344
rect 24580 300 24640 313
rect 24718 305 24778 313
rect 24718 302 24784 305
rect 24718 300 24758 302
rect 2033 287 2061 292
rect 2079 0 2107 300
rect 2217 299 2284 300
rect 2217 0 2245 299
rect 2355 0 2383 300
rect 2493 0 2521 300
rect 2631 0 2659 300
rect 2769 0 2797 300
rect 2907 0 2935 300
rect 3045 299 3112 300
rect 3045 0 3073 299
rect 3183 0 3211 300
rect 3321 0 3349 300
rect 3459 0 3487 300
rect 3597 299 3710 300
rect 3597 0 3625 299
rect 3735 0 3763 300
rect 3873 0 3901 300
rect 4011 0 4039 300
rect 4149 0 4177 300
rect 4287 0 4315 300
rect 4425 0 4453 300
rect 4563 299 4630 300
rect 4563 0 4591 299
rect 4701 0 4729 300
rect 4839 0 4867 300
rect 4977 0 5005 300
rect 5115 0 5143 300
rect 5253 0 5281 300
rect 5391 0 5419 300
rect 5529 0 5557 300
rect 5667 0 5695 300
rect 5805 0 5833 300
rect 5943 0 5971 300
rect 6081 0 6109 300
rect 6219 0 6247 300
rect 6357 0 6385 300
rect 6495 0 6523 300
rect 6633 299 6746 300
rect 6633 0 6661 299
rect 6771 0 6799 300
rect 6909 0 6937 300
rect 7047 0 7075 300
rect 7185 0 7213 300
rect 7323 0 7351 300
rect 7461 299 7528 300
rect 7461 0 7489 299
rect 7599 0 7627 300
rect 7737 0 7765 300
rect 7875 0 7903 300
rect 8013 299 8080 300
rect 8151 299 8218 300
rect 8013 0 8041 299
rect 8151 0 8179 299
rect 8289 0 8317 300
rect 8427 0 8455 300
rect 8565 0 8593 300
rect 8703 0 8731 300
rect 8841 0 8869 300
rect 8979 0 9007 300
rect 9117 0 9145 300
rect 9255 0 9283 300
rect 9393 0 9421 300
rect 9531 0 9559 300
rect 9669 299 9736 300
rect 9669 0 9697 299
rect 9807 0 9835 300
rect 9945 0 9973 300
rect 10083 0 10111 300
rect 10221 0 10249 300
rect 10359 0 10387 300
rect 10497 0 10525 300
rect 10635 0 10663 300
rect 10773 0 10801 300
rect 10911 0 10939 300
rect 11049 0 11077 300
rect 11187 0 11215 300
rect 11325 0 11353 300
rect 11463 0 11491 300
rect 11601 0 11629 300
rect 11739 0 11767 300
rect 11877 0 11905 300
rect 12015 0 12043 300
rect 12153 0 12181 300
rect 12291 299 12358 300
rect 12291 0 12319 299
rect 12429 0 12457 300
rect 12567 0 12595 300
rect 12705 0 12733 300
rect 12843 0 12871 300
rect 12981 0 13009 300
rect 13119 0 13147 300
rect 13257 0 13285 300
rect 13395 0 13423 300
rect 13533 0 13561 300
rect 13671 0 13699 300
rect 13809 0 13837 300
rect 13947 0 13975 300
rect 14085 0 14113 300
rect 14223 0 14251 300
rect 14361 0 14389 300
rect 14499 0 14527 300
rect 14637 0 14665 300
rect 14775 0 14803 300
rect 14913 0 14941 300
rect 15051 0 15079 300
rect 15189 0 15217 300
rect 15327 0 15355 300
rect 15465 0 15493 300
rect 15603 299 15716 300
rect 15603 0 15631 299
rect 15741 0 15769 300
rect 15879 0 15907 300
rect 16017 0 16045 300
rect 16155 0 16183 300
rect 16293 0 16321 300
rect 16431 0 16459 300
rect 16569 0 16597 300
rect 16707 0 16735 300
rect 16845 0 16873 300
rect 16983 0 17011 300
rect 17121 0 17149 300
rect 17259 0 17287 300
rect 17397 0 17425 300
rect 17535 0 17563 300
rect 17673 0 17701 300
rect 17811 0 17839 300
rect 17949 0 17977 300
rect 18087 0 18115 300
rect 18225 0 18253 300
rect 18363 0 18391 300
rect 18501 0 18529 300
rect 18639 299 18752 300
rect 18639 0 18667 299
rect 18777 0 18805 300
rect 18915 299 18982 300
rect 19053 299 19120 300
rect 18915 0 18943 299
rect 19053 0 19081 299
rect 19191 0 19219 300
rect 19329 0 19357 300
rect 19467 0 19495 300
rect 19605 0 19633 300
rect 19743 0 19771 300
rect 19881 0 19909 300
rect 20019 0 20047 300
rect 20157 0 20185 300
rect 20295 0 20323 300
rect 20433 0 20461 300
rect 20571 0 20599 300
rect 20709 0 20737 300
rect 20847 0 20875 300
rect 20985 0 21013 300
rect 21123 0 21151 300
rect 21261 0 21289 300
rect 21399 299 21466 300
rect 21399 0 21427 299
rect 21537 0 21565 300
rect 21675 0 21703 300
rect 21813 0 21841 300
rect 21951 0 21979 300
rect 22089 0 22117 300
rect 22227 0 22255 300
rect 22365 0 22393 300
rect 22503 0 22531 300
rect 22641 0 22669 300
rect 22779 0 22807 300
rect 22917 0 22945 300
rect 23055 299 23122 300
rect 23055 0 23083 299
rect 23193 0 23221 300
rect 23331 0 23359 300
rect 23469 0 23497 300
rect 23607 299 23720 300
rect 23607 0 23635 299
rect 23745 0 23773 300
rect 23883 0 23911 300
rect 24021 0 24049 300
rect 24159 299 24272 300
rect 24159 0 24187 299
rect 24297 0 24325 300
rect 24435 0 24463 300
rect 24573 299 24640 300
rect 24711 299 24758 300
rect 24573 0 24601 299
rect 24711 0 24739 299
rect 24856 300 24962 313
rect 24994 300 25054 313
rect 25132 300 25146 341
rect 25270 300 25284 375
rect 25408 300 25422 681
rect 25448 608 25474 611
rect 25448 579 25474 582
rect 25454 305 25468 579
rect 25448 302 25474 305
rect 24758 273 24784 276
rect 24849 299 24962 300
rect 24987 299 25054 300
rect 24849 0 24877 299
rect 24987 0 25015 299
rect 25125 0 25153 300
rect 25263 0 25291 300
rect 25401 0 25429 300
rect 25546 300 25560 919
rect 27619 829 27669 1347
rect 27619 803 27631 829
rect 27657 803 27669 829
rect 25816 676 25842 679
rect 26506 676 26532 679
rect 25816 647 25842 650
rect 26374 656 26506 670
rect 25678 642 25704 645
rect 25678 613 25704 616
rect 25684 300 25698 613
rect 25822 300 25836 647
rect 26322 642 26348 645
rect 26322 613 26348 616
rect 25862 608 25888 611
rect 25862 579 25888 582
rect 25908 608 25934 611
rect 26184 608 26210 611
rect 25908 579 25934 582
rect 25960 588 26184 602
rect 25868 373 25882 579
rect 25914 407 25928 579
rect 25908 404 25934 407
rect 25908 375 25934 378
rect 25862 370 25888 373
rect 25862 341 25888 344
rect 25960 300 25974 588
rect 26184 579 26210 582
rect 26328 364 26342 613
rect 26098 350 26342 364
rect 26098 300 26112 350
rect 26236 305 26296 313
rect 26236 302 26302 305
rect 26236 300 26276 302
rect 25448 273 25474 276
rect 25539 0 25567 300
rect 25677 0 25705 300
rect 25815 0 25843 300
rect 25953 0 25981 300
rect 26091 0 26119 300
rect 26229 299 26276 300
rect 26229 0 26257 299
rect 26374 300 26388 656
rect 27334 676 27360 679
rect 26506 647 26532 650
rect 26788 639 26940 653
rect 27334 647 27360 650
rect 26644 608 26670 611
rect 26512 588 26644 602
rect 26512 300 26526 588
rect 26644 579 26670 582
rect 26644 438 26670 441
rect 26644 409 26670 412
rect 26650 300 26664 409
rect 26788 300 26802 639
rect 26926 611 26940 639
rect 26874 608 26900 611
rect 26874 579 26900 582
rect 26920 608 26946 611
rect 26920 579 26946 582
rect 27288 608 27314 611
rect 27288 579 27314 582
rect 26880 305 26894 579
rect 26920 472 26946 475
rect 26920 443 26946 446
rect 26874 302 26900 305
rect 26276 273 26302 276
rect 26367 0 26395 300
rect 26505 0 26533 300
rect 26643 0 26671 300
rect 26781 0 26809 300
rect 26926 300 26940 443
rect 27294 441 27308 579
rect 27288 438 27314 441
rect 27288 409 27314 412
rect 27196 404 27222 407
rect 27196 375 27222 378
rect 27058 370 27084 373
rect 27058 341 27084 344
rect 27064 300 27078 341
rect 27202 300 27216 375
rect 27340 300 27354 647
rect 27472 642 27498 645
rect 27472 613 27498 616
rect 27619 634 27669 803
rect 27478 300 27492 613
rect 27564 608 27590 611
rect 27564 579 27590 582
rect 27619 606 27630 634
rect 27658 606 27669 634
rect 30619 1174 30669 1619
rect 30698 1597 30712 1727
rect 30692 1594 30718 1597
rect 30692 1565 30718 1568
rect 30790 1529 30804 1900
rect 30928 1605 30942 1900
rect 31066 1673 31080 1900
rect 31066 1659 31126 1673
rect 30928 1597 31080 1605
rect 30928 1594 31086 1597
rect 30928 1591 31060 1594
rect 31060 1565 31086 1568
rect 31112 1563 31126 1659
rect 31106 1560 31132 1563
rect 31106 1531 31132 1534
rect 31204 1529 31218 1900
rect 31342 1597 31356 1900
rect 31336 1594 31362 1597
rect 31336 1565 31362 1568
rect 31480 1563 31494 1900
rect 31618 1605 31632 1900
rect 31756 1673 31770 1900
rect 31756 1659 31816 1673
rect 31618 1591 31770 1605
rect 31474 1560 31500 1563
rect 31474 1531 31500 1534
rect 30784 1526 30810 1529
rect 30784 1497 30810 1500
rect 31198 1526 31224 1529
rect 31198 1497 31224 1500
rect 31756 1495 31770 1591
rect 31802 1529 31816 1659
rect 31796 1526 31822 1529
rect 31796 1497 31822 1500
rect 31750 1492 31776 1495
rect 31750 1463 31776 1466
rect 31894 1461 31908 1900
rect 32032 1563 32046 1900
rect 32170 1597 32184 1900
rect 32164 1594 32190 1597
rect 32164 1565 32190 1568
rect 32026 1560 32052 1563
rect 32026 1531 32052 1534
rect 32308 1537 32322 1900
rect 32308 1529 32368 1537
rect 32308 1526 32374 1529
rect 32308 1523 32348 1526
rect 32348 1497 32374 1500
rect 31888 1458 31914 1461
rect 31888 1429 31914 1432
rect 32446 1257 32460 1900
rect 32584 1605 32598 1900
rect 32584 1591 32644 1605
rect 32630 1563 32644 1591
rect 32624 1560 32650 1563
rect 32624 1531 32650 1534
rect 32722 1257 32736 1900
rect 32860 1597 32874 1900
rect 32854 1594 32880 1597
rect 32854 1565 32880 1568
rect 32998 1257 33012 1900
rect 33136 1257 33150 1900
rect 33274 1597 33288 1900
rect 33268 1594 33294 1597
rect 33268 1565 33294 1568
rect 33412 1257 33426 1900
rect 33550 1597 33564 1900
rect 33688 1673 33702 1900
rect 33688 1659 33748 1673
rect 33544 1594 33570 1597
rect 33544 1565 33570 1568
rect 33619 1373 33669 1656
rect 33734 1597 33748 1659
rect 33826 1597 33840 1900
rect 33728 1594 33754 1597
rect 33728 1565 33754 1568
rect 33820 1594 33846 1597
rect 33820 1565 33846 1568
rect 33964 1529 33978 1900
rect 33958 1526 33984 1529
rect 33958 1497 33984 1500
rect 33619 1347 33631 1373
rect 33657 1347 33669 1373
rect 32440 1254 32466 1257
rect 32440 1225 32466 1228
rect 32716 1254 32742 1257
rect 32716 1225 32742 1228
rect 32992 1254 33018 1257
rect 32992 1225 33018 1228
rect 33130 1254 33156 1257
rect 33130 1225 33156 1228
rect 33406 1254 33432 1257
rect 33406 1225 33432 1228
rect 30619 1146 30630 1174
rect 30658 1146 30669 1174
rect 30619 1101 30669 1146
rect 30619 1075 30631 1101
rect 30657 1075 30669 1101
rect 27570 475 27584 579
rect 27619 520 27669 606
rect 27748 608 27774 611
rect 27748 579 27774 582
rect 28162 608 28188 611
rect 28162 579 28188 582
rect 27564 472 27590 475
rect 27564 443 27590 446
rect 27754 373 27768 579
rect 28168 407 28182 579
rect 30619 557 30669 1075
rect 30619 531 30631 557
rect 30657 531 30669 557
rect 30619 520 30669 531
rect 33619 829 33669 1347
rect 33619 803 33631 829
rect 33657 803 33669 829
rect 33619 634 33669 803
rect 33619 606 33630 634
rect 33658 606 33669 634
rect 33619 520 33669 606
rect 28162 404 28188 407
rect 28162 375 28188 378
rect 27748 370 27774 373
rect 27748 341 27774 344
rect 26874 273 26900 276
rect 26919 0 26947 300
rect 27057 0 27085 300
rect 27195 0 27223 300
rect 27333 0 27361 300
rect 27471 0 27499 300
<< via2 >>
rect 1481 1856 1509 1884
rect 1849 1652 1877 1680
rect 1895 1516 1923 1544
rect 2033 1856 2061 1884
rect 1987 1788 2015 1816
rect 2033 1244 2061 1272
rect 2125 1380 2153 1408
rect 1389 990 1390 1000
rect 1390 990 1416 1000
rect 1416 990 1417 1000
rect 1389 972 1417 990
rect 1435 836 1463 864
rect 1481 700 1509 728
rect 1803 1040 1831 1068
rect 1757 428 1785 456
rect 1711 292 1739 320
rect 1849 496 1877 524
rect 1895 292 1923 320
rect 2033 292 2061 320
rect 6630 1146 6658 1174
rect 3630 606 3658 634
rect 12630 1146 12658 1174
rect 9630 606 9658 634
rect 18630 1146 18658 1174
rect 15630 606 15658 634
rect 24630 1146 24658 1174
rect 21630 606 21658 634
rect 27630 606 27658 634
rect 30630 1146 30658 1174
rect 33630 606 33658 634
<< metal3 >>
rect 0 2089 300 2104
rect 0 2059 1809 2089
rect 0 2044 300 2059
rect 0 1953 300 1968
rect 0 1923 1441 1953
rect 0 1908 300 1923
rect 1411 1885 1441 1923
rect 1478 1885 1511 1886
rect 1411 1884 1511 1885
rect 1411 1856 1481 1884
rect 1509 1856 1511 1884
rect 1411 1855 1511 1856
rect 1779 1885 1809 2059
rect 2030 1885 2063 1886
rect 1779 1884 2063 1885
rect 1779 1856 2033 1884
rect 2061 1856 2063 1884
rect 1779 1855 2063 1856
rect 1478 1853 1511 1855
rect 2030 1853 2063 1855
rect 0 1817 300 1832
rect 1984 1817 2017 1818
rect 0 1816 2017 1817
rect 0 1788 1987 1816
rect 2015 1788 2017 1816
rect 0 1787 2017 1788
rect 0 1772 300 1787
rect 1984 1785 2017 1787
rect 0 1681 300 1696
rect 1846 1681 1879 1682
rect 0 1680 1879 1681
rect 0 1652 1849 1680
rect 1877 1652 1879 1680
rect 0 1651 1879 1652
rect 0 1636 300 1651
rect 1846 1649 1879 1651
rect 0 1545 300 1560
rect 1892 1545 1925 1546
rect 0 1544 1925 1545
rect 0 1516 1895 1544
rect 1923 1516 1925 1544
rect 0 1515 1925 1516
rect 0 1500 300 1515
rect 1892 1513 1925 1515
rect 0 1409 300 1424
rect 2122 1409 2155 1410
rect 0 1408 2155 1409
rect 0 1380 2125 1408
rect 2153 1380 2155 1408
rect 0 1379 2155 1380
rect 0 1364 300 1379
rect 2122 1377 2155 1379
rect 0 1273 300 1288
rect 2030 1273 2063 1274
rect 0 1272 2063 1273
rect 0 1244 2033 1272
rect 2061 1244 2063 1272
rect 0 1243 2063 1244
rect 0 1228 300 1243
rect 2030 1241 2063 1243
rect 644 1174 34408 1185
rect 0 1137 300 1152
rect 644 1146 6630 1174
rect 6658 1146 12630 1174
rect 12658 1146 18630 1174
rect 18658 1146 24630 1174
rect 24658 1146 30630 1174
rect 30658 1146 34408 1174
rect 0 1107 613 1137
rect 644 1135 34408 1146
rect 0 1092 300 1107
rect 583 1069 613 1107
rect 1800 1069 1833 1070
rect 583 1068 1833 1069
rect 583 1040 1803 1068
rect 1831 1040 1833 1068
rect 583 1039 1833 1040
rect 1800 1037 1833 1039
rect 0 1001 300 1016
rect 1386 1001 1419 1002
rect 0 1000 1419 1001
rect 0 972 1389 1000
rect 1417 972 1419 1000
rect 0 971 1419 972
rect 0 956 300 971
rect 1386 969 1419 971
rect 0 865 300 880
rect 1432 865 1465 866
rect 0 864 1465 865
rect 0 836 1435 864
rect 1463 836 1465 864
rect 0 835 1465 836
rect 0 820 300 835
rect 1432 833 1465 835
rect 0 729 300 744
rect 1478 729 1511 730
rect 0 728 1511 729
rect 0 700 1481 728
rect 1509 700 1511 728
rect 0 699 1511 700
rect 0 684 300 699
rect 1478 697 1511 699
rect 644 634 34408 645
rect 0 593 300 608
rect 644 606 3630 634
rect 3658 606 9630 634
rect 9658 606 15630 634
rect 15658 606 21630 634
rect 21658 606 27630 634
rect 27658 606 33630 634
rect 33658 606 34408 634
rect 644 595 34408 606
rect 0 563 613 593
rect 0 548 300 563
rect 583 525 613 563
rect 1846 525 1879 526
rect 583 524 1879 525
rect 583 496 1849 524
rect 1877 496 1879 524
rect 583 495 1879 496
rect 1846 493 1879 495
rect 0 457 300 472
rect 1754 457 1787 458
rect 0 456 1787 457
rect 0 428 1757 456
rect 1785 428 1787 456
rect 0 427 1787 428
rect 0 412 300 427
rect 1754 425 1787 427
rect 0 321 300 336
rect 1708 321 1741 322
rect 1892 321 1925 322
rect 2030 321 2063 322
rect 0 320 1741 321
rect 0 292 1711 320
rect 1739 292 1741 320
rect 0 291 1741 292
rect 0 276 300 291
rect 1708 289 1741 291
rect 1779 320 1925 321
rect 1779 292 1895 320
rect 1923 292 1925 320
rect 1779 291 1925 292
rect 0 185 300 200
rect 1779 185 1809 291
rect 1892 289 1925 291
rect 1963 320 2063 321
rect 1963 292 2033 320
rect 2061 292 2063 320
rect 1963 291 2063 292
rect 0 155 1809 185
rect 0 140 300 155
rect 0 49 300 64
rect 1963 49 1993 291
rect 2030 289 2063 291
rect 0 19 1993 49
rect 0 4 300 19
use sky130_fd_sc_hd__fill_2  FILLER_3_729 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 34178 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_3_722 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 33856 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[9\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform -1 0 33856 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 34132 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  PHY_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform -1 0 34408 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[99\]
timestamp 1641350499
transform -1 0 33718 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[98\]
timestamp 1641350499
transform -1 0 33580 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[96\]
timestamp 1641350499
transform 1 0 33304 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[93\]
timestamp 1641350499
transform 1 0 33166 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[91\]
timestamp 1641350499
transform 1 0 33028 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[8\]
timestamp 1641350499
transform 1 0 32706 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[89\]
timestamp 1641350499
transform 1 0 32568 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[343\]
timestamp 1641350499
transform -1 0 33028 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1641350499
transform 1 0 32844 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[88\]
timestamp 1641350499
transform 1 0 32430 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[87\]
timestamp 1641350499
transform 1 0 32292 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[86\]
timestamp 1641350499
transform 1 0 32154 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[85\]
timestamp 1641350499
transform 1 0 32016 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[84\]
timestamp 1641350499
transform 1 0 31878 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[83\]
timestamp 1641350499
transform 1 0 31740 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[82\]
timestamp 1641350499
transform 1 0 31602 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[81\]
timestamp 1641350499
transform 1 0 31418 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1641350499
transform 1 0 31556 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[80\]
timestamp 1641350499
transform 1 0 31280 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[7\]
timestamp 1641350499
transform 1 0 31142 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[79\]
timestamp 1641350499
transform 1 0 31004 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[78\]
timestamp 1641350499
transform 1 0 30866 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[77\]
timestamp 1641350499
transform 1 0 30728 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[76\]
timestamp 1641350499
transform 1 0 30590 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[75\]
timestamp 1641350499
transform 1 0 30452 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[74\]
timestamp 1641350499
transform 1 0 30314 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1641350499
transform 1 0 30268 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[73\]
timestamp 1641350499
transform 1 0 30130 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[72\]
timestamp 1641350499
transform 1 0 29992 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[71\]
timestamp 1641350499
transform 1 0 29854 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[70\]
timestamp 1641350499
transform 1 0 29716 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[6\]
timestamp 1641350499
transform 1 0 29578 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[69\]
timestamp 1641350499
transform 1 0 29440 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[68\]
timestamp 1641350499
transform 1 0 29302 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[67\]
timestamp 1641350499
transform 1 0 29164 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[66\]
timestamp 1641350499
transform 1 0 29026 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[65\]
timestamp 1641350499
transform 1 0 28842 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[64\]
timestamp 1641350499
transform 1 0 28704 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[63\]
timestamp 1641350499
transform 1 0 28566 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[62\]
timestamp 1641350499
transform 1 0 28428 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1641350499
transform 1 0 28980 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[61\]
timestamp 1641350499
transform 1 0 28290 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[60\]
timestamp 1641350499
transform 1 0 28152 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[5\]
timestamp 1641350499
transform 1 0 28014 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[59\]
timestamp 1641350499
transform 1 0 27876 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[58\]
timestamp 1641350499
transform 1 0 27738 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[57\]
timestamp 1641350499
transform 1 0 27554 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[56\]
timestamp 1641350499
transform 1 0 27416 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[55\]
timestamp 1641350499
transform 1 0 27278 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1641350499
transform 1 0 27692 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[54\]
timestamp 1641350499
transform 1 0 27140 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[53\]
timestamp 1641350499
transform 1 0 27002 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[52\]
timestamp 1641350499
transform 1 0 26864 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[51\]
timestamp 1641350499
transform 1 0 26726 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[50\]
timestamp 1641350499
transform 1 0 26588 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[4\]
timestamp 1641350499
transform 1 0 26450 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[49\]
timestamp 1641350499
transform 1 0 26266 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[48\]
timestamp 1641350499
transform 1 0 26128 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1641350499
transform 1 0 26404 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[47\]
timestamp 1641350499
transform 1 0 25990 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[46\]
timestamp 1641350499
transform 1 0 25852 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[462\]
timestamp 1641350499
transform 1 0 25714 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[461\]
timestamp 1641350499
transform 1 0 25576 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_3_530
timestamp 1641350499
transform 1 0 25024 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[460\]
timestamp 1641350499
transform 1 0 25438 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[45\]
timestamp 1641350499
transform 1 0 25300 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[459\]
timestamp 1641350499
transform 1 0 25162 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[458\]
timestamp 1641350499
transform 1 0 24886 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1641350499
transform 1 0 25116 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[457\]
timestamp 1641350499
transform 1 0 24748 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[456\]
timestamp 1641350499
transform 1 0 24610 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[455\]
timestamp 1641350499
transform 1 0 24472 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[454\]
timestamp 1641350499
transform 1 0 24334 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[451\]
timestamp 1641350499
transform 1 0 24012 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[450\]
timestamp 1641350499
transform 1 0 23874 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1641350499
transform 1 0 23828 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_3_511 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 24150 0 -1 1632
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  FILLER_3_498
timestamp 1641350499
transform 1 0 23552 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[442\]
timestamp 1641350499
transform 1 0 22862 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[441\]
timestamp 1641350499
transform 1 0 22724 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[440\]
timestamp 1641350499
transform 1 0 22586 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1641350499
transform 1 0 22540 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_3_486 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 23000 0 -1 1632
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[439\]
timestamp 1641350499
transform 1 0 22402 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[438\]
timestamp 1641350499
transform 1 0 22264 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[437\]
timestamp 1641350499
transform 1 0 22126 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[436\]
timestamp 1641350499
transform 1 0 21988 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[435\]
timestamp 1641350499
transform 1 0 21850 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[434\]
timestamp 1641350499
transform 1 0 21712 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[433\]
timestamp 1641350499
transform 1 0 21574 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[432\]
timestamp 1641350499
transform 1 0 21436 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[431\]
timestamp 1641350499
transform 1 0 21298 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[42\]
timestamp 1641350499
transform 1 0 21114 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[429\]
timestamp 1641350499
transform 1 0 20976 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[428\]
timestamp 1641350499
transform 1 0 20838 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1641350499
transform 1 0 21252 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[427\]
timestamp 1641350499
transform 1 0 20700 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[426\]
timestamp 1641350499
transform 1 0 20562 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[425\]
timestamp 1641350499
transform 1 0 20424 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[424\]
timestamp 1641350499
transform 1 0 20286 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[423\]
timestamp 1641350499
transform 1 0 20148 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[422\]
timestamp 1641350499
transform 1 0 20010 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[421\]
timestamp 1641350499
transform 1 0 19826 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[420\]
timestamp 1641350499
transform 1 0 19688 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[41\]
timestamp 1641350499
transform 1 0 19550 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1641350499
transform 1 0 19964 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[419\]
timestamp 1641350499
transform 1 0 19412 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[418\]
timestamp 1641350499
transform 1 0 19274 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[417\]
timestamp 1641350499
transform 1 0 19136 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[416\]
timestamp 1641350499
transform 1 0 18998 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[415\]
timestamp 1641350499
transform 1 0 18860 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[414\]
timestamp 1641350499
transform 1 0 18722 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[412\]
timestamp 1641350499
transform 1 0 18538 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[411\]
timestamp 1641350499
transform 1 0 18400 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1641350499
transform 1 0 18676 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[410\]
timestamp 1641350499
transform 1 0 18262 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[40\]
timestamp 1641350499
transform 1 0 18124 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[409\]
timestamp 1641350499
transform 1 0 17986 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[408\]
timestamp 1641350499
transform 1 0 17848 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[407\]
timestamp 1641350499
transform 1 0 17710 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[406\]
timestamp 1641350499
transform 1 0 17572 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[405\]
timestamp 1641350499
transform 1 0 17434 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[404\]
timestamp 1641350499
transform 1 0 17250 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1641350499
transform 1 0 17388 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[403\]
timestamp 1641350499
transform 1 0 17112 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[402\]
timestamp 1641350499
transform 1 0 16974 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[401\]
timestamp 1641350499
transform 1 0 16836 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[400\]
timestamp 1641350499
transform 1 0 16698 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[3\]
timestamp 1641350499
transform 1 0 16560 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[39\]
timestamp 1641350499
transform 1 0 16422 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[399\]
timestamp 1641350499
transform 1 0 16284 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[398\]
timestamp 1641350499
transform 1 0 16146 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1641350499
transform 1 0 16100 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[397\]
timestamp 1641350499
transform 1 0 15962 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[396\]
timestamp 1641350499
transform 1 0 15824 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[395\]
timestamp 1641350499
transform 1 0 15686 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[394\]
timestamp 1641350499
transform 1 0 15548 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[393\]
timestamp 1641350499
transform 1 0 15410 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[392\]
timestamp 1641350499
transform 1 0 15272 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[391\]
timestamp 1641350499
transform 1 0 15134 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[390\]
timestamp 1641350499
transform 1 0 14996 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[38\]
timestamp 1641350499
transform 1 0 14858 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[388\]
timestamp 1641350499
transform 1 0 14674 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[387\]
timestamp 1641350499
transform 1 0 14536 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[386\]
timestamp 1641350499
transform 1 0 14398 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[385\]
timestamp 1641350499
transform 1 0 14260 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1641350499
transform 1 0 14812 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[384\]
timestamp 1641350499
transform 1 0 14122 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[383\]
timestamp 1641350499
transform 1 0 13984 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[382\]
timestamp 1641350499
transform 1 0 13846 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[381\]
timestamp 1641350499
transform 1 0 13708 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[380\]
timestamp 1641350499
transform 1 0 13570 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[37\]
timestamp 1641350499
transform 1 0 13386 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[379\]
timestamp 1641350499
transform 1 0 13248 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[378\]
timestamp 1641350499
transform 1 0 13110 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1641350499
transform 1 0 13524 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[377\]
timestamp 1641350499
transform 1 0 12972 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[376\]
timestamp 1641350499
transform 1 0 12834 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[375\]
timestamp 1641350499
transform 1 0 12696 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[374\]
timestamp 1641350499
transform 1 0 12558 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[373\]
timestamp 1641350499
transform 1 0 12420 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[372\]
timestamp 1641350499
transform 1 0 12282 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[371\]
timestamp 1641350499
transform 1 0 12098 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[370\]
timestamp 1641350499
transform 1 0 11960 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1641350499
transform 1 0 12236 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[36\]
timestamp 1641350499
transform 1 0 11822 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[369\]
timestamp 1641350499
transform 1 0 11684 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[368\]
timestamp 1641350499
transform 1 0 11546 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[367\]
timestamp 1641350499
transform 1 0 11408 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[366\]
timestamp 1641350499
transform 1 0 11270 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[365\]
timestamp 1641350499
transform 1 0 11132 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[364\]
timestamp 1641350499
transform 1 0 10994 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[363\]
timestamp 1641350499
transform 1 0 10810 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1641350499
transform 1 0 10948 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[362\]
timestamp 1641350499
transform 1 0 10672 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[361\]
timestamp 1641350499
transform 1 0 10534 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[360\]
timestamp 1641350499
transform 1 0 10396 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[35\]
timestamp 1641350499
transform 1 0 10258 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[359\]
timestamp 1641350499
transform 1 0 10120 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[358\]
timestamp 1641350499
transform 1 0 9982 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[357\]
timestamp 1641350499
transform 1 0 9844 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[356\]
timestamp 1641350499
transform 1 0 9706 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[355\]
timestamp 1641350499
transform 1 0 9522 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1641350499
transform 1 0 9660 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[354\]
timestamp 1641350499
transform 1 0 9384 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[353\]
timestamp 1641350499
transform 1 0 9246 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[352\]
timestamp 1641350499
transform 1 0 9108 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[351\]
timestamp 1641350499
transform 1 0 8970 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[350\]
timestamp 1641350499
transform 1 0 8832 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[34\]
timestamp 1641350499
transform 1 0 8694 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[349\]
timestamp 1641350499
transform 1 0 8556 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[348\]
timestamp 1641350499
transform 1 0 8418 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1641350499
transform 1 0 8372 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1641350499
transform 1 0 8280 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[347\]
timestamp 1641350499
transform 1 0 8142 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[346\]
timestamp 1641350499
transform 1 0 8004 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[345\]
timestamp 1641350499
transform 1 0 7866 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[344\]
timestamp 1641350499
transform 1 0 7728 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[15\]
timestamp 1641350499
transform 1 0 7590 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[13\]
timestamp 1641350499
transform 1 0 7452 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[116\]
timestamp 1641350499
transform 1 0 7314 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[114\]
timestamp 1641350499
transform 1 0 7176 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[119\]
timestamp 1641350499
transform 1 0 6762 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[117\]
timestamp 1641350499
transform 1 0 6900 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[115\]
timestamp 1641350499
transform 1 0 6624 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1641350499
transform 1 0 7084 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_3_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 7130 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_3_139
timestamp 1641350499
transform 1 0 7038 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1641350499
transform 1 0 5980 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[124\]
timestamp 1641350499
transform 1 0 6072 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[123\]
timestamp 1641350499
transform 1 0 6210 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[121\]
timestamp 1641350499
transform 1 0 6486 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[11\]
timestamp 1641350499
transform 1 0 6348 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[129\]
timestamp 1641350499
transform 1 0 5382 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[128\]
timestamp 1641350499
transform 1 0 5520 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[127\]
timestamp 1641350499
transform 1 0 5658 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[120\]
timestamp 1641350499
transform 1 0 5842 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1641350499
transform 1 0 5796 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[131\]
timestamp 1641350499
transform 1 0 5106 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[130\]
timestamp 1641350499
transform 1 0 5244 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[126\]
timestamp 1641350499
transform 1 0 4968 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[118\]
timestamp 1641350499
transform 1 0 4830 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[137\]
timestamp 1641350499
transform 1 0 4232 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[136\]
timestamp 1641350499
transform 1 0 4370 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[135\]
timestamp 1641350499
transform 1 0 4554 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[134\]
timestamp 1641350499
transform 1 0 4692 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1641350499
transform 1 0 4508 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[141\]
timestamp 1641350499
transform 1 0 3680 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[140\]
timestamp 1641350499
transform 1 0 3818 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[138\]
timestamp 1641350499
transform 1 0 4094 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[132\]
timestamp 1641350499
transform 1 0 3956 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1641350499
transform 1 0 3128 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[143\]
timestamp 1641350499
transform 1 0 3404 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[142\]
timestamp 1641350499
transform 1 0 3542 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[122\]
timestamp 1641350499
transform 1 0 3266 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1641350499
transform 1 0 3220 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[148\]
timestamp 1641350499
transform 1 0 2668 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[147\]
timestamp 1641350499
transform 1 0 2806 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[139\]
timestamp 1641350499
transform 1 0 2990 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[133\]
timestamp 1641350499
transform 1 0 2530 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_3_50
timestamp 1641350499
transform 1 0 2944 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1641350499
transform 1 0 2484 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1641350499
transform 1 0 1978 0 -1 1632
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[12\]
timestamp 1641350499
transform 1 0 2346 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[10\]
timestamp 1641350499
transform 1 0 2208 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[104\]
timestamp 1641350499
transform 1 0 2070 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1641350499
transform 1 0 1932 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[153\]
timestamp 1641350499
transform -1 0 1380 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[152\]
timestamp 1641350499
transform -1 0 1518 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[149\]
timestamp 1641350499
transform 1 0 1518 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[146\]
timestamp 1641350499
transform -1 0 1794 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[144\]
timestamp 1641350499
transform 1 0 1794 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1641350499
transform 1 0 782 0 -1 1632
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[160\]
timestamp 1641350499
transform 1 0 1104 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1641350499
transform 1 0 644 0 -1 1632
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1641350499
transform 1 0 1058 0 -1 1632
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_2_722 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 33856 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1641350499
transform -1 0 34408 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_2_730
timestamp 1641350499
transform 1 0 34224 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[97\]
timestamp 1641350499
transform -1 0 33304 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_2_710
timestamp 1641350499
transform 1 0 33304 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_2_695
timestamp 1641350499
transform 1 0 32614 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[95\]
timestamp 1641350499
transform -1 0 33166 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[94\]
timestamp 1641350499
transform -1 0 33028 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[92\]
timestamp 1641350499
transform 1 0 32706 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1641350499
transform 1 0 32844 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_2_681
timestamp 1641350499
transform 1 0 31970 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__conb_1  insts\[90\]
timestamp 1641350499
transform 1 0 32476 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  FILLER_2_689
timestamp 1641350499
transform 1 0 32338 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1641350499
transform 1 0 31418 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1641350499
transform 1 0 30866 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1641350499
transform 1 0 30268 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1641350499
transform 1 0 30314 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1641350499
transform 1 0 30222 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1641350499
transform 1 0 29946 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1641350499
transform 1 0 29394 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1641350499
transform 1 0 28842 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1641350499
transform 1 0 28290 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1641350499
transform 1 0 27370 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1641350499
transform 1 0 27692 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1641350499
transform 1 0 27738 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1641350499
transform 1 0 27646 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1641350499
transform 1 0 26818 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1641350499
transform 1 0 26266 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1641350499
transform 1 0 25714 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1641350499
transform 1 0 25116 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1641350499
transform 1 0 25162 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_526
timestamp 1641350499
transform 1 0 24840 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__decap_12  FILLER_2_514
timestamp 1641350499
transform 1 0 24288 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_502
timestamp 1641350499
transform 1 0 23736 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[453\]
timestamp 1641350499
transform 1 0 24150 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[452\]
timestamp 1641350499
transform 1 0 24012 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[44\]
timestamp 1641350499
transform 1 0 23598 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[449\]
timestamp 1641350499
transform 1 0 23460 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[448\]
timestamp 1641350499
transform 1 0 23322 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[447\]
timestamp 1641350499
transform 1 0 23184 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[446\]
timestamp 1641350499
transform 1 0 23046 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[445\]
timestamp 1641350499
transform 1 0 22908 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[444\]
timestamp 1641350499
transform 1 0 22770 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[443\]
timestamp 1641350499
transform 1 0 22632 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1641350499
transform 1 0 22540 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_2_477
timestamp 1641350499
transform 1 0 22586 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1641350499
transform 1 0 22264 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[43\]
timestamp 1641350499
transform 1 0 22126 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_2_466
timestamp 1641350499
transform 1 0 22080 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_454
timestamp 1641350499
transform 1 0 21528 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[430\]
timestamp 1641350499
transform 1 0 20838 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_2_442
timestamp 1641350499
transform 1 0 20976 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_433
timestamp 1641350499
transform 1 0 20562 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1641350499
transform 1 0 19872 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1641350499
transform 1 0 19964 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1641350499
transform 1 0 20010 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1641350499
transform 1 0 19504 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1641350499
transform 1 0 18952 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_386
timestamp 1641350499
transform 1 0 18400 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1641350499
transform 1 0 17986 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[413\]
timestamp 1641350499
transform 1 0 18262 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1641350499
transform 1 0 17388 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1641350499
transform 1 0 17434 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1641350499
transform 1 0 17342 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1641350499
transform 1 0 17066 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1641350499
transform 1 0 16514 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1641350499
transform 1 0 15962 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1641350499
transform 1 0 15410 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1641350499
transform 1 0 14858 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1641350499
transform 1 0 14306 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1641350499
transform 1 0 14536 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[389\]
timestamp 1641350499
transform 1 0 14398 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1641350499
transform 1 0 14812 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1641350499
transform 1 0 13938 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1641350499
transform 1 0 13386 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1641350499
transform 1 0 12834 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1641350499
transform 1 0 11914 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1641350499
transform 1 0 12236 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1641350499
transform 1 0 12282 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1641350499
transform 1 0 12190 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1641350499
transform 1 0 11362 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1641350499
transform 1 0 10810 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1641350499
transform 1 0 10258 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1641350499
transform 1 0 9660 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1641350499
transform 1 0 9706 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1641350499
transform 1 0 9614 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1641350499
transform 1 0 9338 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1641350499
transform 1 0 8786 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1641350499
transform 1 0 8234 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1641350499
transform 1 0 7682 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1641350499
transform 1 0 6624 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1641350499
transform 1 0 6992 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1641350499
transform 1 0 7084 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1641350499
transform 1 0 7130 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_118
timestamp 1641350499
transform 1 0 6072 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1641350499
transform 1 0 5658 0 1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[125\]
timestamp 1641350499
transform 1 0 5934 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1641350499
transform 1 0 5106 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1641350499
transform 1 0 4508 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1641350499
transform 1 0 4554 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1641350499
transform 1 0 3956 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1641350499
transform 1 0 3036 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[330\]
timestamp 1641350499
transform 1 0 3266 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[145\]
timestamp 1641350499
transform 1 0 3128 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_2_60
timestamp 1641350499
transform 1 0 3404 0 1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[154\]
timestamp 1641350499
transform 1 0 2898 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[150\]
timestamp 1641350499
transform 1 0 2760 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[14\]
timestamp 1641350499
transform 1 0 2622 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[102\]
timestamp 1641350499
transform 1 0 2484 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1641350499
transform 1 0 1978 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[101\]
timestamp 1641350499
transform 1 0 2346 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[100\]
timestamp 1641350499
transform 1 0 2208 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[0\]
timestamp 1641350499
transform 1 0 2070 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1641350499
transform 1 0 1932 0 1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[162\]
timestamp 1641350499
transform 1 0 1242 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[159\]
timestamp 1641350499
transform 1 0 1380 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[157\]
timestamp 1641350499
transform 1 0 1518 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[151\]
timestamp 1641350499
transform -1 0 1794 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[105\]
timestamp 1641350499
transform 1 0 1794 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1641350499
transform 1 0 782 0 1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1641350499
transform 1 0 1150 0 1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1641350499
transform 1 0 644 0 1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_1_729
timestamp 1641350499
transform 1 0 34178 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_0_729
timestamp 1641350499
transform 1 0 34178 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1641350499
transform 1 0 33810 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1641350499
transform 1 0 34132 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1641350499
transform 1 0 34132 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1641350499
transform -1 0 34408 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1641350499
transform -1 0 34408 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1641350499
transform 1 0 33994 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1641350499
transform 1 0 34086 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_709
timestamp 1641350499
transform 1 0 33258 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_713
timestamp 1641350499
transform 1 0 33442 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1641350499
transform 1 0 32844 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_697
timestamp 1641350499
transform 1 0 32706 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_701
timestamp 1641350499
transform 1 0 32890 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1641350499
transform 1 0 32706 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1641350499
transform 1 0 32154 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_685
timestamp 1641350499
transform 1 0 32154 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1641350499
transform 1 0 31556 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1641350499
transform 1 0 31556 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1641350499
transform 1 0 31602 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_673
timestamp 1641350499
transform 1 0 31602 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1641350499
transform 1 0 31418 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1641350499
transform 1 0 31510 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1641350499
transform 1 0 31234 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__decap_12  FILLER_0_657
timestamp 1641350499
transform 1 0 30866 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1641350499
transform 1 0 30268 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1641350499
transform 1 0 30682 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_645
timestamp 1641350499
transform 1 0 30314 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_641
timestamp 1641350499
transform 1 0 30130 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1641350499
transform 1 0 30130 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1641350499
transform 1 0 29578 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1641350499
transform 1 0 29026 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_629
timestamp 1641350499
transform 1 0 29578 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1641350499
transform 1 0 29026 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1641350499
transform 1 0 28658 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1641350499
transform 1 0 28980 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1641350499
transform 1 0 28980 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1641350499
transform 1 0 28842 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1641350499
transform 1 0 28934 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[308\]
timestamp 1641350499
transform 1 0 28152 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[239\]
timestamp 1641350499
transform 1 0 28014 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[175\]
timestamp 1641350499
transform 1 0 27876 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1641350499
transform 1 0 28106 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_0_601
timestamp 1641350499
transform 1 0 28290 0 1 544
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[341\]
timestamp 1641350499
transform 1 0 27554 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[331\]
timestamp 1641350499
transform 1 0 27416 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[307\]
timestamp 1641350499
transform 1 0 27278 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[20\]
timestamp 1641350499
transform 1 0 27738 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1641350499
transform 1 0 27692 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1641350499
transform 1 0 27554 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[249\]
timestamp 1641350499
transform 1 0 27140 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[238\]
timestamp 1641350499
transform 1 0 27002 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[225\]
timestamp 1641350499
transform 1 0 26864 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[1\]
timestamp 1641350499
transform 1 0 26726 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1641350499
transform 1 0 27002 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1641350499
transform 1 0 26450 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1641350499
transform 1 0 26404 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1641350499
transform 1 0 26404 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[184\]
timestamp 1641350499
transform 1 0 26450 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[194\]
timestamp 1641350499
transform 1 0 26588 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_553
timestamp 1641350499
transform 1 0 26082 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1641350499
transform 1 0 26266 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[173\]
timestamp 1641350499
transform 1 0 26266 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[323\]
timestamp 1641350499
transform 1 0 26128 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[337\]
timestamp 1641350499
transform 1 0 26128 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[314\]
timestamp 1641350499
transform 1 0 25990 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[306\]
timestamp 1641350499
transform 1 0 25852 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[301\]
timestamp 1641350499
transform 1 0 25714 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[295\]
timestamp 1641350499
transform 1 0 25576 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1641350499
transform 1 0 25530 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[281\]
timestamp 1641350499
transform 1 0 25438 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[275\]
timestamp 1641350499
transform 1 0 25300 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[265\]
timestamp 1641350499
transform 1 0 25162 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[233\]
timestamp 1641350499
transform 1 0 24978 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1641350499
transform 1 0 25116 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1641350499
transform 1 0 24978 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[21\]
timestamp 1641350499
transform 1 0 24840 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[216\]
timestamp 1641350499
transform 1 0 24702 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[211\]
timestamp 1641350499
transform 1 0 24564 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[207\]
timestamp 1641350499
transform 1 0 24426 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[203\]
timestamp 1641350499
transform 1 0 24288 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1641350499
transform 1 0 24426 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1641350499
transform 1 0 23736 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1641350499
transform 1 0 23736 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[199\]
timestamp 1641350499
transform 1 0 24150 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[191\]
timestamp 1641350499
transform 1 0 24012 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[187\]
timestamp 1641350499
transform 1 0 23874 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1641350499
transform 1 0 23828 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1641350499
transform 1 0 23828 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1641350499
transform 1 0 23874 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[322\]
timestamp 1641350499
transform 1 0 23460 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[180\]
timestamp 1641350499
transform 1 0 23598 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[170\]
timestamp 1641350499
transform 1 0 23322 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[167\]
timestamp 1641350499
transform 1 0 23184 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_490
timestamp 1641350499
transform 1 0 23184 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[32\]
timestamp 1641350499
transform 1 0 23046 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[342\]
timestamp 1641350499
transform 1 0 23046 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 1641350499
transform 1 0 22862 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_1_484
timestamp 1641350499
transform 1 0 22908 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[315\]
timestamp 1641350499
transform 1 0 22908 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[326\]
timestamp 1641350499
transform 1 0 22724 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[333\]
timestamp 1641350499
transform 1 0 22770 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_1_479
timestamp 1641350499
transform 1 0 22678 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1641350499
transform 1 0 22540 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[313\]
timestamp 1641350499
transform 1 0 22586 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_1_471
timestamp 1641350499
transform 1 0 22310 0 -1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1641350499
transform 1 0 22448 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[319\]
timestamp 1641350499
transform 1 0 22172 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[311\]
timestamp 1641350499
transform 1 0 22310 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[309\]
timestamp 1641350499
transform 1 0 22172 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[304\]
timestamp 1641350499
transform 1 0 22034 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1641350499
transform 1 0 22126 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_6  FILLER_1_461
timestamp 1641350499
transform 1 0 21850 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[300\]
timestamp 1641350499
transform 1 0 21896 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[298\]
timestamp 1641350499
transform 1 0 21574 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[294\]
timestamp 1641350499
transform 1 0 21436 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[268\]
timestamp 1641350499
transform 1 0 21758 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_458
timestamp 1641350499
transform 1 0 21712 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1641350499
transform 1 0 21298 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1641350499
transform 1 0 20930 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1641350499
transform 1 0 21206 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1641350499
transform 1 0 21252 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1641350499
transform 1 0 21252 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[287\]
timestamp 1641350499
transform 1 0 21022 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[290\]
timestamp 1641350499
transform 1 0 21298 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1641350499
transform 1 0 21160 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[27\]
timestamp 1641350499
transform 1 0 20746 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[283\]
timestamp 1641350499
transform 1 0 20884 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[276\]
timestamp 1641350499
transform 1 0 20608 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[272\]
timestamp 1641350499
transform 1 0 20470 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[269\]
timestamp 1641350499
transform 1 0 20332 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[261\]
timestamp 1641350499
transform 1 0 20194 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1641350499
transform 1 0 20378 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[259\]
timestamp 1641350499
transform 1 0 19826 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[256\]
timestamp 1641350499
transform 1 0 19688 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[253\]
timestamp 1641350499
transform 1 0 19550 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[232\]
timestamp 1641350499
transform 1 0 20056 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1641350499
transform 1 0 19964 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1641350499
transform 1 0 19826 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1641350499
transform 1 0 20010 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[250\]
timestamp 1641350499
transform 1 0 19412 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[248\]
timestamp 1641350499
transform 1 0 19274 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[245\]
timestamp 1641350499
transform 1 0 19136 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[242\]
timestamp 1641350499
transform 1 0 18998 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1641350499
transform 1 0 19274 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[23\]
timestamp 1641350499
transform 1 0 18860 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[237\]
timestamp 1641350499
transform 1 0 18722 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[234\]
timestamp 1641350499
transform 1 0 18538 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[231\]
timestamp 1641350499
transform 1 0 18400 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1641350499
transform 1 0 18676 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1641350499
transform 1 0 18676 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1641350499
transform 1 0 18722 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1641350499
transform 1 0 18630 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[229\]
timestamp 1641350499
transform 1 0 18262 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[226\]
timestamp 1641350499
transform 1 0 18124 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[223\]
timestamp 1641350499
transform 1 0 17986 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[220\]
timestamp 1641350499
transform 1 0 17848 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1641350499
transform 1 0 18078 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[299\]
timestamp 1641350499
transform 1 0 17250 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[218\]
timestamp 1641350499
transform 1 0 17710 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[215\]
timestamp 1641350499
transform 1 0 17572 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[212\]
timestamp 1641350499
transform 1 0 17434 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1641350499
transform 1 0 17388 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1641350499
transform 1 0 17526 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[24\]
timestamp 1641350499
transform 1 0 17112 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[204\]
timestamp 1641350499
transform 1 0 16974 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[201\]
timestamp 1641350499
transform 1 0 16836 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[19\]
timestamp 1641350499
transform 1 0 16698 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_355
timestamp 1641350499
transform 1 0 16974 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_343
timestamp 1641350499
transform 1 0 16422 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[197\]
timestamp 1641350499
transform 1 0 16560 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[286\]
timestamp 1641350499
transform 1 0 16422 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1641350499
transform 1 0 16054 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1641350499
transform 1 0 16146 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1641350499
transform 1 0 16100 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1641350499
transform 1 0 16100 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[186\]
timestamp 1641350499
transform 1 0 16146 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[189\]
timestamp 1641350499
transform 1 0 16284 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[30\]
timestamp 1641350499
transform 1 0 16284 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1641350499
transform 1 0 16008 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[296\]
timestamp 1641350499
transform 1 0 15732 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[289\]
timestamp 1641350499
transform 1 0 15732 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[279\]
timestamp 1641350499
transform 1 0 15456 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[183\]
timestamp 1641350499
transform 1 0 15870 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[178\]
timestamp 1641350499
transform 1 0 15594 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1641350499
transform 1 0 15870 0 -1 1088
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_1_327
timestamp 1641350499
transform 1 0 15686 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__decap_8  FILLER_1_319
timestamp 1641350499
transform 1 0 15318 0 -1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__conb_1  insts\[227\]
timestamp 1641350499
transform 1 0 15042 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[172\]
timestamp 1641350499
transform 1 0 15318 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[16\]
timestamp 1641350499
transform 1 0 15180 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[164\]
timestamp 1641350499
transform 1 0 14904 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1641350499
transform 1 0 14858 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1641350499
transform 1 0 14720 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[33\]
timestamp 1641350499
transform 1 0 14628 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[334\]
timestamp 1641350499
transform 1 0 14582 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[328\]
timestamp 1641350499
transform 1 0 14306 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[266\]
timestamp 1641350499
transform 1 0 14444 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1641350499
transform 1 0 14812 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_307
timestamp 1641350499
transform 1 0 14766 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_3  FILLER_1_301
timestamp 1641350499
transform 1 0 14490 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1641350499
transform 1 0 14122 0 -1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__conb_1  insts\[324\]
timestamp 1641350499
transform 1 0 13892 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[305\]
timestamp 1641350499
transform 1 0 14168 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[257\]
timestamp 1641350499
transform 1 0 14030 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[251\]
timestamp 1641350499
transform 1 0 13754 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_284
timestamp 1641350499
transform 1 0 13708 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1641350499
transform 1 0 13570 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1641350499
transform 1 0 13202 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1641350499
transform 1 0 13478 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1641350499
transform 1 0 13478 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1641350499
transform 1 0 13524 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1641350499
transform 1 0 13524 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[246\]
timestamp 1641350499
transform 1 0 13570 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[320\]
timestamp 1641350499
transform 1 0 13340 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[240\]
timestamp 1641350499
transform 1 0 13202 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[317\]
timestamp 1641350499
transform 1 0 13064 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1641350499
transform 1 0 12558 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[274\]
timestamp 1641350499
transform 1 0 12512 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[235\]
timestamp 1641350499
transform 1 0 12926 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[22\]
timestamp 1641350499
transform 1 0 12650 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[205\]
timestamp 1641350499
transform 1 0 12788 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1641350499
transform 1 0 12650 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[302\]
timestamp 1641350499
transform 1 0 11960 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[224\]
timestamp 1641350499
transform 1 0 12420 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[219\]
timestamp 1641350499
transform 1 0 12098 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[181\]
timestamp 1641350499
transform 1 0 12282 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1641350499
transform 1 0 12236 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1641350499
transform 1 0 12328 0 -1 1088
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_0_245
timestamp 1641350499
transform 1 0 11914 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[29\]
timestamp 1641350499
transform 1 0 11638 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[252\]
timestamp 1641350499
transform 1 0 11362 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[213\]
timestamp 1641350499
transform 1 0 11776 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[208\]
timestamp 1641350499
transform 1 0 11500 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_242
timestamp 1641350499
transform 1 0 11776 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1641350499
transform 1 0 11224 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[198\]
timestamp 1641350499
transform 1 0 10994 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[202\]
timestamp 1641350499
transform 1 0 11224 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[292\]
timestamp 1641350499
transform 1 0 11086 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_0_228
timestamp 1641350499
transform 1 0 11132 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1641350499
transform 1 0 10994 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1641350499
transform 1 0 10810 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1641350499
transform 1 0 10948 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1641350499
transform 1 0 10948 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[244\]
timestamp 1641350499
transform 1 0 10810 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[338\]
timestamp 1641350499
transform 1 0 10120 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[332\]
timestamp 1641350499
transform 1 0 10120 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[318\]
timestamp 1641350499
transform 1 0 10258 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[285\]
timestamp 1641350499
transform 1 0 10534 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[236\]
timestamp 1641350499
transform 1 0 10396 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[192\]
timestamp 1641350499
transform 1 0 10672 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_209
timestamp 1641350499
transform 1 0 10258 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_8  FILLER_1_196
timestamp 1641350499
transform 1 0 9660 0 -1 1088
box -19 -24 387 296
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1641350499
transform 1 0 10028 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1641350499
transform 1 0 9568 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[278\]
timestamp 1641350499
transform 1 0 9982 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[217\]
timestamp 1641350499
transform 1 0 9706 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[176\]
timestamp 1641350499
transform 1 0 9844 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1641350499
transform 1 0 9660 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[339\]
timestamp 1641350499
transform 1 0 9016 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[270\]
timestamp 1641350499
transform 1 0 9430 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[267\]
timestamp 1641350499
transform 1 0 9154 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[165\]
timestamp 1641350499
transform 1 0 9292 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1641350499
transform 1 0 9108 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[325\]
timestamp 1641350499
transform 1 0 8418 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[263\]
timestamp 1641350499
transform 1 0 8878 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[25\]
timestamp 1641350499
transform 1 0 8602 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[258\]
timestamp 1641350499
transform 1 0 8418 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[190\]
timestamp 1641350499
transform 1 0 8740 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1641350499
transform 1 0 8372 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1641350499
transform 1 0 8372 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1641350499
transform 1 0 8556 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_0_172
timestamp 1641350499
transform 1 0 8556 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1641350499
transform 1 0 8280 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1641350499
transform 1 0 8280 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[316\]
timestamp 1641350499
transform 1 0 8004 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[312\]
timestamp 1641350499
transform 1 0 7866 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[254\]
timestamp 1641350499
transform 1 0 8142 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[264\]
timestamp 1641350499
transform 1 0 7452 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[255\]
timestamp 1641350499
transform 1 0 7728 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[247\]
timestamp 1641350499
transform 1 0 7590 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[188\]
timestamp 1641350499
transform 1 0 7176 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[182\]
timestamp 1641350499
transform 1 0 7314 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1641350499
transform 1 0 7728 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_12  FILLER_1_142
timestamp 1641350499
transform 1 0 7176 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__decap_6  FILLER_1_133
timestamp 1641350499
transform 1 0 6762 0 -1 1088
box -19 -24 295 296
use sky130_fd_sc_hd__conb_1  insts\[303\]
timestamp 1641350499
transform 1 0 7038 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[243\]
timestamp 1641350499
transform 1 0 6900 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[230\]
timestamp 1641350499
transform 1 0 6624 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[200\]
timestamp 1641350499
transform 1 0 6762 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1641350499
transform 1 0 7084 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1641350499
transform 1 0 7130 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1641350499
transform 1 0 7038 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_0_119
timestamp 1641350499
transform 1 0 6118 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[340\]
timestamp 1641350499
transform 1 0 6072 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[310\]
timestamp 1641350499
transform 1 0 6486 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[241\]
timestamp 1641350499
transform 1 0 6348 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[193\]
timestamp 1641350499
transform 1 0 5980 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[163\]
timestamp 1641350499
transform 1 0 6210 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_121
timestamp 1641350499
transform 1 0 6210 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1641350499
transform 1 0 6026 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[273\]
timestamp 1641350499
transform 1 0 5474 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[171\]
timestamp 1641350499
transform 1 0 5612 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[166\]
timestamp 1641350499
transform 1 0 5842 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1641350499
transform 1 0 5796 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_11
timestamp 1641350499
transform 1 0 5796 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1641350499
transform 1 0 5842 0 -1 1088
box -19 -24 203 296
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1641350499
transform 1 0 5612 0 -1 1088
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1641350499
transform 1 0 5750 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1641350499
transform 1 0 4968 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[336\]
timestamp 1641350499
transform 1 0 4922 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[335\]
timestamp 1641350499
transform 1 0 5198 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[293\]
timestamp 1641350499
transform 1 0 5060 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[196\]
timestamp 1641350499
transform 1 0 4830 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[174\]
timestamp 1641350499
transform 1 0 5336 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1641350499
transform 1 0 5060 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1641350499
transform 1 0 4876 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[329\]
timestamp 1641350499
transform 1 0 4232 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[195\]
timestamp 1641350499
transform 1 0 4692 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[179\]
timestamp 1641350499
transform 1 0 4370 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[169\]
timestamp 1641350499
transform 1 0 4554 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1641350499
transform 1 0 4508 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1641350499
transform 1 0 4324 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__conb_1  insts\[282\]
timestamp 1641350499
transform 1 0 3634 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[271\]
timestamp 1641350499
transform 1 0 3772 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[221\]
timestamp 1641350499
transform 1 0 3910 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[168\]
timestamp 1641350499
transform 1 0 4048 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1641350499
transform 1 0 3772 0 -1 1088
box -19 -24 571 296
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1641350499
transform 1 0 4186 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1641350499
transform 1 0 3726 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[26\]
timestamp 1641350499
transform 1 0 3588 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1641350499
transform 1 0 3542 0 -1 1088
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[185\]
timestamp 1641350499
transform 1 0 3450 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[31\]
timestamp 1641350499
transform 1 0 3404 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1641350499
transform 1 0 3266 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1641350499
transform 1 0 3220 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1641350499
transform 1 0 3220 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[177\]
timestamp 1641350499
transform 1 0 3312 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[291\]
timestamp 1641350499
transform 1 0 3266 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1641350499
transform 1 0 3174 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1641350499
transform 1 0 3174 0 -1 1088
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[214\]
timestamp 1641350499
transform 1 0 3036 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[277\]
timestamp 1641350499
transform 1 0 3036 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[262\]
timestamp 1641350499
transform 1 0 2760 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[222\]
timestamp 1641350499
transform 1 0 2898 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[209\]
timestamp 1641350499
transform 1 0 2898 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[206\]
timestamp 1641350499
transform 1 0 2760 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[18\]
timestamp 1641350499
transform 1 0 2622 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[161\]
timestamp 1641350499
transform 1 0 2622 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[112\]
timestamp 1641350499
transform 1 0 2484 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[108\]
timestamp 1641350499
transform 1 0 2484 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1641350499
transform 1 0 1978 0 1 544
box -19 -24 111 296
use sky130_fd_sc_hd__conb_1  insts\[155\]
timestamp 1641350499
transform 1 0 1932 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[111\]
timestamp 1641350499
transform 1 0 2346 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[110\]
timestamp 1641350499
transform 1 0 2208 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[109\]
timestamp 1641350499
transform 1 0 2070 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[107\]
timestamp 1641350499
transform 1 0 2346 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[106\]
timestamp 1641350499
transform 1 0 2208 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[103\]
timestamp 1641350499
transform 1 0 2070 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1641350499
transform 1 0 1932 0 1 544
box -19 -24 65 296
use sky130_fd_sc_hd__conb_1  insts\[113\]
timestamp 1641350499
transform 1 0 1794 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[156\]
timestamp 1641350499
transform 1 0 1794 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[158\]
timestamp 1641350499
transform 1 0 1656 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[17\]
timestamp 1641350499
transform 1 0 1656 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[210\]
timestamp 1641350499
transform 1 0 1518 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[280\]
timestamp 1641350499
transform 1 0 1518 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[228\]
timestamp 1641350499
transform 1 0 1380 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[260\]
timestamp 1641350499
transform 1 0 1242 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[284\]
timestamp 1641350499
transform 1 0 1380 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[28\]
timestamp 1641350499
transform -1 0 1380 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[327\]
timestamp 1641350499
transform -1 0 1104 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[321\]
timestamp 1641350499
transform 1 0 1104 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[2\]
timestamp 1641350499
transform -1 0 966 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[297\]
timestamp 1641350499
transform -1 0 1104 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__conb_1  insts\[288\]
timestamp 1641350499
transform -1 0 1242 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1641350499
transform 1 0 644 0 -1 1088
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1641350499
transform 1 0 644 0 1 544
box -19 -24 157 296
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1641350499
transform 1 0 782 0 -1 1088
box -19 -24 203 296
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp 1641350499
transform 1 0 782 0 1 544
box -19 -24 65 296
<< labels >>
rlabel metal3 s 0 1908 300 1968 6 HI[0]
port 0 nsew signal tristate
rlabel metal3 s 0 1772 300 1832 6 HI[100]
port 1 nsew signal tristate
rlabel metal3 s 0 1636 300 1696 6 HI[101]
port 2 nsew signal tristate
rlabel metal3 s 0 1500 300 1560 6 HI[102]
port 3 nsew signal tristate
rlabel metal3 s 0 1364 300 1424 6 HI[103]
port 4 nsew signal tristate
rlabel metal3 s 0 1228 300 1288 6 HI[104]
port 5 nsew signal tristate
rlabel metal3 s 0 1092 300 1152 6 HI[105]
port 6 nsew signal tristate
rlabel metal3 s 0 956 300 1016 6 HI[106]
port 7 nsew signal tristate
rlabel metal3 s 0 820 300 880 6 HI[107]
port 8 nsew signal tristate
rlabel metal3 s 0 684 300 744 6 HI[108]
port 9 nsew signal tristate
rlabel metal3 s 0 548 300 608 6 HI[109]
port 10 nsew signal tristate
rlabel metal3 s 0 2044 300 2104 6 HI[10]
port 11 nsew signal tristate
rlabel metal3 s 0 412 300 472 6 HI[110]
port 12 nsew signal tristate
rlabel metal3 s 0 140 300 200 6 HI[111]
port 13 nsew signal tristate
rlabel metal3 s 0 4 300 64 6 HI[112]
port 14 nsew signal tristate
rlabel metal3 s 0 276 300 336 6 HI[113]
port 15 nsew signal tristate
rlabel metal2 s 7047 1900 7075 2200 6 HI[114]
port 16 nsew signal tristate
rlabel metal2 s 6495 1900 6523 2200 6 HI[115]
port 17 nsew signal tristate
rlabel metal2 s 6909 1900 6937 2200 6 HI[116]
port 18 nsew signal tristate
rlabel metal2 s 6771 1900 6799 2200 6 HI[117]
port 19 nsew signal tristate
rlabel metal2 s 4701 1900 4729 2200 6 HI[118]
port 20 nsew signal tristate
rlabel metal2 s 6633 1900 6661 2200 6 HI[119]
port 21 nsew signal tristate
rlabel metal2 s 6219 1900 6247 2200 6 HI[11]
port 22 nsew signal tristate
rlabel metal2 s 5667 1900 5695 2200 6 HI[120]
port 23 nsew signal tristate
rlabel metal2 s 6357 1900 6385 2200 6 HI[121]
port 24 nsew signal tristate
rlabel metal2 s 3183 1900 3211 2200 6 HI[122]
port 25 nsew signal tristate
rlabel metal2 s 6081 1900 6109 2200 6 HI[123]
port 26 nsew signal tristate
rlabel metal2 s 5943 1900 5971 2200 6 HI[124]
port 27 nsew signal tristate
rlabel metal2 s 5805 1900 5833 2200 6 HI[125]
port 28 nsew signal tristate
rlabel metal2 s 4839 1900 4867 2200 6 HI[126]
port 29 nsew signal tristate
rlabel metal2 s 5529 1900 5557 2200 6 HI[127]
port 30 nsew signal tristate
rlabel metal2 s 5391 1900 5419 2200 6 HI[128]
port 31 nsew signal tristate
rlabel metal2 s 5253 1900 5281 2200 6 HI[129]
port 32 nsew signal tristate
rlabel metal2 s 285 1900 313 2200 6 HI[12]
port 33 nsew signal tristate
rlabel metal2 s 5115 1900 5143 2200 6 HI[130]
port 34 nsew signal tristate
rlabel metal2 s 4977 1900 5005 2200 6 HI[131]
port 35 nsew signal tristate
rlabel metal2 s 3873 1900 3901 2200 6 HI[132]
port 36 nsew signal tristate
rlabel metal2 s 2493 1900 2521 2200 6 HI[133]
port 37 nsew signal tristate
rlabel metal2 s 4563 1900 4591 2200 6 HI[134]
port 38 nsew signal tristate
rlabel metal2 s 4425 1900 4453 2200 6 HI[135]
port 39 nsew signal tristate
rlabel metal2 s 4287 1900 4315 2200 6 HI[136]
port 40 nsew signal tristate
rlabel metal2 s 4149 1900 4177 2200 6 HI[137]
port 41 nsew signal tristate
rlabel metal2 s 4011 1900 4039 2200 6 HI[138]
port 42 nsew signal tristate
rlabel metal2 s 2907 1900 2935 2200 6 HI[139]
port 43 nsew signal tristate
rlabel metal2 s 7185 1900 7213 2200 6 HI[13]
port 44 nsew signal tristate
rlabel metal2 s 3735 1900 3763 2200 6 HI[140]
port 45 nsew signal tristate
rlabel metal2 s 3597 1900 3625 2200 6 HI[141]
port 46 nsew signal tristate
rlabel metal2 s 3459 1900 3487 2200 6 HI[142]
port 47 nsew signal tristate
rlabel metal2 s 3321 1900 3349 2200 6 HI[143]
port 48 nsew signal tristate
rlabel metal2 s 9 1900 37 2200 6 HI[144]
port 49 nsew signal tristate
rlabel metal2 s 3045 1900 3073 2200 6 HI[145]
port 50 nsew signal tristate
rlabel metal2 s 1803 1900 1831 2200 6 HI[146]
port 51 nsew signal tristate
rlabel metal2 s 2769 1900 2797 2200 6 HI[147]
port 52 nsew signal tristate
rlabel metal2 s 2631 1900 2659 2200 6 HI[148]
port 53 nsew signal tristate
rlabel metal2 s 147 1900 175 2200 6 HI[149]
port 54 nsew signal tristate
rlabel metal2 s 2217 1900 2245 2200 6 HI[14]
port 55 nsew signal tristate
rlabel metal2 s 2355 1900 2383 2200 6 HI[150]
port 56 nsew signal tristate
rlabel metal2 s 1941 1900 1969 2200 6 HI[151]
port 57 nsew signal tristate
rlabel metal2 s 2079 1900 2107 2200 6 HI[152]
port 58 nsew signal tristate
rlabel metal2 s 1665 1900 1693 2200 6 HI[153]
port 59 nsew signal tristate
rlabel metal2 s 561 1900 589 2200 6 HI[154]
port 60 nsew signal tristate
rlabel metal2 s 1527 1900 1555 2200 6 HI[155]
port 61 nsew signal tristate
rlabel metal2 s 1389 1900 1417 2200 6 HI[156]
port 62 nsew signal tristate
rlabel metal2 s 1251 1900 1279 2200 6 HI[157]
port 63 nsew signal tristate
rlabel metal2 s 1113 1900 1141 2200 6 HI[158]
port 64 nsew signal tristate
rlabel metal2 s 975 1900 1003 2200 6 HI[159]
port 65 nsew signal tristate
rlabel metal2 s 7323 1900 7351 2200 6 HI[15]
port 66 nsew signal tristate
rlabel metal2 s 699 1900 727 2200 6 HI[160]
port 67 nsew signal tristate
rlabel metal2 s 837 1900 865 2200 6 HI[161]
port 68 nsew signal tristate
rlabel metal2 s 423 1900 451 2200 6 HI[162]
port 69 nsew signal tristate
rlabel metal2 s 5943 0 5971 300 6 HI[163]
port 70 nsew signal tristate
rlabel metal2 s 14499 0 14527 300 6 HI[164]
port 71 nsew signal tristate
rlabel metal2 s 8979 0 9007 300 6 HI[165]
port 72 nsew signal tristate
rlabel metal2 s 5529 0 5557 300 6 HI[166]
port 73 nsew signal tristate
rlabel metal2 s 22641 0 22669 300 6 HI[167]
port 74 nsew signal tristate
rlabel metal2 s 3873 0 3901 300 6 HI[168]
port 75 nsew signal tristate
rlabel metal2 s 4287 0 4315 300 6 HI[169]
port 76 nsew signal tristate
rlabel metal2 s 14775 0 14803 300 6 HI[16]
port 77 nsew signal tristate
rlabel metal2 s 22779 0 22807 300 6 HI[170]
port 78 nsew signal tristate
rlabel metal2 s 5391 0 5419 300 6 HI[171]
port 79 nsew signal tristate
rlabel metal2 s 14913 0 14941 300 6 HI[172]
port 80 nsew signal tristate
rlabel metal2 s 25677 0 25705 300 6 HI[173]
port 81 nsew signal tristate
rlabel metal2 s 5115 0 5143 300 6 HI[174]
port 82 nsew signal tristate
rlabel metal2 s 27333 0 27361 300 6 HI[175]
port 83 nsew signal tristate
rlabel metal2 s 9531 0 9559 300 6 HI[176]
port 84 nsew signal tristate
rlabel metal2 s 3183 0 3211 300 6 HI[177]
port 85 nsew signal tristate
rlabel metal2 s 15189 0 15217 300 6 HI[178]
port 86 nsew signal tristate
rlabel metal2 s 4149 0 4177 300 6 HI[179]
port 87 nsew signal tristate
rlabel metal2 s 147 0 175 300 6 HI[17]
port 88 nsew signal tristate
rlabel metal2 s 23055 0 23083 300 6 HI[180]
port 89 nsew signal tristate
rlabel metal2 s 11877 0 11905 300 6 HI[181]
port 90 nsew signal tristate
rlabel metal2 s 7047 0 7075 300 6 HI[182]
port 91 nsew signal tristate
rlabel metal2 s 15465 0 15493 300 6 HI[183]
port 92 nsew signal tristate
rlabel metal2 s 25815 0 25843 300 6 HI[184]
port 93 nsew signal tristate
rlabel metal2 s 3045 0 3073 300 6 HI[185]
port 94 nsew signal tristate
rlabel metal2 s 15603 0 15631 300 6 HI[186]
port 95 nsew signal tristate
rlabel metal2 s 23193 0 23221 300 6 HI[187]
port 96 nsew signal tristate
rlabel metal2 s 6909 0 6937 300 6 HI[188]
port 97 nsew signal tristate
rlabel metal2 s 15741 0 15769 300 6 HI[189]
port 98 nsew signal tristate
rlabel metal2 s 1389 0 1417 300 6 HI[18]
port 99 nsew signal tristate
rlabel metal2 s 8427 0 8455 300 6 HI[190]
port 100 nsew signal tristate
rlabel metal2 s 23331 0 23359 300 6 HI[191]
port 101 nsew signal tristate
rlabel metal2 s 10359 0 10387 300 6 HI[192]
port 102 nsew signal tristate
rlabel metal2 s 5667 0 5695 300 6 HI[193]
port 103 nsew signal tristate
rlabel metal2 s 25953 0 25981 300 6 HI[194]
port 104 nsew signal tristate
rlabel metal2 s 4425 0 4453 300 6 HI[195]
port 105 nsew signal tristate
rlabel metal2 s 4563 0 4591 300 6 HI[196]
port 106 nsew signal tristate
rlabel metal2 s 16155 0 16183 300 6 HI[197]
port 107 nsew signal tristate
rlabel metal2 s 10635 0 10663 300 6 HI[198]
port 108 nsew signal tristate
rlabel metal2 s 23469 0 23497 300 6 HI[199]
port 109 nsew signal tristate
rlabel metal2 s 16293 0 16321 300 6 HI[19]
port 110 nsew signal tristate
rlabel metal2 s 26091 0 26119 300 6 HI[1]
port 111 nsew signal tristate
rlabel metal2 s 6495 0 6523 300 6 HI[200]
port 112 nsew signal tristate
rlabel metal2 s 16431 0 16459 300 6 HI[201]
port 113 nsew signal tristate
rlabel metal2 s 10911 0 10939 300 6 HI[202]
port 114 nsew signal tristate
rlabel metal2 s 23607 0 23635 300 6 HI[203]
port 115 nsew signal tristate
rlabel metal2 s 16569 0 16597 300 6 HI[204]
port 116 nsew signal tristate
rlabel metal2 s 12429 0 12457 300 6 HI[205]
port 117 nsew signal tristate
rlabel metal2 s 2493 0 2521 300 6 HI[206]
port 118 nsew signal tristate
rlabel metal2 s 23745 0 23773 300 6 HI[207]
port 119 nsew signal tristate
rlabel metal2 s 11187 0 11215 300 6 HI[208]
port 120 nsew signal tristate
rlabel metal2 s 423 0 451 300 6 HI[209]
port 121 nsew signal tristate
rlabel metal2 s 27057 0 27085 300 6 HI[20]
port 122 nsew signal tristate
rlabel metal2 s 1113 0 1141 300 6 HI[210]
port 123 nsew signal tristate
rlabel metal2 s 23883 0 23911 300 6 HI[211]
port 124 nsew signal tristate
rlabel metal2 s 16983 0 17011 300 6 HI[212]
port 125 nsew signal tristate
rlabel metal2 s 11463 0 11491 300 6 HI[213]
port 126 nsew signal tristate
rlabel metal2 s 2217 0 2245 300 6 HI[214]
port 127 nsew signal tristate
rlabel metal2 s 17121 0 17149 300 6 HI[215]
port 128 nsew signal tristate
rlabel metal2 s 24021 0 24049 300 6 HI[216]
port 129 nsew signal tristate
rlabel metal2 s 9255 0 9283 300 6 HI[217]
port 130 nsew signal tristate
rlabel metal2 s 17259 0 17287 300 6 HI[218]
port 131 nsew signal tristate
rlabel metal2 s 11739 0 11767 300 6 HI[219]
port 132 nsew signal tristate
rlabel metal2 s 24159 0 24187 300 6 HI[21]
port 133 nsew signal tristate
rlabel metal2 s 17397 0 17425 300 6 HI[220]
port 134 nsew signal tristate
rlabel metal2 s 3735 0 3763 300 6 HI[221]
port 135 nsew signal tristate
rlabel metal2 s 2769 0 2797 300 6 HI[222]
port 136 nsew signal tristate
rlabel metal2 s 17535 0 17563 300 6 HI[223]
port 137 nsew signal tristate
rlabel metal2 s 12015 0 12043 300 6 HI[224]
port 138 nsew signal tristate
rlabel metal2 s 26229 0 26257 300 6 HI[225]
port 139 nsew signal tristate
rlabel metal2 s 17673 0 17701 300 6 HI[226]
port 140 nsew signal tristate
rlabel metal2 s 14361 0 14389 300 6 HI[227]
port 141 nsew signal tristate
rlabel metal2 s 9 0 37 300 6 HI[228]
port 142 nsew signal tristate
rlabel metal2 s 17811 0 17839 300 6 HI[229]
port 143 nsew signal tristate
rlabel metal2 s 12291 0 12319 300 6 HI[22]
port 144 nsew signal tristate
rlabel metal2 s 6357 0 6385 300 6 HI[230]
port 145 nsew signal tristate
rlabel metal2 s 17949 0 17977 300 6 HI[231]
port 146 nsew signal tristate
rlabel metal2 s 19605 0 19633 300 6 HI[232]
port 147 nsew signal tristate
rlabel metal2 s 24297 0 24325 300 6 HI[233]
port 148 nsew signal tristate
rlabel metal2 s 18087 0 18115 300 6 HI[234]
port 149 nsew signal tristate
rlabel metal2 s 12567 0 12595 300 6 HI[235]
port 150 nsew signal tristate
rlabel metal2 s 10083 0 10111 300 6 HI[236]
port 151 nsew signal tristate
rlabel metal2 s 18225 0 18253 300 6 HI[237]
port 152 nsew signal tristate
rlabel metal2 s 26367 0 26395 300 6 HI[238]
port 153 nsew signal tristate
rlabel metal2 s 27471 0 27499 300 6 HI[239]
port 154 nsew signal tristate
rlabel metal2 s 18363 0 18391 300 6 HI[23]
port 155 nsew signal tristate
rlabel metal2 s 12843 0 12871 300 6 HI[240]
port 156 nsew signal tristate
rlabel metal2 s 6081 0 6109 300 6 HI[241]
port 157 nsew signal tristate
rlabel metal2 s 18501 0 18529 300 6 HI[242]
port 158 nsew signal tristate
rlabel metal2 s 6633 0 6661 300 6 HI[243]
port 159 nsew signal tristate
rlabel metal2 s 10497 0 10525 300 6 HI[244]
port 160 nsew signal tristate
rlabel metal2 s 18639 0 18667 300 6 HI[245]
port 161 nsew signal tristate
rlabel metal2 s 13119 0 13147 300 6 HI[246]
port 162 nsew signal tristate
rlabel metal2 s 7323 0 7351 300 6 HI[247]
port 163 nsew signal tristate
rlabel metal2 s 18777 0 18805 300 6 HI[248]
port 164 nsew signal tristate
rlabel metal2 s 26505 0 26533 300 6 HI[249]
port 165 nsew signal tristate
rlabel metal2 s 16707 0 16735 300 6 HI[24]
port 166 nsew signal tristate
rlabel metal2 s 18915 0 18943 300 6 HI[250]
port 167 nsew signal tristate
rlabel metal2 s 13395 0 13423 300 6 HI[251]
port 168 nsew signal tristate
rlabel metal2 s 11049 0 11077 300 6 HI[252]
port 169 nsew signal tristate
rlabel metal2 s 19053 0 19081 300 6 HI[253]
port 170 nsew signal tristate
rlabel metal2 s 7875 0 7903 300 6 HI[254]
port 171 nsew signal tristate
rlabel metal2 s 7461 0 7489 300 6 HI[255]
port 172 nsew signal tristate
rlabel metal2 s 19191 0 19219 300 6 HI[256]
port 173 nsew signal tristate
rlabel metal2 s 13671 0 13699 300 6 HI[257]
port 174 nsew signal tristate
rlabel metal2 s 8151 0 8179 300 6 HI[258]
port 175 nsew signal tristate
rlabel metal2 s 19329 0 19357 300 6 HI[259]
port 176 nsew signal tristate
rlabel metal2 s 8289 0 8317 300 6 HI[25]
port 177 nsew signal tristate
rlabel metal2 s 975 0 1003 300 6 HI[260]
port 178 nsew signal tristate
rlabel metal2 s 19467 0 19495 300 6 HI[261]
port 179 nsew signal tristate
rlabel metal2 s 837 0 865 300 6 HI[262]
port 180 nsew signal tristate
rlabel metal2 s 8565 0 8593 300 6 HI[263]
port 181 nsew signal tristate
rlabel metal2 s 7185 0 7213 300 6 HI[264]
port 182 nsew signal tristate
rlabel metal2 s 24435 0 24463 300 6 HI[265]
port 183 nsew signal tristate
rlabel metal2 s 14085 0 14113 300 6 HI[266]
port 184 nsew signal tristate
rlabel metal2 s 8841 0 8869 300 6 HI[267]
port 185 nsew signal tristate
rlabel metal2 s 21261 0 21289 300 6 HI[268]
port 186 nsew signal tristate
rlabel metal2 s 19743 0 19771 300 6 HI[269]
port 187 nsew signal tristate
rlabel metal2 s 3321 0 3349 300 6 HI[26]
port 188 nsew signal tristate
rlabel metal2 s 9117 0 9145 300 6 HI[270]
port 189 nsew signal tristate
rlabel metal2 s 3597 0 3625 300 6 HI[271]
port 190 nsew signal tristate
rlabel metal2 s 19881 0 19909 300 6 HI[272]
port 191 nsew signal tristate
rlabel metal2 s 5253 0 5281 300 6 HI[273]
port 192 nsew signal tristate
rlabel metal2 s 12153 0 12181 300 6 HI[274]
port 193 nsew signal tristate
rlabel metal2 s 24573 0 24601 300 6 HI[275]
port 194 nsew signal tristate
rlabel metal2 s 20019 0 20047 300 6 HI[276]
port 195 nsew signal tristate
rlabel metal2 s 2631 0 2659 300 6 HI[277]
port 196 nsew signal tristate
rlabel metal2 s 9669 0 9697 300 6 HI[278]
port 197 nsew signal tristate
rlabel metal2 s 14637 0 14665 300 6 HI[279]
port 198 nsew signal tristate
rlabel metal2 s 20157 0 20185 300 6 HI[27]
port 199 nsew signal tristate
rlabel metal2 s 1527 0 1555 300 6 HI[280]
port 200 nsew signal tristate
rlabel metal2 s 24711 0 24739 300 6 HI[281]
port 201 nsew signal tristate
rlabel metal2 s 3459 0 3487 300 6 HI[282]
port 202 nsew signal tristate
rlabel metal2 s 20295 0 20323 300 6 HI[283]
port 203 nsew signal tristate
rlabel metal2 s 699 0 727 300 6 HI[284]
port 204 nsew signal tristate
rlabel metal2 s 10221 0 10249 300 6 HI[285]
port 205 nsew signal tristate
rlabel metal2 s 16017 0 16045 300 6 HI[286]
port 206 nsew signal tristate
rlabel metal2 s 20433 0 20461 300 6 HI[287]
port 207 nsew signal tristate
rlabel metal2 s 1665 0 1693 300 6 HI[288]
port 208 nsew signal tristate
rlabel metal2 s 15051 0 15079 300 6 HI[289]
port 209 nsew signal tristate
rlabel metal2 s 1941 0 1969 300 6 HI[28]
port 210 nsew signal tristate
rlabel metal2 s 20571 0 20599 300 6 HI[290]
port 211 nsew signal tristate
rlabel metal2 s 2355 0 2383 300 6 HI[291]
port 212 nsew signal tristate
rlabel metal2 s 10773 0 10801 300 6 HI[292]
port 213 nsew signal tristate
rlabel metal2 s 4839 0 4867 300 6 HI[293]
port 214 nsew signal tristate
rlabel metal2 s 20709 0 20737 300 6 HI[294]
port 215 nsew signal tristate
rlabel metal2 s 24849 0 24877 300 6 HI[295]
port 216 nsew signal tristate
rlabel metal2 s 15327 0 15355 300 6 HI[296]
port 217 nsew signal tristate
rlabel metal2 s 1251 0 1279 300 6 HI[297]
port 218 nsew signal tristate
rlabel metal2 s 20847 0 20875 300 6 HI[298]
port 219 nsew signal tristate
rlabel metal2 s 16845 0 16873 300 6 HI[299]
port 220 nsew signal tristate
rlabel metal2 s 11325 0 11353 300 6 HI[29]
port 221 nsew signal tristate
rlabel metal2 s 2079 0 2107 300 6 HI[2]
port 222 nsew signal tristate
rlabel metal2 s 20985 0 21013 300 6 HI[300]
port 223 nsew signal tristate
rlabel metal2 s 24987 0 25015 300 6 HI[301]
port 224 nsew signal tristate
rlabel metal2 s 11601 0 11629 300 6 HI[302]
port 225 nsew signal tristate
rlabel metal2 s 6771 0 6799 300 6 HI[303]
port 226 nsew signal tristate
rlabel metal2 s 21123 0 21151 300 6 HI[304]
port 227 nsew signal tristate
rlabel metal2 s 13809 0 13837 300 6 HI[305]
port 228 nsew signal tristate
rlabel metal2 s 25125 0 25153 300 6 HI[306]
port 229 nsew signal tristate
rlabel metal2 s 26643 0 26671 300 6 HI[307]
port 230 nsew signal tristate
rlabel metal2 s 27195 0 27223 300 6 HI[308]
port 231 nsew signal tristate
rlabel metal2 s 21537 0 21565 300 6 HI[309]
port 232 nsew signal tristate
rlabel metal2 s 15879 0 15907 300 6 HI[30]
port 233 nsew signal tristate
rlabel metal2 s 6219 0 6247 300 6 HI[310]
port 234 nsew signal tristate
rlabel metal2 s 21399 0 21427 300 6 HI[311]
port 235 nsew signal tristate
rlabel metal2 s 7599 0 7627 300 6 HI[312]
port 236 nsew signal tristate
rlabel metal2 s 21813 0 21841 300 6 HI[313]
port 237 nsew signal tristate
rlabel metal2 s 25263 0 25291 300 6 HI[314]
port 238 nsew signal tristate
rlabel metal2 s 22365 0 22393 300 6 HI[315]
port 239 nsew signal tristate
rlabel metal2 s 7737 0 7765 300 6 HI[316]
port 240 nsew signal tristate
rlabel metal2 s 12705 0 12733 300 6 HI[317]
port 241 nsew signal tristate
rlabel metal2 s 9945 0 9973 300 6 HI[318]
port 242 nsew signal tristate
rlabel metal2 s 21675 0 21703 300 6 HI[319]
port 243 nsew signal tristate
rlabel metal2 s 285 0 313 300 6 HI[31]
port 244 nsew signal tristate
rlabel metal2 s 12981 0 13009 300 6 HI[320]
port 245 nsew signal tristate
rlabel metal2 s 561 0 589 300 6 HI[321]
port 246 nsew signal tristate
rlabel metal2 s 22917 0 22945 300 6 HI[322]
port 247 nsew signal tristate
rlabel metal2 s 25401 0 25429 300 6 HI[323]
port 248 nsew signal tristate
rlabel metal2 s 13257 0 13285 300 6 HI[324]
port 249 nsew signal tristate
rlabel metal2 s 8013 0 8041 300 6 HI[325]
port 250 nsew signal tristate
rlabel metal2 s 21951 0 21979 300 6 HI[326]
port 251 nsew signal tristate
rlabel metal2 s 1803 0 1831 300 6 HI[327]
port 252 nsew signal tristate
rlabel metal2 s 13533 0 13561 300 6 HI[328]
port 253 nsew signal tristate
rlabel metal2 s 4011 0 4039 300 6 HI[329]
port 254 nsew signal tristate
rlabel metal2 s 22089 0 22117 300 6 HI[32]
port 255 nsew signal tristate
rlabel metal2 s 2907 0 2935 300 6 HI[330]
port 256 nsew signal tristate
rlabel metal2 s 26781 0 26809 300 6 HI[331]
port 257 nsew signal tristate
rlabel metal2 s 9393 0 9421 300 6 HI[332]
port 258 nsew signal tristate
rlabel metal2 s 22227 0 22255 300 6 HI[333]
port 259 nsew signal tristate
rlabel metal2 s 13947 0 13975 300 6 HI[334]
port 260 nsew signal tristate
rlabel metal2 s 4977 0 5005 300 6 HI[335]
port 261 nsew signal tristate
rlabel metal2 s 4701 0 4729 300 6 HI[336]
port 262 nsew signal tristate
rlabel metal2 s 25539 0 25567 300 6 HI[337]
port 263 nsew signal tristate
rlabel metal2 s 9807 0 9835 300 6 HI[338]
port 264 nsew signal tristate
rlabel metal2 s 8703 0 8731 300 6 HI[339]
port 265 nsew signal tristate
rlabel metal2 s 14223 0 14251 300 6 HI[33]
port 266 nsew signal tristate
rlabel metal2 s 5805 0 5833 300 6 HI[340]
port 267 nsew signal tristate
rlabel metal2 s 26919 0 26947 300 6 HI[341]
port 268 nsew signal tristate
rlabel metal2 s 22503 0 22531 300 6 HI[342]
port 269 nsew signal tristate
rlabel metal2 s 33957 1900 33985 2200 6 HI[343]
port 270 nsew signal tristate
rlabel metal2 s 7461 1900 7489 2200 6 HI[344]
port 271 nsew signal tristate
rlabel metal2 s 7599 1900 7627 2200 6 HI[345]
port 272 nsew signal tristate
rlabel metal2 s 7737 1900 7765 2200 6 HI[346]
port 273 nsew signal tristate
rlabel metal2 s 7875 1900 7903 2200 6 HI[347]
port 274 nsew signal tristate
rlabel metal2 s 8013 1900 8041 2200 6 HI[348]
port 275 nsew signal tristate
rlabel metal2 s 8151 1900 8179 2200 6 HI[349]
port 276 nsew signal tristate
rlabel metal2 s 8289 1900 8317 2200 6 HI[34]
port 277 nsew signal tristate
rlabel metal2 s 8427 1900 8455 2200 6 HI[350]
port 278 nsew signal tristate
rlabel metal2 s 8565 1900 8593 2200 6 HI[351]
port 279 nsew signal tristate
rlabel metal2 s 8703 1900 8731 2200 6 HI[352]
port 280 nsew signal tristate
rlabel metal2 s 8841 1900 8869 2200 6 HI[353]
port 281 nsew signal tristate
rlabel metal2 s 8979 1900 9007 2200 6 HI[354]
port 282 nsew signal tristate
rlabel metal2 s 9117 1900 9145 2200 6 HI[355]
port 283 nsew signal tristate
rlabel metal2 s 9255 1900 9283 2200 6 HI[356]
port 284 nsew signal tristate
rlabel metal2 s 9393 1900 9421 2200 6 HI[357]
port 285 nsew signal tristate
rlabel metal2 s 9531 1900 9559 2200 6 HI[358]
port 286 nsew signal tristate
rlabel metal2 s 9669 1900 9697 2200 6 HI[359]
port 287 nsew signal tristate
rlabel metal2 s 9807 1900 9835 2200 6 HI[35]
port 288 nsew signal tristate
rlabel metal2 s 9945 1900 9973 2200 6 HI[360]
port 289 nsew signal tristate
rlabel metal2 s 10083 1900 10111 2200 6 HI[361]
port 290 nsew signal tristate
rlabel metal2 s 10221 1900 10249 2200 6 HI[362]
port 291 nsew signal tristate
rlabel metal2 s 10359 1900 10387 2200 6 HI[363]
port 292 nsew signal tristate
rlabel metal2 s 10497 1900 10525 2200 6 HI[364]
port 293 nsew signal tristate
rlabel metal2 s 10635 1900 10663 2200 6 HI[365]
port 294 nsew signal tristate
rlabel metal2 s 10773 1900 10801 2200 6 HI[366]
port 295 nsew signal tristate
rlabel metal2 s 10911 1900 10939 2200 6 HI[367]
port 296 nsew signal tristate
rlabel metal2 s 11049 1900 11077 2200 6 HI[368]
port 297 nsew signal tristate
rlabel metal2 s 11187 1900 11215 2200 6 HI[369]
port 298 nsew signal tristate
rlabel metal2 s 11325 1900 11353 2200 6 HI[36]
port 299 nsew signal tristate
rlabel metal2 s 11463 1900 11491 2200 6 HI[370]
port 300 nsew signal tristate
rlabel metal2 s 11601 1900 11629 2200 6 HI[371]
port 301 nsew signal tristate
rlabel metal2 s 11739 1900 11767 2200 6 HI[372]
port 302 nsew signal tristate
rlabel metal2 s 11877 1900 11905 2200 6 HI[373]
port 303 nsew signal tristate
rlabel metal2 s 12015 1900 12043 2200 6 HI[374]
port 304 nsew signal tristate
rlabel metal2 s 12153 1900 12181 2200 6 HI[375]
port 305 nsew signal tristate
rlabel metal2 s 12291 1900 12319 2200 6 HI[376]
port 306 nsew signal tristate
rlabel metal2 s 12429 1900 12457 2200 6 HI[377]
port 307 nsew signal tristate
rlabel metal2 s 12567 1900 12595 2200 6 HI[378]
port 308 nsew signal tristate
rlabel metal2 s 12705 1900 12733 2200 6 HI[379]
port 309 nsew signal tristate
rlabel metal2 s 12843 1900 12871 2200 6 HI[37]
port 310 nsew signal tristate
rlabel metal2 s 12981 1900 13009 2200 6 HI[380]
port 311 nsew signal tristate
rlabel metal2 s 13119 1900 13147 2200 6 HI[381]
port 312 nsew signal tristate
rlabel metal2 s 13257 1900 13285 2200 6 HI[382]
port 313 nsew signal tristate
rlabel metal2 s 13395 1900 13423 2200 6 HI[383]
port 314 nsew signal tristate
rlabel metal2 s 13533 1900 13561 2200 6 HI[384]
port 315 nsew signal tristate
rlabel metal2 s 13671 1900 13699 2200 6 HI[385]
port 316 nsew signal tristate
rlabel metal2 s 13809 1900 13837 2200 6 HI[386]
port 317 nsew signal tristate
rlabel metal2 s 13947 1900 13975 2200 6 HI[387]
port 318 nsew signal tristate
rlabel metal2 s 14085 1900 14113 2200 6 HI[388]
port 319 nsew signal tristate
rlabel metal2 s 14223 1900 14251 2200 6 HI[389]
port 320 nsew signal tristate
rlabel metal2 s 14361 1900 14389 2200 6 HI[38]
port 321 nsew signal tristate
rlabel metal2 s 14499 1900 14527 2200 6 HI[390]
port 322 nsew signal tristate
rlabel metal2 s 14637 1900 14665 2200 6 HI[391]
port 323 nsew signal tristate
rlabel metal2 s 14775 1900 14803 2200 6 HI[392]
port 324 nsew signal tristate
rlabel metal2 s 14913 1900 14941 2200 6 HI[393]
port 325 nsew signal tristate
rlabel metal2 s 15051 1900 15079 2200 6 HI[394]
port 326 nsew signal tristate
rlabel metal2 s 15189 1900 15217 2200 6 HI[395]
port 327 nsew signal tristate
rlabel metal2 s 15327 1900 15355 2200 6 HI[396]
port 328 nsew signal tristate
rlabel metal2 s 15465 1900 15493 2200 6 HI[397]
port 329 nsew signal tristate
rlabel metal2 s 15603 1900 15631 2200 6 HI[398]
port 330 nsew signal tristate
rlabel metal2 s 15741 1900 15769 2200 6 HI[399]
port 331 nsew signal tristate
rlabel metal2 s 15879 1900 15907 2200 6 HI[39]
port 332 nsew signal tristate
rlabel metal2 s 16017 1900 16045 2200 6 HI[3]
port 333 nsew signal tristate
rlabel metal2 s 16155 1900 16183 2200 6 HI[400]
port 334 nsew signal tristate
rlabel metal2 s 16293 1900 16321 2200 6 HI[401]
port 335 nsew signal tristate
rlabel metal2 s 16431 1900 16459 2200 6 HI[402]
port 336 nsew signal tristate
rlabel metal2 s 16569 1900 16597 2200 6 HI[403]
port 337 nsew signal tristate
rlabel metal2 s 16707 1900 16735 2200 6 HI[404]
port 338 nsew signal tristate
rlabel metal2 s 16845 1900 16873 2200 6 HI[405]
port 339 nsew signal tristate
rlabel metal2 s 16983 1900 17011 2200 6 HI[406]
port 340 nsew signal tristate
rlabel metal2 s 17121 1900 17149 2200 6 HI[407]
port 341 nsew signal tristate
rlabel metal2 s 17259 1900 17287 2200 6 HI[408]
port 342 nsew signal tristate
rlabel metal2 s 17397 1900 17425 2200 6 HI[409]
port 343 nsew signal tristate
rlabel metal2 s 17535 1900 17563 2200 6 HI[40]
port 344 nsew signal tristate
rlabel metal2 s 17673 1900 17701 2200 6 HI[410]
port 345 nsew signal tristate
rlabel metal2 s 17811 1900 17839 2200 6 HI[411]
port 346 nsew signal tristate
rlabel metal2 s 17949 1900 17977 2200 6 HI[412]
port 347 nsew signal tristate
rlabel metal2 s 18087 1900 18115 2200 6 HI[413]
port 348 nsew signal tristate
rlabel metal2 s 18225 1900 18253 2200 6 HI[414]
port 349 nsew signal tristate
rlabel metal2 s 18363 1900 18391 2200 6 HI[415]
port 350 nsew signal tristate
rlabel metal2 s 18501 1900 18529 2200 6 HI[416]
port 351 nsew signal tristate
rlabel metal2 s 18639 1900 18667 2200 6 HI[417]
port 352 nsew signal tristate
rlabel metal2 s 18777 1900 18805 2200 6 HI[418]
port 353 nsew signal tristate
rlabel metal2 s 18915 1900 18943 2200 6 HI[419]
port 354 nsew signal tristate
rlabel metal2 s 19053 1900 19081 2200 6 HI[41]
port 355 nsew signal tristate
rlabel metal2 s 19191 1900 19219 2200 6 HI[420]
port 356 nsew signal tristate
rlabel metal2 s 19329 1900 19357 2200 6 HI[421]
port 357 nsew signal tristate
rlabel metal2 s 19467 1900 19495 2200 6 HI[422]
port 358 nsew signal tristate
rlabel metal2 s 19605 1900 19633 2200 6 HI[423]
port 359 nsew signal tristate
rlabel metal2 s 19743 1900 19771 2200 6 HI[424]
port 360 nsew signal tristate
rlabel metal2 s 19881 1900 19909 2200 6 HI[425]
port 361 nsew signal tristate
rlabel metal2 s 20019 1900 20047 2200 6 HI[426]
port 362 nsew signal tristate
rlabel metal2 s 20157 1900 20185 2200 6 HI[427]
port 363 nsew signal tristate
rlabel metal2 s 20295 1900 20323 2200 6 HI[428]
port 364 nsew signal tristate
rlabel metal2 s 20433 1900 20461 2200 6 HI[429]
port 365 nsew signal tristate
rlabel metal2 s 20571 1900 20599 2200 6 HI[42]
port 366 nsew signal tristate
rlabel metal2 s 20709 1900 20737 2200 6 HI[430]
port 367 nsew signal tristate
rlabel metal2 s 20847 1900 20875 2200 6 HI[431]
port 368 nsew signal tristate
rlabel metal2 s 20985 1900 21013 2200 6 HI[432]
port 369 nsew signal tristate
rlabel metal2 s 21123 1900 21151 2200 6 HI[433]
port 370 nsew signal tristate
rlabel metal2 s 21261 1900 21289 2200 6 HI[434]
port 371 nsew signal tristate
rlabel metal2 s 21399 1900 21427 2200 6 HI[435]
port 372 nsew signal tristate
rlabel metal2 s 21537 1900 21565 2200 6 HI[436]
port 373 nsew signal tristate
rlabel metal2 s 21675 1900 21703 2200 6 HI[437]
port 374 nsew signal tristate
rlabel metal2 s 21813 1900 21841 2200 6 HI[438]
port 375 nsew signal tristate
rlabel metal2 s 21951 1900 21979 2200 6 HI[439]
port 376 nsew signal tristate
rlabel metal2 s 22089 1900 22117 2200 6 HI[43]
port 377 nsew signal tristate
rlabel metal2 s 22227 1900 22255 2200 6 HI[440]
port 378 nsew signal tristate
rlabel metal2 s 22365 1900 22393 2200 6 HI[441]
port 379 nsew signal tristate
rlabel metal2 s 22503 1900 22531 2200 6 HI[442]
port 380 nsew signal tristate
rlabel metal2 s 22641 1900 22669 2200 6 HI[443]
port 381 nsew signal tristate
rlabel metal2 s 22779 1900 22807 2200 6 HI[444]
port 382 nsew signal tristate
rlabel metal2 s 22917 1900 22945 2200 6 HI[445]
port 383 nsew signal tristate
rlabel metal2 s 23055 1900 23083 2200 6 HI[446]
port 384 nsew signal tristate
rlabel metal2 s 23193 1900 23221 2200 6 HI[447]
port 385 nsew signal tristate
rlabel metal2 s 23331 1900 23359 2200 6 HI[448]
port 386 nsew signal tristate
rlabel metal2 s 23469 1900 23497 2200 6 HI[449]
port 387 nsew signal tristate
rlabel metal2 s 23607 1900 23635 2200 6 HI[44]
port 388 nsew signal tristate
rlabel metal2 s 23745 1900 23773 2200 6 HI[450]
port 389 nsew signal tristate
rlabel metal2 s 23883 1900 23911 2200 6 HI[451]
port 390 nsew signal tristate
rlabel metal2 s 24021 1900 24049 2200 6 HI[452]
port 391 nsew signal tristate
rlabel metal2 s 24159 1900 24187 2200 6 HI[453]
port 392 nsew signal tristate
rlabel metal2 s 24297 1900 24325 2200 6 HI[454]
port 393 nsew signal tristate
rlabel metal2 s 24435 1900 24463 2200 6 HI[455]
port 394 nsew signal tristate
rlabel metal2 s 24573 1900 24601 2200 6 HI[456]
port 395 nsew signal tristate
rlabel metal2 s 24711 1900 24739 2200 6 HI[457]
port 396 nsew signal tristate
rlabel metal2 s 24849 1900 24877 2200 6 HI[458]
port 397 nsew signal tristate
rlabel metal2 s 24987 1900 25015 2200 6 HI[459]
port 398 nsew signal tristate
rlabel metal2 s 25125 1900 25153 2200 6 HI[45]
port 399 nsew signal tristate
rlabel metal2 s 25263 1900 25291 2200 6 HI[460]
port 400 nsew signal tristate
rlabel metal2 s 25401 1900 25429 2200 6 HI[461]
port 401 nsew signal tristate
rlabel metal2 s 25539 1900 25567 2200 6 HI[462]
port 402 nsew signal tristate
rlabel metal2 s 25677 1900 25705 2200 6 HI[46]
port 403 nsew signal tristate
rlabel metal2 s 25815 1900 25843 2200 6 HI[47]
port 404 nsew signal tristate
rlabel metal2 s 25953 1900 25981 2200 6 HI[48]
port 405 nsew signal tristate
rlabel metal2 s 26091 1900 26119 2200 6 HI[49]
port 406 nsew signal tristate
rlabel metal2 s 26229 1900 26257 2200 6 HI[4]
port 407 nsew signal tristate
rlabel metal2 s 26367 1900 26395 2200 6 HI[50]
port 408 nsew signal tristate
rlabel metal2 s 26505 1900 26533 2200 6 HI[51]
port 409 nsew signal tristate
rlabel metal2 s 26643 1900 26671 2200 6 HI[52]
port 410 nsew signal tristate
rlabel metal2 s 26781 1900 26809 2200 6 HI[53]
port 411 nsew signal tristate
rlabel metal2 s 26919 1900 26947 2200 6 HI[54]
port 412 nsew signal tristate
rlabel metal2 s 27057 1900 27085 2200 6 HI[55]
port 413 nsew signal tristate
rlabel metal2 s 27195 1900 27223 2200 6 HI[56]
port 414 nsew signal tristate
rlabel metal2 s 27333 1900 27361 2200 6 HI[57]
port 415 nsew signal tristate
rlabel metal2 s 27471 1900 27499 2200 6 HI[58]
port 416 nsew signal tristate
rlabel metal2 s 27609 1900 27637 2200 6 HI[59]
port 417 nsew signal tristate
rlabel metal2 s 27747 1900 27775 2200 6 HI[5]
port 418 nsew signal tristate
rlabel metal2 s 27885 1900 27913 2200 6 HI[60]
port 419 nsew signal tristate
rlabel metal2 s 28023 1900 28051 2200 6 HI[61]
port 420 nsew signal tristate
rlabel metal2 s 28161 1900 28189 2200 6 HI[62]
port 421 nsew signal tristate
rlabel metal2 s 28299 1900 28327 2200 6 HI[63]
port 422 nsew signal tristate
rlabel metal2 s 28437 1900 28465 2200 6 HI[64]
port 423 nsew signal tristate
rlabel metal2 s 28575 1900 28603 2200 6 HI[65]
port 424 nsew signal tristate
rlabel metal2 s 28713 1900 28741 2200 6 HI[66]
port 425 nsew signal tristate
rlabel metal2 s 28851 1900 28879 2200 6 HI[67]
port 426 nsew signal tristate
rlabel metal2 s 28989 1900 29017 2200 6 HI[68]
port 427 nsew signal tristate
rlabel metal2 s 29127 1900 29155 2200 6 HI[69]
port 428 nsew signal tristate
rlabel metal2 s 29265 1900 29293 2200 6 HI[6]
port 429 nsew signal tristate
rlabel metal2 s 29403 1900 29431 2200 6 HI[70]
port 430 nsew signal tristate
rlabel metal2 s 29541 1900 29569 2200 6 HI[71]
port 431 nsew signal tristate
rlabel metal2 s 29679 1900 29707 2200 6 HI[72]
port 432 nsew signal tristate
rlabel metal2 s 29817 1900 29845 2200 6 HI[73]
port 433 nsew signal tristate
rlabel metal2 s 29955 1900 29983 2200 6 HI[74]
port 434 nsew signal tristate
rlabel metal2 s 30093 1900 30121 2200 6 HI[75]
port 435 nsew signal tristate
rlabel metal2 s 30231 1900 30259 2200 6 HI[76]
port 436 nsew signal tristate
rlabel metal2 s 30369 1900 30397 2200 6 HI[77]
port 437 nsew signal tristate
rlabel metal2 s 30507 1900 30535 2200 6 HI[78]
port 438 nsew signal tristate
rlabel metal2 s 30645 1900 30673 2200 6 HI[79]
port 439 nsew signal tristate
rlabel metal2 s 30783 1900 30811 2200 6 HI[7]
port 440 nsew signal tristate
rlabel metal2 s 30921 1900 30949 2200 6 HI[80]
port 441 nsew signal tristate
rlabel metal2 s 31059 1900 31087 2200 6 HI[81]
port 442 nsew signal tristate
rlabel metal2 s 31197 1900 31225 2200 6 HI[82]
port 443 nsew signal tristate
rlabel metal2 s 31335 1900 31363 2200 6 HI[83]
port 444 nsew signal tristate
rlabel metal2 s 31473 1900 31501 2200 6 HI[84]
port 445 nsew signal tristate
rlabel metal2 s 31611 1900 31639 2200 6 HI[85]
port 446 nsew signal tristate
rlabel metal2 s 31749 1900 31777 2200 6 HI[86]
port 447 nsew signal tristate
rlabel metal2 s 31887 1900 31915 2200 6 HI[87]
port 448 nsew signal tristate
rlabel metal2 s 32025 1900 32053 2200 6 HI[88]
port 449 nsew signal tristate
rlabel metal2 s 32163 1900 32191 2200 6 HI[89]
port 450 nsew signal tristate
rlabel metal2 s 32301 1900 32329 2200 6 HI[8]
port 451 nsew signal tristate
rlabel metal2 s 32439 1900 32467 2200 6 HI[90]
port 452 nsew signal tristate
rlabel metal2 s 32577 1900 32605 2200 6 HI[91]
port 453 nsew signal tristate
rlabel metal2 s 32715 1900 32743 2200 6 HI[92]
port 454 nsew signal tristate
rlabel metal2 s 32853 1900 32881 2200 6 HI[93]
port 455 nsew signal tristate
rlabel metal2 s 32991 1900 33019 2200 6 HI[94]
port 456 nsew signal tristate
rlabel metal2 s 33129 1900 33157 2200 6 HI[95]
port 457 nsew signal tristate
rlabel metal2 s 33267 1900 33295 2200 6 HI[96]
port 458 nsew signal tristate
rlabel metal2 s 33405 1900 33433 2200 6 HI[97]
port 459 nsew signal tristate
rlabel metal2 s 33543 1900 33571 2200 6 HI[98]
port 460 nsew signal tristate
rlabel metal2 s 33681 1900 33709 2200 6 HI[99]
port 461 nsew signal tristate
rlabel metal2 s 33819 1900 33847 2200 6 HI[9]
port 462 nsew signal tristate
rlabel metal3 s 644 595 34408 645 6 vccd1
port 463 nsew power input
rlabel metal2 s 3619 520 3669 1656 6 vccd1
port 463 nsew power input
rlabel metal2 s 9619 520 9669 1656 6 vccd1
port 463 nsew power input
rlabel metal2 s 15619 520 15669 1656 6 vccd1
port 463 nsew power input
rlabel metal2 s 21619 520 21669 1656 6 vccd1
port 463 nsew power input
rlabel metal2 s 27619 520 27669 1656 6 vccd1
port 463 nsew power input
rlabel metal2 s 33619 520 33669 1656 6 vccd1
port 463 nsew power input
rlabel metal3 s 644 1135 34408 1185 6 vssd1
port 464 nsew ground input
rlabel metal2 s 6619 520 6669 1656 6 vssd1
port 464 nsew ground input
rlabel metal2 s 12619 520 12669 1656 6 vssd1
port 464 nsew ground input
rlabel metal2 s 18619 520 18669 1656 6 vssd1
port 464 nsew ground input
rlabel metal2 s 24619 520 24669 1656 6 vssd1
port 464 nsew ground input
rlabel metal2 s 30619 520 30669 1656 6 vssd1
port 464 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 35000 2200
<< end >>
