* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_2 abstract view
.subckt sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for gpio_logic_high abstract view
.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
X_131_ _131_/CLK hold1/A resetn vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__dfrtp_2
X_062_ _105_/Q user_gpio_oeb vssd vssd vccd vccd _062_/X sky130_fd_sc_hd__and2b_2
XANTENNA__132__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_114_ _101__10/Y hold1/X _085_/X _086_/Y vssd vssd vccd vccd pad_gpio_dm[2] _114_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_130_ _133_/A _130_/D resetn vssd vssd vccd vccd hold1/A sky130_fd_sc_hd__dfrtp_2
X_061_ pad_gpio_inenb _111_/Q vssd vssd vccd vccd _061_/Y sky130_fd_sc_hd__nand2b_2
X_113_ _100__9/Y _130_/D _083_/X _084_/Y vssd vssd vccd vccd pad_gpio_dm[1] _113_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
Xclkbuf_1_0__f_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _100__9/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__135__A pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_104__13 _100__9/A vssd vssd vccd vccd _104__13/Y sky130_fd_sc_hd__inv_2
X_094__3 _134_/A vssd vssd vccd vccd _094__3/Y sky130_fd_sc_hd__inv_2
XFILLER_18_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xhold10 _124_/Q vssd vssd vccd vccd _125_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__122__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_112_ _099__8/Y hold8/X _081_/X _082_/Y vssd vssd vccd vccd pad_gpio_dm[0] _065_/A1
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__065__A0 mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__061__A_N pad_gpio_inenb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__084__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_111_ _098__7/Y hold5/X _079_/X _080_/Y vssd vssd vccd vccd _111_/Q _111_/Q_N sky130_fd_sc_hd__dfbbn_2
XANTENNA__067__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold11 _125_/Q vssd vssd vccd vccd _126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__075__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_79 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__131__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__072__B gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__074__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_110_ _097__6/Y hold9/X _077_/X _078_/Y vssd vssd vccd vccd pad_gpio_ib_mode_sel
+ _110_/Q_N sky130_fd_sc_hd__dfbbn_2
Xhold12 _123_/Q vssd vssd vccd vccd _124_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__067__B gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__083__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__080__B gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__064__C mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__075__B gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__091__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold13 _129_/Q vssd vssd vccd vccd _130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_097__6 _100__9/A vssd vssd vccd vccd _097__6/Y sky130_fd_sc_hd__inv_2
XANTENNA__083__B gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__078__B gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__064__A_N pad_gpio_dm[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__089__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__125__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__091__B gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__086__B gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__089__B gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
XANTENNA__119__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_079_ resetn gpio_defaults[1] vssd vssd vccd vccd _079_/X sky130_fd_sc_hd__or2_2
XANTENNA__128__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__090__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_078_ resetn gpio_defaults[4] vssd vssd vccd vccd _078_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_7_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__080__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_100__9 _100__9/A vssd vssd vccd vccd _100__9/Y sky130_fd_sc_hd__inv_2
X_077_ resetn gpio_defaults[4] vssd vssd vccd vccd _077_/X sky130_fd_sc_hd__or2_2
X_129_ _133_/A hold8/X resetn vssd vssd vccd vccd _129_/Q sky130_fd_sc_hd__dfrtp_2
X_103__12 _100__9/A vssd vssd vccd vccd _103__12/Y sky130_fd_sc_hd__inv_2
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_076_ resetn gpio_defaults[3] vssd vssd vccd vccd _076_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_10_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__070__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_128_ _133_/A hold2/X resetn vssd vssd vccd vccd hold8/A sky130_fd_sc_hd__dfrtp_2
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__121__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_092_ resetn gpio_defaults[7] vssd vssd vccd vccd _092_/Y sky130_fd_sc_hd__nand2b_2
Xgpio_in_buf _058_/Y gpio_in_buf/TE vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_075_ resetn gpio_defaults[3] vssd vssd vccd vccd _075_/X sky130_fd_sc_hd__or2_2
X_058_ pad_gpio_in vssd vssd vccd vccd _058_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_serial_load_A serial_load vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_127_ _133_/A hold7/X resetn vssd vssd vccd vccd hold2/A sky130_fd_sc_hd__dfrtp_2
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_074_ resetn gpio_defaults[9] vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__nand2b_2
X_091_ resetn gpio_defaults[7] vssd vssd vccd vccd _091_/X sky130_fd_sc_hd__or2_2
X_126_ _126_/CLK _126_/D resetn vssd vssd vccd vccd hold7/A sky130_fd_sc_hd__dfrtp_2
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_095__4 _134_/A vssd vssd vccd vccd _095__4/Y sky130_fd_sc_hd__inv_2
XFILLER_13_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_109_ _096__5/Y hold4/X _075_/X _076_/Y vssd vssd vccd vccd pad_gpio_inenb _109_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__130__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_60 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ resetn gpio_defaults[6] vssd vssd vccd vccd _090_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__073__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__062__B user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_073_ resetn gpio_defaults[9] vssd vssd vccd vccd _073_/X sky130_fd_sc_hd__or2_2
XFILLER_2_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_125_ _126_/CLK _125_/D resetn vssd vssd vccd vccd _125_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__070__B gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_108_ _095__4/Y hold2/X _073_/X _074_/Y vssd vssd vccd vccd pad_gpio_vtrip_sel _108_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__081__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_61 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_072_ resetn gpio_defaults[8] vssd vssd vccd vccd _072_/Y sky130_fd_sc_hd__nand2b_2
XTAP_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__086__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__068__B gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__073__B gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_124_ _126_/CLK _124_/D resetn vssd vssd vccd vccd _124_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__079__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_107_ _094__3/Y hold7/X _071_/X _072_/Y vssd vssd vccd vccd pad_gpio_slow_sel _107_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__124__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_060__14 _133_/A vssd vssd vccd vccd _131_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__076__B gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__081__B gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_62 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_071_ resetn gpio_defaults[8] vssd vssd vccd vccd _071_/X sky130_fd_sc_hd__or2_2
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__087__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_40 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_106_ _093__2/Y hold3/X _069_/X _070_/Y vssd vssd vccd vccd pad_gpio_holdover _106_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
X_123_ _126_/CLK hold9/X resetn vssd vssd vccd vccd _123_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__084__B gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__079__B gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__076__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_070_ resetn gpio_defaults[2] vssd vssd vccd vccd _070_/Y sky130_fd_sc_hd__nand2b_2
XTAP_63 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__118__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__092__B gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__087__B gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_41 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_098__7 _134_/A vssd vssd vccd vccd _098__7/Y sky130_fd_sc_hd__inv_2
X_122_ _126_/CLK hold4/X resetn vssd vssd vccd vccd hold9/A sky130_fd_sc_hd__dfrtp_2
XFILLER_2_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_105_ _059__1/Y hold6/X _067_/X _068_/Y vssd vssd vccd vccd _105_/Q _105_/Q_N sky130_fd_sc_hd__dfbbn_2
XTAP_64 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ _126_/CLK hold3/X resetn vssd vssd vccd vccd hold4/A sky130_fd_sc_hd__dfrtp_2
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_65 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_54 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ _126_/CLK hold5/X resetn vssd vssd vccd vccd hold3/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__127__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd vssd vccd vccd hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_55 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_102__11 _100__9/A vssd vssd vccd vccd _102__11/Y sky130_fd_sc_hd__inv_2
Xhold2 hold2/A vssd vssd vccd vccd hold2/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_serial_load serial_load vssd vssd vccd vccd clkbuf_0_serial_load/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_56 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
XFILLER_2_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold3 hold3/A vssd vssd vccd vccd hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_57 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__120__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd vssd vccd vccd hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__092__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_58 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_093__2 _134_/A vssd vssd vccd vccd _093__2/Y sky130_fd_sc_hd__inv_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xhold5 hold5/A vssd vssd vccd vccd hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__082__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_59 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd vssd vccd vccd hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_089_ resetn gpio_defaults[6] vssd vssd vccd vccd _089_/X sky130_fd_sc_hd__or2_2
XTAP_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__072__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__063__A2 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__118__D serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_088_ resetn gpio_defaults[5] vssd vssd vccd vccd _088_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__058__A pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd vssd vccd vccd hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__071__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_39 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__066__A0 user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__123__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _134_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__069__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_087_ resetn gpio_defaults[5] vssd vssd vccd vccd _087_/X sky130_fd_sc_hd__or2_2
Xhold8 hold8/A vssd vssd vccd vccd hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_096__5 _134_/A vssd vssd vccd vccd _096__5/Y sky130_fd_sc_hd__inv_2
XANTENNA__071__B gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__077__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_086_ resetn gpio_defaults[12] vssd vssd vccd vccd _086_/Y sky130_fd_sc_hd__nand2b_2
XANTENNA__074__B gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_11_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__085__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_069_ resetn gpio_defaults[2] vssd vssd vccd vccd _069_/X sky130_fd_sc_hd__or2_2
XANTENNA__069__B gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd vssd vccd vccd hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__082__B gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__077__B gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__085__B gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_085_ resetn gpio_defaults[12] vssd vssd vccd vccd _085_/X sky130_fd_sc_hd__or2_2
XANTENNA__090__B gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_068_ resetn gpio_defaults[0] vssd vssd vccd vccd _068_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_50 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__088__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__088__B gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_067_ resetn gpio_defaults[0] vssd vssd vccd vccd _067_/X sky130_fd_sc_hd__or2_2
XFILLER_8_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_084_ resetn gpio_defaults[11] vssd vssd vccd vccd _084_/Y sky130_fd_sc_hd__nand2b_2
X_119_ _126_/CLK hold6/X resetn vssd vssd vccd vccd hold5/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__126__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_101__10 _134_/A vssd vssd vccd vccd _101__10/Y sky130_fd_sc_hd__inv_2
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__078__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_083_ resetn gpio_defaults[11] vssd vssd vccd vccd _083_/X sky130_fd_sc_hd__or2_2
X_099__8 _100__9/A vssd vssd vccd vccd _099__8/Y sky130_fd_sc_hd__inv_2
XFILLER_18_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_118_ _133_/A serial_data_in resetn vssd vssd vccd vccd hold6/A sky130_fd_sc_hd__dfrtp_2
X_066_ user_gpio_out _065_/X _105_/Q vssd vssd vccd vccd pad_gpio_out sky130_fd_sc_hd__mux2_1
X_135_ pad_gpio_in _061_/Y vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_2
XFILLER_0_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_134_ _134_/A vssd vssd vccd vccd serial_load_out sky130_fd_sc_hd__buf_2
X_059__1 _134_/A vssd vssd vccd vccd _059__1/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_082_ resetn gpio_defaults[10] vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__nand2b_2
X_065_ mgmt_gpio_out _065_/A1 _065_/S vssd vssd vccd vccd _065_/X sky130_fd_sc_hd__mux2_1
XANTENNA__068__A_N resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_117_ _104__13/Y _126_/D _091_/X _092_/Y vssd vssd vccd vccd pad_gpio_ana_pol _117_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_081_ resetn gpio_defaults[10] vssd vssd vccd vccd _081_/X sky130_fd_sc_hd__or2_2
X_133_ _133_/A vssd vssd vccd vccd serial_clock_out sky130_fd_sc_hd__buf_2
X_064_ pad_gpio_dm[2] pad_gpio_dm[1] mgmt_gpio_oeb vssd vssd vccd vccd _065_/S sky130_fd_sc_hd__and3b_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_116_ _103__12/Y _125_/D _089_/X _090_/Y vssd vssd vccd vccd pad_gpio_ana_sel _116_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA_clkbuf_0_serial_clock_A serial_clock vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_080_ resetn gpio_defaults[1] vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__nand2b_2
X_132_ resetn vssd vssd vccd vccd resetn_out sky130_fd_sc_hd__buf_2
X_063_ _111_/Q mgmt_gpio_oeb _105_/Q _062_/X vssd vssd vccd vccd pad_gpio_outenb sky130_fd_sc_hd__a31o_2
XANTENNA__129__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_115_ _102__11/Y _124_/D _087_/X _088_/Y vssd vssd vccd vccd pad_gpio_ana_en _115_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
.ends

