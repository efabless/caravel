VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_defaults_block
  CLASS BLOCK ;
  FOREIGN gpio_defaults_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.000 BY 28.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 13.400 5.200 14.800 22.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.060 16.340 16.340 17.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 4.000 5.200 5.400 22.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.060 8.940 16.340 10.340 ;
    END
  END VPWR
  PIN gpio_defaults[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 3.770 25.000 4.050 31.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 21.120 3.000 21.720 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 3.770 -3.000 4.050 3.000 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 5.610 -3.000 5.890 3.000 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 5.610 25.000 5.890 31.000 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 4.800 3.000 5.400 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 6.160 3.000 6.760 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 7.520 3.000 8.120 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 11.600 3.000 12.200 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 12.960 3.000 13.560 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 14.320 3.000 14.920 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 18.400 3.000 19.000 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT -3.000 19.760 3.000 20.360 ;
    END
  END gpio_defaults[9]
  OBS
      LAYER li1 ;
        RECT 0.000 0.000 17.000 28.000 ;
      LAYER met1 ;
        RECT 0.000 0.000 17.000 28.000 ;
      LAYER met2 ;
        RECT 0.000 0.000 17.000 28.000 ;
      LAYER met3 ;
        RECT 0.000 0.000 17.000 28.000 ;
  END
END gpio_defaults_block
END LIBRARY

