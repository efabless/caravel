module user_id_textblock ();
endmodule
