VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 75.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.040 5.200 42.640 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 5.200 82.640 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.050 94.540 42.650 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 5.200 62.640 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 21.050 94.540 22.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 61.050 94.540 62.650 ;
    END
  END VPWR
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 71.000 27.970 75.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 71.000 35.330 75.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 71.000 42.690 75.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 71.000 50.050 75.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 71.000 57.410 75.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 71.000 64.770 75.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 71.000 72.130 75.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 71.000 79.490 75.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 71.000 86.850 75.000 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 71.000 94.210 75.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 67.360 100.000 67.960 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.120 100.000 55.720 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 42.880 100.000 43.480 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 18.400 100.000 19.000 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.160 100.000 6.760 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 71.000 5.890 75.000 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 71.000 13.250 75.000 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 71.000 20.610 75.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END resetb
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 94.300 68.085 ;
      LAYER met1 ;
        RECT 5.520 4.460 94.300 68.640 ;
      LAYER met2 ;
        RECT 6.170 70.720 12.690 71.810 ;
        RECT 13.530 70.720 20.050 71.810 ;
        RECT 20.890 70.720 27.410 71.810 ;
        RECT 28.250 70.720 34.770 71.810 ;
        RECT 35.610 70.720 42.130 71.810 ;
        RECT 42.970 70.720 49.490 71.810 ;
        RECT 50.330 70.720 56.850 71.810 ;
        RECT 57.690 70.720 64.210 71.810 ;
        RECT 65.050 70.720 71.570 71.810 ;
        RECT 72.410 70.720 78.930 71.810 ;
        RECT 79.770 70.720 86.290 71.810 ;
        RECT 87.130 70.720 93.650 71.810 ;
        RECT 5.890 4.280 94.210 70.720 ;
        RECT 5.890 3.670 24.650 4.280 ;
        RECT 25.490 3.670 74.330 4.280 ;
        RECT 75.170 3.670 94.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 66.960 95.600 68.165 ;
        RECT 4.000 64.280 96.000 66.960 ;
        RECT 4.400 62.880 96.000 64.280 ;
        RECT 4.000 60.200 96.000 62.880 ;
        RECT 4.400 58.800 96.000 60.200 ;
        RECT 4.000 56.120 96.000 58.800 ;
        RECT 4.400 54.720 95.600 56.120 ;
        RECT 4.000 52.040 96.000 54.720 ;
        RECT 4.400 50.640 96.000 52.040 ;
        RECT 4.000 47.960 96.000 50.640 ;
        RECT 4.400 46.560 96.000 47.960 ;
        RECT 4.000 43.880 96.000 46.560 ;
        RECT 4.400 42.480 95.600 43.880 ;
        RECT 4.000 39.800 96.000 42.480 ;
        RECT 4.400 38.400 96.000 39.800 ;
        RECT 4.000 35.720 96.000 38.400 ;
        RECT 4.400 34.320 96.000 35.720 ;
        RECT 4.000 31.640 96.000 34.320 ;
        RECT 4.400 30.240 95.600 31.640 ;
        RECT 4.000 27.560 96.000 30.240 ;
        RECT 4.400 26.160 96.000 27.560 ;
        RECT 4.000 23.480 96.000 26.160 ;
        RECT 4.400 22.080 96.000 23.480 ;
        RECT 4.000 19.400 96.000 22.080 ;
        RECT 4.400 18.000 95.600 19.400 ;
        RECT 4.000 15.320 96.000 18.000 ;
        RECT 4.400 13.920 96.000 15.320 ;
        RECT 4.000 11.240 96.000 13.920 ;
        RECT 4.400 9.840 96.000 11.240 ;
        RECT 4.000 7.160 96.000 9.840 ;
        RECT 4.400 5.760 95.600 7.160 ;
        RECT 4.000 5.275 96.000 5.760 ;
  END
END digital_pll
END LIBRARY

