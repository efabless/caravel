magic
tech sky130A
magscale 1 2
timestamp 1665595735
<< nwell >>
rect 330 4613 7582 4934
rect 330 3525 7582 4091
rect 330 2437 7582 3003
rect 330 1349 7582 1915
<< obsli1 >>
rect 368 1071 7544 4913
<< obsm1 >>
rect 368 1040 7699 4944
<< metal2 >>
rect 478 5200 534 6000
rect 846 5200 902 6000
rect 1214 5200 1270 6000
rect 1582 5200 1638 6000
rect 1950 5200 2006 6000
rect 2318 5200 2374 6000
rect 2686 5200 2742 6000
rect 3054 5200 3110 6000
rect 3422 5200 3478 6000
rect 3790 5200 3846 6000
rect 4158 5200 4214 6000
rect 4526 5200 4582 6000
rect 4894 5200 4950 6000
rect 5262 5200 5318 6000
rect 5630 5200 5686 6000
rect 5998 5200 6054 6000
rect 6366 5200 6422 6000
rect 6734 5200 6790 6000
rect 7102 5200 7158 6000
rect 7470 5200 7526 6000
rect 478 0 534 800
rect 846 0 902 800
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
<< obsm2 >>
rect 590 5144 790 5250
rect 958 5144 1158 5250
rect 1326 5144 1526 5250
rect 1694 5144 1894 5250
rect 2062 5144 2262 5250
rect 2430 5144 2630 5250
rect 2798 5144 2998 5250
rect 3166 5144 3366 5250
rect 3534 5144 3734 5250
rect 3902 5144 4102 5250
rect 4270 5144 4470 5250
rect 4638 5144 4838 5250
rect 5006 5144 5206 5250
rect 5374 5144 5574 5250
rect 5742 5144 5942 5250
rect 6110 5144 6310 5250
rect 6478 5144 6678 5250
rect 6846 5144 7046 5250
rect 7214 5144 7414 5250
rect 7582 5144 7693 5250
rect 480 856 7693 5144
rect 590 800 790 856
rect 958 800 1158 856
rect 1326 800 1526 856
rect 1694 800 1894 856
rect 2062 800 2262 856
rect 2430 800 2630 856
rect 2798 800 2998 856
rect 3166 800 3366 856
rect 3534 800 3734 856
rect 3902 800 4102 856
rect 4270 800 4470 856
rect 4638 800 4838 856
rect 5006 800 5206 856
rect 5374 800 5574 856
rect 5742 800 5942 856
rect 6110 800 6310 856
rect 6478 800 6678 856
rect 6846 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7693 856
<< obsm3 >>
rect 1106 1055 7697 4929
<< metal4 >>
rect 1104 1040 1424 4944
rect 2000 1040 2320 4944
rect 2897 1040 3217 4944
rect 3793 1040 4113 4944
rect 4690 1040 5010 4944
rect 5586 1040 5906 4944
rect 6483 1040 6803 4944
rect 7379 1040 7699 4944
<< labels >>
rlabel metal4 s 2000 1040 2320 4944 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3793 1040 4113 4944 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5586 1040 5906 4944 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7379 1040 7699 4944 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1104 1040 1424 4944 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 2897 1040 3217 4944 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4690 1040 5010 4944 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6483 1040 6803 4944 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 478 0 534 800 6 in[0]
port 3 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 in[10]
port 4 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 in[11]
port 5 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 in[12]
port 6 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 in[13]
port 7 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 in[14]
port 8 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 in[15]
port 9 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 in[16]
port 10 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 in[17]
port 11 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 in[18]
port 12 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 in[19]
port 13 nsew signal input
rlabel metal2 s 846 0 902 800 6 in[1]
port 14 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 in[2]
port 15 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 in[3]
port 16 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 in[4]
port 17 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 in[5]
port 18 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 in[6]
port 19 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 in[7]
port 20 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 in[8]
port 21 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 in[9]
port 22 nsew signal input
rlabel metal2 s 478 5200 534 6000 6 out[0]
port 23 nsew signal output
rlabel metal2 s 4158 5200 4214 6000 6 out[10]
port 24 nsew signal output
rlabel metal2 s 4526 5200 4582 6000 6 out[11]
port 25 nsew signal output
rlabel metal2 s 4894 5200 4950 6000 6 out[12]
port 26 nsew signal output
rlabel metal2 s 5262 5200 5318 6000 6 out[13]
port 27 nsew signal output
rlabel metal2 s 5630 5200 5686 6000 6 out[14]
port 28 nsew signal output
rlabel metal2 s 5998 5200 6054 6000 6 out[15]
port 29 nsew signal output
rlabel metal2 s 6366 5200 6422 6000 6 out[16]
port 30 nsew signal output
rlabel metal2 s 6734 5200 6790 6000 6 out[17]
port 31 nsew signal output
rlabel metal2 s 7102 5200 7158 6000 6 out[18]
port 32 nsew signal output
rlabel metal2 s 7470 5200 7526 6000 6 out[19]
port 33 nsew signal output
rlabel metal2 s 846 5200 902 6000 6 out[1]
port 34 nsew signal output
rlabel metal2 s 1214 5200 1270 6000 6 out[2]
port 35 nsew signal output
rlabel metal2 s 1582 5200 1638 6000 6 out[3]
port 36 nsew signal output
rlabel metal2 s 1950 5200 2006 6000 6 out[4]
port 37 nsew signal output
rlabel metal2 s 2318 5200 2374 6000 6 out[5]
port 38 nsew signal output
rlabel metal2 s 2686 5200 2742 6000 6 out[6]
port 39 nsew signal output
rlabel metal2 s 3054 5200 3110 6000 6 out[7]
port 40 nsew signal output
rlabel metal2 s 3422 5200 3478 6000 6 out[8]
port 41 nsew signal output
rlabel metal2 s 3790 5200 3846 6000 6 out[9]
port 42 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8000 6000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 107194
string GDS_FILE /home/hosni/My_forks/caravel/openlane/buff8x20/runs/RUN_2022.10.12_17.28.33/results/signoff/buff8x20.magic.gds
string GDS_START 29274
<< end >>

