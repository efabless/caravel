magic
tech sky130A
magscale 1 2
timestamp 1675162489
<< viali >>
rect 1593 4233 1627 4267
rect 949 3961 983 3995
rect 2329 3689 2363 3723
rect 1501 3553 1535 3587
rect 1317 3009 1351 3043
rect 1961 2873 1995 2907
rect 1501 2601 1535 2635
rect 2329 2397 2363 2431
rect 2237 1785 2271 1819
rect 949 1717 983 1751
rect 1593 1717 1627 1751
rect 1593 1513 1627 1547
rect 949 1377 983 1411
<< metal1 >>
rect 460 4378 3220 4400
rect 460 4326 2698 4378
rect 2750 4326 2762 4378
rect 2814 4326 2826 4378
rect 2878 4326 2890 4378
rect 2942 4326 3220 4378
rect 460 4304 3220 4326
rect 1302 4224 1308 4276
rect 1360 4264 1366 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1360 4236 1593 4264
rect 1360 4224 1366 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 937 3995 995 4001
rect 937 3961 949 3995
rect 983 3992 995 3995
rect 1118 3992 1124 4004
rect 983 3964 1124 3992
rect 983 3961 995 3964
rect 937 3955 995 3961
rect 1118 3952 1124 3964
rect 1176 3952 1182 4004
rect 460 3834 3220 3856
rect 460 3782 818 3834
rect 870 3782 882 3834
rect 934 3782 946 3834
rect 998 3782 1010 3834
rect 1062 3782 3220 3834
rect 460 3760 3220 3782
rect 1302 3680 1308 3732
rect 1360 3720 1366 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1360 3692 2329 3720
rect 1360 3680 1366 3692
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 2317 3683 2375 3689
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1489 3587 1547 3593
rect 1489 3584 1501 3587
rect 1452 3556 1501 3584
rect 1452 3544 1458 3556
rect 1489 3553 1501 3556
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 460 3290 3220 3312
rect 460 3238 2698 3290
rect 2750 3238 2762 3290
rect 2814 3238 2826 3290
rect 2878 3238 2890 3290
rect 2942 3238 3220 3290
rect 460 3216 3220 3238
rect 658 3000 664 3052
rect 716 3040 722 3052
rect 1305 3043 1363 3049
rect 1305 3040 1317 3043
rect 716 3012 1317 3040
rect 716 3000 722 3012
rect 1305 3009 1317 3012
rect 1351 3009 1363 3043
rect 1305 3003 1363 3009
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 1949 2907 2007 2913
rect 1949 2904 1961 2907
rect 1176 2876 1961 2904
rect 1176 2864 1182 2876
rect 1949 2873 1961 2876
rect 1995 2873 2007 2907
rect 1949 2867 2007 2873
rect 460 2746 3220 2768
rect 460 2694 818 2746
rect 870 2694 882 2746
rect 934 2694 946 2746
rect 998 2694 1010 2746
rect 1062 2694 3220 2746
rect 460 2672 3220 2694
rect 1302 2592 1308 2644
rect 1360 2632 1366 2644
rect 1489 2635 1547 2641
rect 1489 2632 1501 2635
rect 1360 2604 1501 2632
rect 1360 2592 1366 2604
rect 1489 2601 1501 2604
rect 1535 2601 1547 2635
rect 1489 2595 1547 2601
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 1268 2400 2329 2428
rect 1268 2388 1274 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 460 2202 3220 2224
rect 460 2150 2698 2202
rect 2750 2150 2762 2202
rect 2814 2150 2826 2202
rect 2878 2150 2890 2202
rect 2942 2150 3220 2202
rect 460 2128 3220 2150
rect 566 1776 572 1828
rect 624 1816 630 1828
rect 2225 1819 2283 1825
rect 2225 1816 2237 1819
rect 624 1788 2237 1816
rect 624 1776 630 1788
rect 2225 1785 2237 1788
rect 2271 1785 2283 1819
rect 2225 1779 2283 1785
rect 658 1708 664 1760
rect 716 1748 722 1760
rect 937 1751 995 1757
rect 937 1748 949 1751
rect 716 1720 949 1748
rect 716 1708 722 1720
rect 937 1717 949 1720
rect 983 1717 995 1751
rect 937 1711 995 1717
rect 1210 1708 1216 1760
rect 1268 1748 1274 1760
rect 1581 1751 1639 1757
rect 1581 1748 1593 1751
rect 1268 1720 1593 1748
rect 1268 1708 1274 1720
rect 1581 1717 1593 1720
rect 1627 1717 1639 1751
rect 1581 1711 1639 1717
rect 460 1658 3220 1680
rect 460 1606 818 1658
rect 870 1606 882 1658
rect 934 1606 946 1658
rect 998 1606 1010 1658
rect 1062 1606 3220 1658
rect 460 1584 3220 1606
rect 1302 1504 1308 1556
rect 1360 1544 1366 1556
rect 1581 1547 1639 1553
rect 1581 1544 1593 1547
rect 1360 1516 1593 1544
rect 1360 1504 1366 1516
rect 1581 1513 1593 1516
rect 1627 1513 1639 1547
rect 1581 1507 1639 1513
rect 937 1411 995 1417
rect 937 1377 949 1411
rect 983 1408 995 1411
rect 1118 1408 1124 1420
rect 983 1380 1124 1408
rect 983 1377 995 1380
rect 937 1371 995 1377
rect 1118 1368 1124 1380
rect 1176 1368 1182 1420
rect 460 1114 3220 1136
rect 460 1062 2698 1114
rect 2750 1062 2762 1114
rect 2814 1062 2826 1114
rect 2878 1062 2890 1114
rect 2942 1062 3220 1114
rect 460 1040 3220 1062
<< via1 >>
rect 2698 4326 2750 4378
rect 2762 4326 2814 4378
rect 2826 4326 2878 4378
rect 2890 4326 2942 4378
rect 1308 4224 1360 4276
rect 1124 3952 1176 4004
rect 818 3782 870 3834
rect 882 3782 934 3834
rect 946 3782 998 3834
rect 1010 3782 1062 3834
rect 1308 3680 1360 3732
rect 1400 3544 1452 3596
rect 2698 3238 2750 3290
rect 2762 3238 2814 3290
rect 2826 3238 2878 3290
rect 2890 3238 2942 3290
rect 664 3000 716 3052
rect 1124 2864 1176 2916
rect 818 2694 870 2746
rect 882 2694 934 2746
rect 946 2694 998 2746
rect 1010 2694 1062 2746
rect 1308 2592 1360 2644
rect 1216 2388 1268 2440
rect 2698 2150 2750 2202
rect 2762 2150 2814 2202
rect 2826 2150 2878 2202
rect 2890 2150 2942 2202
rect 572 1776 624 1828
rect 664 1708 716 1760
rect 1216 1708 1268 1760
rect 818 1606 870 1658
rect 882 1606 934 1658
rect 946 1606 998 1658
rect 1010 1606 1062 1658
rect 1308 1504 1360 1556
rect 1124 1368 1176 1420
rect 2698 1062 2750 1114
rect 2762 1062 2814 1114
rect 2826 1062 2878 1114
rect 2890 1062 2942 1114
<< metal2 >>
rect 754 5114 810 6200
rect 676 5086 810 5114
rect 676 3058 704 5086
rect 754 5000 810 5086
rect 1122 5114 1178 6200
rect 1122 5086 1256 5114
rect 1122 5000 1178 5086
rect 800 3834 1080 4400
rect 1122 4040 1178 4049
rect 1122 3975 1124 3984
rect 1176 3975 1178 3984
rect 1124 3946 1176 3952
rect 800 3782 818 3834
rect 870 3782 882 3834
rect 934 3782 946 3834
rect 998 3782 1010 3834
rect 1062 3782 1080 3834
rect 664 3052 716 3058
rect 664 2994 716 3000
rect 800 2746 1080 3782
rect 1228 3618 1256 5086
rect 2680 4378 2960 4400
rect 2680 4326 2698 4378
rect 2750 4326 2762 4378
rect 2814 4326 2826 4378
rect 2878 4326 2890 4378
rect 2942 4326 2960 4378
rect 1306 4312 1362 4321
rect 1306 4247 1308 4256
rect 1360 4247 1362 4256
rect 1308 4218 1360 4224
rect 1306 3768 1362 3777
rect 1306 3703 1308 3712
rect 1360 3703 1362 3712
rect 1308 3674 1360 3680
rect 1228 3602 1440 3618
rect 1228 3596 1452 3602
rect 1228 3590 1400 3596
rect 1400 3538 1452 3544
rect 2680 3516 2960 4326
rect 2680 3460 2712 3516
rect 2768 3460 2792 3516
rect 2848 3460 2872 3516
rect 2928 3460 2960 3516
rect 2680 3436 2960 3460
rect 2680 3380 2712 3436
rect 2768 3380 2792 3436
rect 2848 3380 2872 3436
rect 2928 3380 2960 3436
rect 2680 3356 2960 3380
rect 2680 3300 2712 3356
rect 2768 3300 2792 3356
rect 2848 3300 2872 3356
rect 2928 3300 2960 3356
rect 2680 3290 2960 3300
rect 2680 3238 2698 3290
rect 2750 3238 2762 3290
rect 2814 3238 2826 3290
rect 2878 3238 2890 3290
rect 2942 3238 2960 3290
rect 1122 2952 1178 2961
rect 1122 2887 1124 2896
rect 1176 2887 1178 2896
rect 1124 2858 1176 2864
rect 800 2694 818 2746
rect 870 2694 882 2746
rect 934 2694 946 2746
rect 998 2694 1010 2746
rect 1062 2694 1080 2746
rect 800 2036 1080 2694
rect 1306 2680 1362 2689
rect 1306 2615 1308 2624
rect 1360 2615 1362 2624
rect 1308 2586 1360 2592
rect 1216 2440 1268 2446
rect 1214 2408 1216 2417
rect 1268 2408 1270 2417
rect 1214 2343 1270 2352
rect 800 1980 832 2036
rect 888 1980 912 2036
rect 968 1980 992 2036
rect 1048 1980 1080 2036
rect 800 1956 1080 1980
rect 800 1900 832 1956
rect 888 1900 912 1956
rect 968 1900 992 1956
rect 1048 1900 1080 1956
rect 800 1876 1080 1900
rect 572 1828 624 1834
rect 572 1770 624 1776
rect 800 1820 832 1876
rect 888 1820 912 1876
rect 968 1820 992 1876
rect 1048 1820 1080 1876
rect 584 490 612 1770
rect 664 1760 716 1766
rect 664 1702 716 1708
rect 676 1193 704 1702
rect 800 1658 1080 1820
rect 2680 2202 2960 3238
rect 2680 2150 2698 2202
rect 2750 2150 2762 2202
rect 2814 2150 2826 2202
rect 2878 2150 2890 2202
rect 2942 2150 2960 2202
rect 1216 1760 1268 1766
rect 1216 1702 1268 1708
rect 800 1606 818 1658
rect 870 1606 882 1658
rect 934 1606 946 1658
rect 998 1606 1010 1658
rect 1062 1606 1080 1658
rect 662 1184 718 1193
rect 662 1119 718 1128
rect 800 1040 1080 1606
rect 1124 1420 1176 1426
rect 1124 1362 1176 1368
rect 1136 1329 1164 1362
rect 1122 1320 1178 1329
rect 1122 1255 1178 1264
rect 754 490 810 600
rect 584 462 810 490
rect 754 -600 810 462
rect 1122 490 1178 600
rect 1228 490 1256 1702
rect 1306 1592 1362 1601
rect 1306 1527 1308 1536
rect 1360 1527 1362 1536
rect 1308 1498 1360 1504
rect 2680 1114 2960 2150
rect 2680 1062 2698 1114
rect 2750 1062 2762 1114
rect 2814 1062 2826 1114
rect 2878 1062 2890 1114
rect 2942 1062 2960 1114
rect 2680 1040 2960 1062
rect 1122 462 1256 490
rect 1122 -600 1178 462
<< via2 >>
rect 1122 4004 1178 4040
rect 1122 3984 1124 4004
rect 1124 3984 1176 4004
rect 1176 3984 1178 4004
rect 1306 4276 1362 4312
rect 1306 4256 1308 4276
rect 1308 4256 1360 4276
rect 1360 4256 1362 4276
rect 1306 3732 1362 3768
rect 1306 3712 1308 3732
rect 1308 3712 1360 3732
rect 1360 3712 1362 3732
rect 2712 3460 2768 3516
rect 2792 3460 2848 3516
rect 2872 3460 2928 3516
rect 2712 3380 2768 3436
rect 2792 3380 2848 3436
rect 2872 3380 2928 3436
rect 2712 3300 2768 3356
rect 2792 3300 2848 3356
rect 2872 3300 2928 3356
rect 1122 2916 1178 2952
rect 1122 2896 1124 2916
rect 1124 2896 1176 2916
rect 1176 2896 1178 2916
rect 1306 2644 1362 2680
rect 1306 2624 1308 2644
rect 1308 2624 1360 2644
rect 1360 2624 1362 2644
rect 1214 2388 1216 2408
rect 1216 2388 1268 2408
rect 1268 2388 1270 2408
rect 1214 2352 1270 2388
rect 832 1980 888 2036
rect 912 1980 968 2036
rect 992 1980 1048 2036
rect 832 1900 888 1956
rect 912 1900 968 1956
rect 992 1900 1048 1956
rect 832 1820 888 1876
rect 912 1820 968 1876
rect 992 1820 1048 1876
rect 662 1128 718 1184
rect 1122 1264 1178 1320
rect 1306 1556 1362 1592
rect 1306 1536 1308 1556
rect 1308 1536 1360 1556
rect 1360 1536 1362 1556
<< metal3 >>
rect -600 4314 600 4344
rect 1301 4314 1367 4317
rect -600 4312 1367 4314
rect -600 4256 1306 4312
rect 1362 4256 1367 4312
rect -600 4254 1367 4256
rect -600 4224 600 4254
rect 1301 4251 1367 4254
rect -600 4042 600 4072
rect 1117 4042 1183 4045
rect -600 4040 1183 4042
rect -600 3984 1122 4040
rect 1178 3984 1183 4040
rect -600 3982 1183 3984
rect -600 3952 600 3982
rect 1117 3979 1183 3982
rect -600 3770 600 3800
rect 1301 3770 1367 3773
rect -600 3768 1367 3770
rect -600 3712 1306 3768
rect 1362 3712 1367 3768
rect -600 3710 1367 3712
rect -600 3680 600 3710
rect 1301 3707 1367 3710
rect 412 3516 3268 3548
rect 412 3460 2712 3516
rect 2768 3460 2792 3516
rect 2848 3460 2872 3516
rect 2928 3460 3268 3516
rect 412 3436 3268 3460
rect 412 3380 2712 3436
rect 2768 3380 2792 3436
rect 2848 3380 2872 3436
rect 2928 3380 3268 3436
rect 412 3356 3268 3380
rect 412 3300 2712 3356
rect 2768 3300 2792 3356
rect 2848 3300 2872 3356
rect 2928 3300 3268 3356
rect 412 3268 3268 3300
rect -600 2954 600 2984
rect 1117 2954 1183 2957
rect -600 2952 1183 2954
rect -600 2896 1122 2952
rect 1178 2896 1183 2952
rect -600 2894 1183 2896
rect -600 2864 600 2894
rect 1117 2891 1183 2894
rect -600 2682 600 2712
rect 1301 2682 1367 2685
rect -600 2680 1367 2682
rect -600 2624 1306 2680
rect 1362 2624 1367 2680
rect -600 2622 1367 2624
rect -600 2592 600 2622
rect 1301 2619 1367 2622
rect -600 2410 600 2440
rect 1209 2410 1275 2413
rect -600 2408 1275 2410
rect -600 2352 1214 2408
rect 1270 2352 1275 2408
rect -600 2350 1275 2352
rect -600 2320 600 2350
rect 1209 2347 1275 2350
rect 412 2036 3268 2068
rect 412 1980 832 2036
rect 888 1980 912 2036
rect 968 1980 992 2036
rect 1048 1980 3268 2036
rect 412 1956 3268 1980
rect 412 1900 832 1956
rect 888 1900 912 1956
rect 968 1900 992 1956
rect 1048 1900 3268 1956
rect 412 1876 3268 1900
rect 412 1820 832 1876
rect 888 1820 912 1876
rect 968 1820 992 1876
rect 1048 1820 3268 1876
rect 412 1788 3268 1820
rect -600 1594 600 1624
rect 1301 1594 1367 1597
rect -600 1592 1367 1594
rect -600 1536 1306 1592
rect 1362 1536 1367 1592
rect -600 1534 1367 1536
rect -600 1504 600 1534
rect 1301 1531 1367 1534
rect -600 1322 600 1352
rect 1117 1322 1183 1325
rect -600 1320 1183 1322
rect -600 1264 1122 1320
rect 1178 1264 1183 1320
rect -600 1262 1183 1264
rect -600 1232 600 1262
rect 1117 1259 1183 1262
rect 657 1186 723 1189
rect 657 1184 858 1186
rect 657 1128 662 1184
rect 718 1128 858 1184
rect 657 1126 858 1128
rect 657 1123 723 1126
rect -600 1050 600 1080
rect 798 1050 858 1126
rect -600 990 858 1050
rect -600 960 600 990
use sky130_fd_sc_hd__fill_2  FILLER_0_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1196 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1673029049
transform 1 0 1840 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2116 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2852 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1673029049
transform 1 0 736 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1673029049
transform 1 0 1196 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1673029049
transform 1 0 1840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1673029049
transform 1 0 2484 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_26
timestamp 1673029049
transform 1 0 2852 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1673029049
transform 1 0 736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_14 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1673029049
transform 1 0 2116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1673029049
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 736 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1673029049
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp 1673029049
transform 1 0 2208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1673029049
transform 1 0 736 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp 1673029049
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1673029049
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1673029049
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1673029049
transform 1 0 736 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1673029049
transform 1 0 1196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1673029049
transform 1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_18
timestamp 1673029049
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1673029049
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 3220 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1673029049
transform 1 0 2024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1673029049
transform 1 0 2024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1673029049
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[1\]
timestamp 1673029049
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[2\]
timestamp 1673029049
transform -1 0 1196 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[3\]
timestamp 1673029049
transform -1 0 1196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[4\]
timestamp 1673029049
transform -1 0 1840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[5\]
timestamp 1673029049
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[6\]
timestamp 1673029049
transform -1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[7\]
timestamp 1673029049
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[8\]
timestamp 1673029049
transform -1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[9\]
timestamp 1673029049
transform -1 0 1196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[10\]
timestamp 1673029049
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[11\]
timestamp 1673029049
transform -1 0 2484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[12\]
timestamp 1673029049
transform -1 0 1840 0 -1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 2680 1040 2960 4400 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 412 3268 3268 3548 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 800 1040 1080 4400 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 412 1788 3268 2068 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 754 5000 810 6200 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 2 nsew signal tristate
flabel metal3 s -600 4224 600 4344 0 FreeSans 480 0 0 0 gpio_defaults[10]
port 3 nsew signal tristate
flabel metal2 s 754 -600 810 600 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 4 nsew signal tristate
flabel metal2 s 1122 -600 1178 600 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 5 nsew signal tristate
flabel metal2 s 1122 5000 1178 6200 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 6 nsew signal tristate
flabel metal3 s -600 960 600 1080 0 FreeSans 480 0 0 0 gpio_defaults[2]
port 7 nsew signal tristate
flabel metal3 s -600 1232 600 1352 0 FreeSans 480 0 0 0 gpio_defaults[3]
port 8 nsew signal tristate
flabel metal3 s -600 1504 600 1624 0 FreeSans 480 0 0 0 gpio_defaults[4]
port 9 nsew signal tristate
flabel metal3 s -600 2320 600 2440 0 FreeSans 480 0 0 0 gpio_defaults[5]
port 10 nsew signal tristate
flabel metal3 s -600 2592 600 2712 0 FreeSans 480 0 0 0 gpio_defaults[6]
port 11 nsew signal tristate
flabel metal3 s -600 2864 600 2984 0 FreeSans 480 0 0 0 gpio_defaults[7]
port 12 nsew signal tristate
flabel metal3 s -600 3680 600 3800 0 FreeSans 480 0 0 0 gpio_defaults[8]
port 13 nsew signal tristate
flabel metal3 s -600 3952 600 4072 0 FreeSans 480 0 0 0 gpio_defaults[9]
port 14 nsew signal tristate
rlabel metal1 1840 4352 1840 4352 0 VGND
rlabel metal1 1840 3808 1840 3808 0 VPWR
rlabel metal1 1472 4250 1472 4250 0 gpio_defaults_high\[10\]
rlabel metal1 1472 3570 1472 3570 0 gpio_defaults_high\[1\]
rlabel metal1 1012 3026 1012 3026 0 gpio_defaults_low\[0\]
rlabel metal2 683 476 683 476 0 gpio_defaults_low\[11\]
rlabel metal2 1203 476 1203 476 0 gpio_defaults_low\[12\]
rlabel metal3 659 1020 659 1020 0 gpio_defaults_low\[2\]
rlabel metal3 820 1292 820 1292 0 gpio_defaults_low\[3\]
rlabel metal1 1472 1530 1472 1530 0 gpio_defaults_low\[4\]
rlabel metal3 866 2380 866 2380 0 gpio_defaults_low\[5\]
rlabel metal1 1426 2618 1426 2618 0 gpio_defaults_low\[6\]
rlabel metal3 820 2924 820 2924 0 gpio_defaults_low\[7\]
rlabel metal1 1840 3706 1840 3706 0 gpio_defaults_low\[8\]
rlabel metal3 820 4012 820 4012 0 gpio_defaults_low\[9\]
<< properties >>
string FIXED_BBOX 0 0 3400 5600
<< end >>
