magic
tech sky130A
magscale 1 2
timestamp 1665362231
<< nwell >>
rect 1066 29637 378894 30203
rect 1066 28549 378894 29115
rect 1066 27461 378894 28027
rect 1066 26373 378894 26939
rect 1066 25285 378894 25851
rect 1066 24197 378894 24763
rect 1066 23109 378894 23675
rect 1066 22021 378894 22587
rect 1066 20933 378894 21499
rect 1066 19845 378894 20411
rect 1066 18757 378894 19323
rect 1066 17669 378894 18235
rect 1066 16581 378894 17147
rect 1066 15493 133714 16059
rect 1066 14405 133714 14971
rect 1066 13317 133714 13883
rect 1066 12229 133714 12795
rect 1066 11386 133714 11707
rect 1066 11141 64070 11386
rect 1066 10053 64070 10619
rect 1066 8965 64070 9531
rect 1066 7877 64070 8443
rect 1066 6789 64070 7355
rect 1066 5701 64070 6267
rect 1066 4613 378894 5179
rect 1066 3525 378894 4091
rect 1066 2437 378894 3003
rect 1066 1349 378894 1915
<< obsli1 >>
rect 1104 1071 378856 30481
<< obsm1 >>
rect 26206 32000 142384 32008
rect 144886 32000 147674 32008
rect 1104 8 378856 32000
<< metal2 >>
rect 8482 31200 8538 32400
rect 9218 31200 9274 32400
rect 9954 31200 10010 32400
rect 10690 31200 10746 32400
rect 11426 31200 11482 32400
rect 12162 31200 12218 32400
rect 12898 31200 12954 32400
rect 13634 31200 13690 32400
rect 14370 31200 14426 32400
rect 15106 31200 15162 32400
rect 15842 31200 15898 32400
rect 16578 31200 16634 32400
rect 17314 31200 17370 32400
rect 18050 31200 18106 32400
rect 18786 31200 18842 32400
rect 19522 31200 19578 32400
rect 20258 31200 20314 32400
rect 20994 31200 21050 32400
rect 21730 31200 21786 32400
rect 22466 31200 22522 32400
rect 23202 31200 23258 32400
rect 23938 31200 23994 32400
rect 24674 31200 24730 32400
rect 25410 31200 25466 32400
rect 26146 31200 26202 32400
rect 26882 31200 26938 32400
rect 27618 31200 27674 32400
rect 28354 31200 28410 32400
rect 29090 31200 29146 32400
rect 29826 31200 29882 32400
rect 30562 31200 30618 32400
rect 31298 31200 31354 32400
rect 32034 31200 32090 32400
rect 32770 31200 32826 32400
rect 33506 31200 33562 32400
rect 34242 31200 34298 32400
rect 34978 31200 35034 32400
rect 35714 31200 35770 32400
rect 36450 31200 36506 32400
rect 37186 31200 37242 32400
rect 37922 31200 37978 32400
rect 38658 31200 38714 32400
rect 39394 31200 39450 32400
rect 40130 31200 40186 32400
rect 40866 31200 40922 32400
rect 41602 31200 41658 32400
rect 42338 31200 42394 32400
rect 43074 31200 43130 32400
rect 43810 31200 43866 32400
rect 44546 31200 44602 32400
rect 45282 31200 45338 32400
rect 46018 31200 46074 32400
rect 46754 31200 46810 32400
rect 47490 31200 47546 32400
rect 48226 31200 48282 32400
rect 48962 31200 49018 32400
rect 49698 31200 49754 32400
rect 50434 31200 50490 32400
rect 51170 31200 51226 32400
rect 51906 31200 51962 32400
rect 52642 31200 52698 32400
rect 53378 31200 53434 32400
rect 54114 31200 54170 32400
rect 54850 31200 54906 32400
rect 55586 31200 55642 32400
rect 56322 31200 56378 32400
rect 57058 31200 57114 32400
rect 57794 31200 57850 32400
rect 58530 31200 58586 32400
rect 59266 31200 59322 32400
rect 60002 31200 60058 32400
rect 60738 31200 60794 32400
rect 61474 31200 61530 32400
rect 62210 31200 62266 32400
rect 62946 31200 63002 32400
rect 63682 31200 63738 32400
rect 64418 31200 64474 32400
rect 65154 31200 65210 32400
rect 65890 31200 65946 32400
rect 66626 31200 66682 32400
rect 67362 31200 67418 32400
rect 68098 31200 68154 32400
rect 68834 31200 68890 32400
rect 69570 31200 69626 32400
rect 70306 31200 70362 32400
rect 71042 31200 71098 32400
rect 71778 31200 71834 32400
rect 72514 31200 72570 32400
rect 73250 31200 73306 32400
rect 73986 31200 74042 32400
rect 74722 31200 74778 32400
rect 75458 31200 75514 32400
rect 76194 31200 76250 32400
rect 76930 31200 76986 32400
rect 77666 31200 77722 32400
rect 78402 31200 78458 32400
rect 79138 31200 79194 32400
rect 79874 31200 79930 32400
rect 80610 31200 80666 32400
rect 81346 31200 81402 32400
rect 82082 31200 82138 32400
rect 82818 31200 82874 32400
rect 83554 31200 83610 32400
rect 84290 31200 84346 32400
rect 85026 31200 85082 32400
rect 85762 31200 85818 32400
rect 86498 31200 86554 32400
rect 87234 31200 87290 32400
rect 87970 31200 88026 32400
rect 88706 31200 88762 32400
rect 89442 31200 89498 32400
rect 90178 31200 90234 32400
rect 90914 31200 90970 32400
rect 91650 31200 91706 32400
rect 92386 31200 92442 32400
rect 93122 31200 93178 32400
rect 93858 31200 93914 32400
rect 94594 31200 94650 32400
rect 95330 31200 95386 32400
rect 96066 31200 96122 32400
rect 96802 31200 96858 32400
rect 97538 31200 97594 32400
rect 98274 31200 98330 32400
rect 99010 31200 99066 32400
rect 99746 31200 99802 32400
rect 100482 31200 100538 32400
rect 101218 31200 101274 32400
rect 101954 31200 102010 32400
rect 102690 31200 102746 32400
rect 103426 31200 103482 32400
rect 104162 31200 104218 32400
rect 104898 31200 104954 32400
rect 105634 31200 105690 32400
rect 106370 31200 106426 32400
rect 107106 31200 107162 32400
rect 107842 31200 107898 32400
rect 108578 31200 108634 32400
rect 109314 31200 109370 32400
rect 110050 31200 110106 32400
rect 110786 31200 110842 32400
rect 111522 31200 111578 32400
rect 112258 31200 112314 32400
rect 112994 31200 113050 32400
rect 113730 31200 113786 32400
rect 114466 31200 114522 32400
rect 115202 31200 115258 32400
rect 115938 31200 115994 32400
rect 116674 31200 116730 32400
rect 117410 31200 117466 32400
rect 118146 31200 118202 32400
rect 118882 31200 118938 32400
rect 119618 31200 119674 32400
rect 120354 31200 120410 32400
rect 121090 31200 121146 32400
rect 121826 31200 121882 32400
rect 122562 31200 122618 32400
rect 123298 31200 123354 32400
rect 124034 31200 124090 32400
rect 124770 31200 124826 32400
rect 125506 31200 125562 32400
rect 126242 31200 126298 32400
rect 126978 31200 127034 32400
rect 127714 31200 127770 32400
rect 128450 31200 128506 32400
rect 129186 31200 129242 32400
rect 129922 31200 129978 32400
rect 130658 31200 130714 32400
rect 131394 31200 131450 32400
rect 132130 31200 132186 32400
rect 132866 31200 132922 32400
rect 133602 31200 133658 32400
rect 134338 31200 134394 32400
rect 135074 31200 135130 32400
rect 135810 31200 135866 32400
rect 136546 31200 136602 32400
rect 137282 31200 137338 32400
rect 138018 31200 138074 32400
rect 138754 31200 138810 32400
rect 139490 31200 139546 32400
rect 140226 31200 140282 32400
rect 140962 31200 141018 32400
rect 141698 31200 141754 32400
rect 142434 31200 142490 32400
rect 143170 31200 143226 32400
rect 143906 31200 143962 32400
rect 144642 31200 144698 32400
rect 145378 31200 145434 32400
rect 146114 31200 146170 32400
rect 146850 31200 146906 32400
rect 147586 31200 147642 32400
rect 148322 31200 148378 32400
rect 149058 31200 149114 32400
rect 149794 31200 149850 32400
rect 150530 31200 150586 32400
rect 151266 31200 151322 32400
rect 152002 31200 152058 32400
rect 152738 31200 152794 32400
rect 153474 31200 153530 32400
rect 154210 31200 154266 32400
rect 154946 31200 155002 32400
rect 155682 31200 155738 32400
rect 156418 31200 156474 32400
rect 157154 31200 157210 32400
rect 157890 31200 157946 32400
rect 158626 31200 158682 32400
rect 159362 31200 159418 32400
rect 160098 31200 160154 32400
rect 160834 31200 160890 32400
rect 161570 31200 161626 32400
rect 162306 31200 162362 32400
rect 163042 31200 163098 32400
rect 163778 31200 163834 32400
rect 164514 31200 164570 32400
rect 165250 31200 165306 32400
rect 165986 31200 166042 32400
rect 166722 31200 166778 32400
rect 167458 31200 167514 32400
rect 168194 31200 168250 32400
rect 168930 31200 168986 32400
rect 169666 31200 169722 32400
rect 170402 31200 170458 32400
rect 171138 31200 171194 32400
rect 171874 31200 171930 32400
rect 172610 31200 172666 32400
rect 173346 31200 173402 32400
rect 174082 31200 174138 32400
rect 174818 31200 174874 32400
rect 175554 31200 175610 32400
rect 176290 31200 176346 32400
rect 177026 31200 177082 32400
rect 177762 31200 177818 32400
rect 178498 31200 178554 32400
rect 179234 31200 179290 32400
rect 179970 31200 180026 32400
rect 180706 31200 180762 32400
rect 181442 31200 181498 32400
rect 182178 31200 182234 32400
rect 182914 31200 182970 32400
rect 183650 31200 183706 32400
rect 184386 31200 184442 32400
rect 185122 31200 185178 32400
rect 185858 31200 185914 32400
rect 186594 31200 186650 32400
rect 187330 31200 187386 32400
rect 188066 31200 188122 32400
rect 188802 31200 188858 32400
rect 189538 31200 189594 32400
rect 190274 31200 190330 32400
rect 191010 31200 191066 32400
rect 191746 31200 191802 32400
rect 192482 31200 192538 32400
rect 193218 31200 193274 32400
rect 193954 31200 194010 32400
rect 194690 31200 194746 32400
rect 195426 31200 195482 32400
rect 196162 31200 196218 32400
rect 196898 31200 196954 32400
rect 197634 31200 197690 32400
rect 198370 31200 198426 32400
rect 199106 31200 199162 32400
rect 199842 31200 199898 32400
rect 200578 31200 200634 32400
rect 201314 31200 201370 32400
rect 202050 31200 202106 32400
rect 202786 31200 202842 32400
rect 203522 31200 203578 32400
rect 204258 31200 204314 32400
rect 204994 31200 205050 32400
rect 205730 31200 205786 32400
rect 206466 31200 206522 32400
rect 207202 31200 207258 32400
rect 207938 31200 207994 32400
rect 208674 31200 208730 32400
rect 209410 31200 209466 32400
rect 210146 31200 210202 32400
rect 210882 31200 210938 32400
rect 211618 31200 211674 32400
rect 212354 31200 212410 32400
rect 213090 31200 213146 32400
rect 213826 31200 213882 32400
rect 214562 31200 214618 32400
rect 215298 31200 215354 32400
rect 216034 31200 216090 32400
rect 216770 31200 216826 32400
rect 217506 31200 217562 32400
rect 218242 31200 218298 32400
rect 218978 31200 219034 32400
rect 219714 31200 219770 32400
rect 220450 31200 220506 32400
rect 221186 31200 221242 32400
rect 221922 31200 221978 32400
rect 222658 31200 222714 32400
rect 223394 31200 223450 32400
rect 224130 31200 224186 32400
rect 224866 31200 224922 32400
rect 225602 31200 225658 32400
rect 226338 31200 226394 32400
rect 227074 31200 227130 32400
rect 227810 31200 227866 32400
rect 228546 31200 228602 32400
rect 229282 31200 229338 32400
rect 230018 31200 230074 32400
rect 230754 31200 230810 32400
rect 231490 31200 231546 32400
rect 232226 31200 232282 32400
rect 232962 31200 233018 32400
rect 233698 31200 233754 32400
rect 234434 31200 234490 32400
rect 235170 31200 235226 32400
rect 235906 31200 235962 32400
rect 236642 31200 236698 32400
rect 237378 31200 237434 32400
rect 238114 31200 238170 32400
rect 238850 31200 238906 32400
rect 239586 31200 239642 32400
rect 240322 31200 240378 32400
rect 241058 31200 241114 32400
rect 241794 31200 241850 32400
rect 242530 31200 242586 32400
rect 243266 31200 243322 32400
rect 244002 31200 244058 32400
rect 244738 31200 244794 32400
rect 245474 31200 245530 32400
rect 246210 31200 246266 32400
rect 246946 31200 247002 32400
rect 247682 31200 247738 32400
rect 248418 31200 248474 32400
rect 249154 31200 249210 32400
rect 249890 31200 249946 32400
rect 250626 31200 250682 32400
rect 251362 31200 251418 32400
rect 252098 31200 252154 32400
rect 252834 31200 252890 32400
rect 253570 31200 253626 32400
rect 254306 31200 254362 32400
rect 255042 31200 255098 32400
rect 255778 31200 255834 32400
rect 256514 31200 256570 32400
rect 257250 31200 257306 32400
rect 257986 31200 258042 32400
rect 258722 31200 258778 32400
rect 259458 31200 259514 32400
rect 260194 31200 260250 32400
rect 260930 31200 260986 32400
rect 261666 31200 261722 32400
rect 262402 31200 262458 32400
rect 263138 31200 263194 32400
rect 263874 31200 263930 32400
rect 264610 31200 264666 32400
rect 265346 31200 265402 32400
rect 266082 31200 266138 32400
rect 266818 31200 266874 32400
rect 267554 31200 267610 32400
rect 268290 31200 268346 32400
rect 269026 31200 269082 32400
rect 269762 31200 269818 32400
rect 270498 31200 270554 32400
rect 271234 31200 271290 32400
rect 271970 31200 272026 32400
rect 272706 31200 272762 32400
rect 273442 31200 273498 32400
rect 274178 31200 274234 32400
rect 274914 31200 274970 32400
rect 275650 31200 275706 32400
rect 276386 31200 276442 32400
rect 277122 31200 277178 32400
rect 277858 31200 277914 32400
rect 278594 31200 278650 32400
rect 279330 31200 279386 32400
rect 280066 31200 280122 32400
rect 280802 31200 280858 32400
rect 281538 31200 281594 32400
rect 282274 31200 282330 32400
rect 283010 31200 283066 32400
rect 283746 31200 283802 32400
rect 284482 31200 284538 32400
rect 285218 31200 285274 32400
rect 285954 31200 286010 32400
rect 286690 31200 286746 32400
rect 287426 31200 287482 32400
rect 288162 31200 288218 32400
rect 288898 31200 288954 32400
rect 289634 31200 289690 32400
rect 290370 31200 290426 32400
rect 291106 31200 291162 32400
rect 291842 31200 291898 32400
rect 292578 31200 292634 32400
rect 293314 31200 293370 32400
rect 294050 31200 294106 32400
rect 294786 31200 294842 32400
rect 295522 31200 295578 32400
rect 296258 31200 296314 32400
rect 296994 31200 297050 32400
rect 297730 31200 297786 32400
rect 298466 31200 298522 32400
rect 299202 31200 299258 32400
rect 299938 31200 299994 32400
rect 300674 31200 300730 32400
rect 301410 31200 301466 32400
rect 302146 31200 302202 32400
rect 302882 31200 302938 32400
rect 303618 31200 303674 32400
rect 304354 31200 304410 32400
rect 305090 31200 305146 32400
rect 305826 31200 305882 32400
rect 306562 31200 306618 32400
rect 307298 31200 307354 32400
rect 308034 31200 308090 32400
rect 308770 31200 308826 32400
rect 309506 31200 309562 32400
rect 310242 31200 310298 32400
rect 310978 31200 311034 32400
rect 311714 31200 311770 32400
rect 312450 31200 312506 32400
rect 313186 31200 313242 32400
rect 313922 31200 313978 32400
rect 314658 31200 314714 32400
rect 315394 31200 315450 32400
rect 316130 31200 316186 32400
rect 316866 31200 316922 32400
rect 317602 31200 317658 32400
rect 318338 31200 318394 32400
rect 319074 31200 319130 32400
rect 319810 31200 319866 32400
rect 320546 31200 320602 32400
rect 321282 31200 321338 32400
rect 322018 31200 322074 32400
rect 322754 31200 322810 32400
rect 323490 31200 323546 32400
rect 324226 31200 324282 32400
rect 324962 31200 325018 32400
rect 325698 31200 325754 32400
rect 326434 31200 326490 32400
rect 327170 31200 327226 32400
rect 327906 31200 327962 32400
rect 328642 31200 328698 32400
rect 329378 31200 329434 32400
rect 330114 31200 330170 32400
rect 330850 31200 330906 32400
rect 331586 31200 331642 32400
rect 332322 31200 332378 32400
rect 333058 31200 333114 32400
rect 333794 31200 333850 32400
rect 334530 31200 334586 32400
rect 335266 31200 335322 32400
rect 336002 31200 336058 32400
rect 336738 31200 336794 32400
rect 337474 31200 337530 32400
rect 338210 31200 338266 32400
rect 338946 31200 339002 32400
rect 339682 31200 339738 32400
rect 340418 31200 340474 32400
rect 341154 31200 341210 32400
rect 341890 31200 341946 32400
rect 342626 31200 342682 32400
rect 343362 31200 343418 32400
rect 344098 31200 344154 32400
rect 344834 31200 344890 32400
rect 345570 31200 345626 32400
rect 346306 31200 346362 32400
rect 347042 31200 347098 32400
rect 347778 31200 347834 32400
rect 348514 31200 348570 32400
rect 349250 31200 349306 32400
rect 349986 31200 350042 32400
rect 350722 31200 350778 32400
rect 351458 31200 351514 32400
rect 352194 31200 352250 32400
rect 352930 31200 352986 32400
rect 353666 31200 353722 32400
rect 354402 31200 354458 32400
rect 355138 31200 355194 32400
rect 355874 31200 355930 32400
rect 356610 31200 356666 32400
rect 357346 31200 357402 32400
rect 358082 31200 358138 32400
rect 358818 31200 358874 32400
rect 359554 31200 359610 32400
rect 360290 31200 360346 32400
rect 361026 31200 361082 32400
rect 361762 31200 361818 32400
rect 362498 31200 362554 32400
rect 363234 31200 363290 32400
rect 363970 31200 364026 32400
rect 364706 31200 364762 32400
rect 365442 31200 365498 32400
rect 366178 31200 366234 32400
rect 366914 31200 366970 32400
rect 367650 31200 367706 32400
rect 368386 31200 368442 32400
rect 369122 31200 369178 32400
rect 369858 31200 369914 32400
rect 370594 31200 370650 32400
rect 371330 31200 371386 32400
rect 19890 -400 19946 800
rect 20442 -400 20498 800
rect 20994 -400 21050 800
rect 21546 -400 21602 800
rect 22098 -400 22154 800
rect 22650 -400 22706 800
rect 23202 -400 23258 800
rect 23754 -400 23810 800
rect 24306 -400 24362 800
rect 24858 -400 24914 800
rect 25410 -400 25466 800
rect 25962 -400 26018 800
rect 26514 -400 26570 800
rect 27066 -400 27122 800
rect 27618 -400 27674 800
rect 28170 -400 28226 800
rect 28722 -400 28778 800
rect 29274 -400 29330 800
rect 29826 -400 29882 800
rect 30378 -400 30434 800
rect 30930 -400 30986 800
rect 31482 -400 31538 800
rect 32034 -400 32090 800
rect 32586 -400 32642 800
rect 33138 -400 33194 800
rect 33690 -400 33746 800
rect 34242 -400 34298 800
rect 34794 -400 34850 800
rect 35346 -400 35402 800
rect 35898 -400 35954 800
rect 36450 -400 36506 800
rect 37002 -400 37058 800
rect 37554 -400 37610 800
rect 38106 -400 38162 800
rect 38658 -400 38714 800
rect 39210 -400 39266 800
rect 39762 -400 39818 800
rect 40314 -400 40370 800
rect 40866 -400 40922 800
rect 41418 -400 41474 800
rect 41970 -400 42026 800
rect 42522 -400 42578 800
rect 43074 -400 43130 800
rect 43626 -400 43682 800
rect 44178 -400 44234 800
rect 44730 -400 44786 800
rect 45282 -400 45338 800
rect 45834 -400 45890 800
rect 46386 -400 46442 800
rect 46938 -400 46994 800
rect 47490 -400 47546 800
rect 48042 -400 48098 800
rect 48594 -400 48650 800
rect 49146 -400 49202 800
rect 49698 -400 49754 800
rect 50250 -400 50306 800
rect 50802 -400 50858 800
rect 51354 -400 51410 800
rect 51906 -400 51962 800
rect 52458 -400 52514 800
rect 53010 -400 53066 800
rect 53562 -400 53618 800
rect 54114 -400 54170 800
rect 54666 -400 54722 800
rect 55218 -400 55274 800
rect 55770 -400 55826 800
rect 56322 -400 56378 800
rect 56874 -400 56930 800
rect 57426 -400 57482 800
rect 57978 -400 58034 800
rect 58530 -400 58586 800
rect 59082 -400 59138 800
rect 59634 -400 59690 800
rect 60186 -400 60242 800
rect 60738 -400 60794 800
rect 61290 -400 61346 800
rect 61842 -400 61898 800
rect 62394 -400 62450 800
rect 62946 -400 63002 800
rect 63498 -400 63554 800
rect 64050 -400 64106 800
rect 64602 -400 64658 800
rect 65154 -400 65210 800
rect 65706 -400 65762 800
rect 66258 -400 66314 800
rect 66810 -400 66866 800
rect 67362 -400 67418 800
rect 67914 -400 67970 800
rect 68466 -400 68522 800
rect 69018 -400 69074 800
rect 69570 -400 69626 800
rect 70122 -400 70178 800
rect 70674 -400 70730 800
rect 71226 -400 71282 800
rect 71778 -400 71834 800
rect 72330 -400 72386 800
rect 72882 -400 72938 800
rect 73434 -400 73490 800
rect 73986 -400 74042 800
rect 74538 -400 74594 800
rect 75090 -400 75146 800
rect 75642 -400 75698 800
rect 76194 -400 76250 800
rect 76746 -400 76802 800
rect 77298 -400 77354 800
rect 77850 -400 77906 800
rect 78402 -400 78458 800
rect 78954 -400 79010 800
rect 79506 -400 79562 800
rect 80058 -400 80114 800
rect 80610 -400 80666 800
rect 81162 -400 81218 800
rect 81714 -400 81770 800
rect 82266 -400 82322 800
rect 82818 -400 82874 800
rect 83370 -400 83426 800
rect 83922 -400 83978 800
rect 84474 -400 84530 800
rect 85026 -400 85082 800
rect 85578 -400 85634 800
rect 86130 -400 86186 800
rect 86682 -400 86738 800
rect 87234 -400 87290 800
rect 87786 -400 87842 800
rect 88338 -400 88394 800
rect 88890 -400 88946 800
rect 89442 -400 89498 800
rect 89994 -400 90050 800
rect 90546 -400 90602 800
rect 91098 -400 91154 800
rect 91650 -400 91706 800
rect 92202 -400 92258 800
rect 92754 -400 92810 800
rect 93306 -400 93362 800
rect 93858 -400 93914 800
rect 94410 -400 94466 800
rect 94962 -400 95018 800
rect 95514 -400 95570 800
rect 96066 -400 96122 800
rect 96618 -400 96674 800
rect 97170 -400 97226 800
rect 97722 -400 97778 800
rect 98274 -400 98330 800
rect 98826 -400 98882 800
rect 99378 -400 99434 800
rect 99930 -400 99986 800
rect 100482 -400 100538 800
rect 101034 -400 101090 800
rect 101586 -400 101642 800
rect 102138 -400 102194 800
rect 102690 -400 102746 800
rect 103242 -400 103298 800
rect 103794 -400 103850 800
rect 104346 -400 104402 800
rect 104898 -400 104954 800
rect 105450 -400 105506 800
rect 106002 -400 106058 800
rect 106554 -400 106610 800
rect 107106 -400 107162 800
rect 107658 -400 107714 800
rect 108210 -400 108266 800
rect 108762 -400 108818 800
rect 109314 -400 109370 800
rect 109866 -400 109922 800
rect 110418 -400 110474 800
rect 110970 -400 111026 800
rect 111522 -400 111578 800
rect 112074 -400 112130 800
rect 112626 -400 112682 800
rect 113178 -400 113234 800
rect 113730 -400 113786 800
rect 114282 -400 114338 800
rect 114834 -400 114890 800
rect 115386 -400 115442 800
rect 115938 -400 115994 800
rect 116490 -400 116546 800
rect 117042 -400 117098 800
rect 117594 -400 117650 800
rect 118146 -400 118202 800
rect 118698 -400 118754 800
rect 119250 -400 119306 800
rect 119802 -400 119858 800
rect 120354 -400 120410 800
rect 120906 -400 120962 800
rect 121458 -400 121514 800
rect 122010 -400 122066 800
rect 122562 -400 122618 800
rect 123114 -400 123170 800
rect 123666 -400 123722 800
rect 124218 -400 124274 800
rect 124770 -400 124826 800
rect 125322 -400 125378 800
rect 125874 -400 125930 800
rect 126426 -400 126482 800
rect 126978 -400 127034 800
rect 127530 -400 127586 800
rect 128082 -400 128138 800
rect 128634 -400 128690 800
rect 129186 -400 129242 800
rect 129738 -400 129794 800
rect 130290 -400 130346 800
rect 130842 -400 130898 800
rect 131394 -400 131450 800
rect 131946 -400 132002 800
rect 132498 -400 132554 800
rect 133050 -400 133106 800
rect 133602 -400 133658 800
rect 134154 -400 134210 800
rect 134706 -400 134762 800
rect 135258 -400 135314 800
rect 135810 -400 135866 800
rect 136362 -400 136418 800
rect 136914 -400 136970 800
rect 137466 -400 137522 800
rect 138018 -400 138074 800
rect 138570 -400 138626 800
rect 139122 -400 139178 800
rect 139674 -400 139730 800
rect 140226 -400 140282 800
rect 140778 -400 140834 800
rect 141330 -400 141386 800
rect 141882 -400 141938 800
rect 142434 -400 142490 800
rect 142986 -400 143042 800
rect 143538 -400 143594 800
rect 144090 -400 144146 800
rect 144642 -400 144698 800
rect 145194 -400 145250 800
rect 145746 -400 145802 800
rect 146298 -400 146354 800
rect 146850 -400 146906 800
rect 147402 -400 147458 800
rect 147954 -400 148010 800
rect 148506 -400 148562 800
rect 149058 -400 149114 800
rect 149610 -400 149666 800
rect 150162 -400 150218 800
rect 150714 -400 150770 800
rect 151266 -400 151322 800
rect 151818 -400 151874 800
rect 152370 -400 152426 800
rect 152922 -400 152978 800
rect 153474 -400 153530 800
rect 154026 -400 154082 800
rect 154578 -400 154634 800
rect 155130 -400 155186 800
rect 155682 -400 155738 800
rect 156234 -400 156290 800
rect 156786 -400 156842 800
rect 157338 -400 157394 800
rect 157890 -400 157946 800
rect 158442 -400 158498 800
rect 158994 -400 159050 800
rect 159546 -400 159602 800
rect 160098 -400 160154 800
rect 160650 -400 160706 800
rect 161202 -400 161258 800
rect 161754 -400 161810 800
rect 162306 -400 162362 800
rect 162858 -400 162914 800
rect 163410 -400 163466 800
rect 163962 -400 164018 800
rect 164514 -400 164570 800
rect 165066 -400 165122 800
rect 165618 -400 165674 800
rect 166170 -400 166226 800
rect 166722 -400 166778 800
rect 167274 -400 167330 800
rect 167826 -400 167882 800
rect 168378 -400 168434 800
rect 168930 -400 168986 800
rect 169482 -400 169538 800
rect 170034 -400 170090 800
rect 170586 -400 170642 800
rect 171138 -400 171194 800
rect 171690 -400 171746 800
rect 172242 -400 172298 800
rect 172794 -400 172850 800
rect 173346 -400 173402 800
rect 173898 -400 173954 800
rect 174450 -400 174506 800
rect 175002 -400 175058 800
rect 175554 -400 175610 800
rect 176106 -400 176162 800
rect 176658 -400 176714 800
rect 177210 -400 177266 800
rect 177762 -400 177818 800
rect 178314 -400 178370 800
rect 178866 -400 178922 800
rect 179418 -400 179474 800
rect 179970 -400 180026 800
rect 180522 -400 180578 800
rect 181074 -400 181130 800
rect 181626 -400 181682 800
rect 182178 -400 182234 800
rect 182730 -400 182786 800
rect 183282 -400 183338 800
rect 183834 -400 183890 800
rect 184386 -400 184442 800
rect 184938 -400 184994 800
rect 185490 -400 185546 800
rect 186042 -400 186098 800
rect 186594 -400 186650 800
rect 187146 -400 187202 800
rect 187698 -400 187754 800
rect 188250 -400 188306 800
rect 188802 -400 188858 800
rect 189354 -400 189410 800
rect 189906 -400 189962 800
rect 190458 -400 190514 800
rect 191010 -400 191066 800
rect 191562 -400 191618 800
rect 192114 -400 192170 800
rect 192666 -400 192722 800
rect 193218 -400 193274 800
rect 193770 -400 193826 800
rect 194322 -400 194378 800
rect 194874 -400 194930 800
rect 195426 -400 195482 800
rect 195978 -400 196034 800
rect 196530 -400 196586 800
rect 197082 -400 197138 800
rect 197634 -400 197690 800
rect 198186 -400 198242 800
rect 198738 -400 198794 800
rect 199290 -400 199346 800
rect 199842 -400 199898 800
rect 200394 -400 200450 800
rect 200946 -400 201002 800
rect 201498 -400 201554 800
rect 202050 -400 202106 800
rect 202602 -400 202658 800
rect 203154 -400 203210 800
rect 203706 -400 203762 800
rect 204258 -400 204314 800
rect 204810 -400 204866 800
rect 205362 -400 205418 800
rect 205914 -400 205970 800
rect 206466 -400 206522 800
rect 207018 -400 207074 800
rect 207570 -400 207626 800
rect 208122 -400 208178 800
rect 208674 -400 208730 800
rect 209226 -400 209282 800
rect 209778 -400 209834 800
rect 210330 -400 210386 800
rect 210882 -400 210938 800
rect 211434 -400 211490 800
rect 211986 -400 212042 800
rect 212538 -400 212594 800
rect 213090 -400 213146 800
rect 213642 -400 213698 800
rect 214194 -400 214250 800
rect 214746 -400 214802 800
rect 215298 -400 215354 800
rect 215850 -400 215906 800
rect 216402 -400 216458 800
rect 216954 -400 217010 800
rect 217506 -400 217562 800
rect 218058 -400 218114 800
rect 218610 -400 218666 800
rect 219162 -400 219218 800
rect 219714 -400 219770 800
rect 220266 -400 220322 800
rect 220818 -400 220874 800
rect 221370 -400 221426 800
rect 221922 -400 221978 800
rect 222474 -400 222530 800
rect 223026 -400 223082 800
rect 223578 -400 223634 800
rect 224130 -400 224186 800
rect 224682 -400 224738 800
rect 225234 -400 225290 800
rect 225786 -400 225842 800
rect 226338 -400 226394 800
rect 226890 -400 226946 800
rect 227442 -400 227498 800
rect 227994 -400 228050 800
rect 228546 -400 228602 800
rect 229098 -400 229154 800
rect 229650 -400 229706 800
rect 230202 -400 230258 800
rect 230754 -400 230810 800
rect 231306 -400 231362 800
rect 231858 -400 231914 800
rect 232410 -400 232466 800
rect 232962 -400 233018 800
rect 233514 -400 233570 800
rect 234066 -400 234122 800
rect 234618 -400 234674 800
rect 235170 -400 235226 800
rect 235722 -400 235778 800
rect 236274 -400 236330 800
rect 236826 -400 236882 800
rect 237378 -400 237434 800
rect 237930 -400 237986 800
rect 238482 -400 238538 800
rect 239034 -400 239090 800
rect 239586 -400 239642 800
rect 240138 -400 240194 800
rect 240690 -400 240746 800
rect 241242 -400 241298 800
rect 241794 -400 241850 800
rect 242346 -400 242402 800
rect 242898 -400 242954 800
rect 243450 -400 243506 800
rect 244002 -400 244058 800
rect 244554 -400 244610 800
rect 245106 -400 245162 800
rect 245658 -400 245714 800
rect 246210 -400 246266 800
rect 246762 -400 246818 800
rect 247314 -400 247370 800
rect 247866 -400 247922 800
rect 248418 -400 248474 800
rect 248970 -400 249026 800
rect 249522 -400 249578 800
rect 250074 -400 250130 800
rect 250626 -400 250682 800
rect 251178 -400 251234 800
rect 251730 -400 251786 800
rect 252282 -400 252338 800
rect 252834 -400 252890 800
rect 253386 -400 253442 800
rect 253938 -400 253994 800
rect 254490 -400 254546 800
rect 255042 -400 255098 800
rect 255594 -400 255650 800
rect 256146 -400 256202 800
rect 256698 -400 256754 800
rect 257250 -400 257306 800
rect 257802 -400 257858 800
rect 258354 -400 258410 800
rect 258906 -400 258962 800
rect 259458 -400 259514 800
rect 260010 -400 260066 800
rect 260562 -400 260618 800
rect 261114 -400 261170 800
rect 261666 -400 261722 800
rect 262218 -400 262274 800
rect 262770 -400 262826 800
rect 263322 -400 263378 800
rect 263874 -400 263930 800
rect 264426 -400 264482 800
rect 264978 -400 265034 800
rect 265530 -400 265586 800
rect 266082 -400 266138 800
rect 266634 -400 266690 800
rect 267186 -400 267242 800
rect 267738 -400 267794 800
rect 268290 -400 268346 800
rect 268842 -400 268898 800
rect 269394 -400 269450 800
rect 269946 -400 270002 800
rect 270498 -400 270554 800
rect 271050 -400 271106 800
rect 271602 -400 271658 800
rect 272154 -400 272210 800
rect 272706 -400 272762 800
rect 273258 -400 273314 800
rect 273810 -400 273866 800
rect 274362 -400 274418 800
rect 274914 -400 274970 800
rect 275466 -400 275522 800
rect 276018 -400 276074 800
rect 276570 -400 276626 800
rect 277122 -400 277178 800
rect 277674 -400 277730 800
rect 278226 -400 278282 800
rect 278778 -400 278834 800
rect 279330 -400 279386 800
rect 279882 -400 279938 800
rect 280434 -400 280490 800
rect 280986 -400 281042 800
rect 281538 -400 281594 800
rect 282090 -400 282146 800
rect 282642 -400 282698 800
rect 283194 -400 283250 800
rect 283746 -400 283802 800
rect 284298 -400 284354 800
rect 284850 -400 284906 800
rect 285402 -400 285458 800
rect 285954 -400 286010 800
rect 286506 -400 286562 800
rect 287058 -400 287114 800
rect 287610 -400 287666 800
rect 288162 -400 288218 800
rect 288714 -400 288770 800
rect 289266 -400 289322 800
rect 289818 -400 289874 800
rect 290370 -400 290426 800
rect 290922 -400 290978 800
rect 291474 -400 291530 800
rect 292026 -400 292082 800
rect 292578 -400 292634 800
rect 293130 -400 293186 800
rect 293682 -400 293738 800
rect 294234 -400 294290 800
rect 294786 -400 294842 800
rect 295338 -400 295394 800
rect 295890 -400 295946 800
rect 296442 -400 296498 800
rect 296994 -400 297050 800
rect 297546 -400 297602 800
rect 298098 -400 298154 800
rect 298650 -400 298706 800
rect 299202 -400 299258 800
rect 299754 -400 299810 800
rect 300306 -400 300362 800
rect 300858 -400 300914 800
rect 301410 -400 301466 800
rect 301962 -400 302018 800
rect 302514 -400 302570 800
rect 303066 -400 303122 800
rect 303618 -400 303674 800
rect 304170 -400 304226 800
rect 304722 -400 304778 800
rect 305274 -400 305330 800
rect 305826 -400 305882 800
rect 306378 -400 306434 800
rect 306930 -400 306986 800
rect 307482 -400 307538 800
rect 308034 -400 308090 800
rect 308586 -400 308642 800
rect 309138 -400 309194 800
rect 309690 -400 309746 800
rect 310242 -400 310298 800
rect 310794 -400 310850 800
rect 311346 -400 311402 800
rect 311898 -400 311954 800
rect 312450 -400 312506 800
rect 313002 -400 313058 800
rect 313554 -400 313610 800
rect 314106 -400 314162 800
rect 314658 -400 314714 800
rect 315210 -400 315266 800
rect 315762 -400 315818 800
rect 316314 -400 316370 800
rect 316866 -400 316922 800
rect 317418 -400 317474 800
rect 317970 -400 318026 800
rect 318522 -400 318578 800
rect 319074 -400 319130 800
rect 319626 -400 319682 800
rect 320178 -400 320234 800
rect 320730 -400 320786 800
rect 321282 -400 321338 800
rect 321834 -400 321890 800
rect 322386 -400 322442 800
rect 322938 -400 322994 800
rect 323490 -400 323546 800
rect 324042 -400 324098 800
rect 324594 -400 324650 800
rect 325146 -400 325202 800
rect 325698 -400 325754 800
rect 326250 -400 326306 800
rect 326802 -400 326858 800
rect 327354 -400 327410 800
rect 327906 -400 327962 800
rect 328458 -400 328514 800
rect 329010 -400 329066 800
rect 329562 -400 329618 800
rect 330114 -400 330170 800
rect 330666 -400 330722 800
rect 331218 -400 331274 800
rect 331770 -400 331826 800
rect 332322 -400 332378 800
rect 332874 -400 332930 800
rect 333426 -400 333482 800
rect 333978 -400 334034 800
rect 334530 -400 334586 800
rect 335082 -400 335138 800
rect 335634 -400 335690 800
rect 336186 -400 336242 800
rect 336738 -400 336794 800
rect 337290 -400 337346 800
rect 337842 -400 337898 800
rect 338394 -400 338450 800
rect 338946 -400 339002 800
rect 339498 -400 339554 800
rect 340050 -400 340106 800
rect 340602 -400 340658 800
rect 341154 -400 341210 800
rect 341706 -400 341762 800
rect 342258 -400 342314 800
rect 342810 -400 342866 800
rect 343362 -400 343418 800
rect 343914 -400 343970 800
rect 344466 -400 344522 800
rect 345018 -400 345074 800
rect 345570 -400 345626 800
rect 346122 -400 346178 800
rect 346674 -400 346730 800
rect 347226 -400 347282 800
rect 347778 -400 347834 800
rect 348330 -400 348386 800
rect 348882 -400 348938 800
rect 349434 -400 349490 800
rect 349986 -400 350042 800
rect 350538 -400 350594 800
rect 351090 -400 351146 800
rect 351642 -400 351698 800
rect 352194 -400 352250 800
rect 352746 -400 352802 800
rect 353298 -400 353354 800
rect 353850 -400 353906 800
rect 354402 -400 354458 800
rect 354954 -400 355010 800
rect 355506 -400 355562 800
rect 356058 -400 356114 800
rect 356610 -400 356666 800
rect 357162 -400 357218 800
rect 357714 -400 357770 800
rect 358266 -400 358322 800
rect 358818 -400 358874 800
rect 359370 -400 359426 800
rect 359922 -400 359978 800
<< obsm2 >>
rect 5036 31144 8426 31958
rect 8594 31144 9162 31958
rect 9330 31144 9898 31958
rect 10066 31144 10634 31958
rect 10802 31144 11370 31958
rect 11538 31144 12106 31958
rect 12274 31144 12842 31958
rect 13010 31144 13578 31958
rect 13746 31144 14314 31958
rect 14482 31144 15050 31958
rect 15218 31144 15786 31958
rect 15954 31144 16522 31958
rect 16690 31144 17258 31958
rect 17426 31144 17994 31958
rect 18162 31144 18730 31958
rect 18898 31144 19466 31958
rect 19634 31144 20202 31958
rect 20370 31144 20938 31958
rect 21106 31144 21674 31958
rect 21842 31144 22410 31958
rect 22578 31144 23146 31958
rect 23314 31144 23882 31958
rect 24050 31144 24618 31958
rect 24786 31144 25354 31958
rect 25522 31144 26090 31958
rect 26258 31144 26826 31958
rect 26994 31144 27562 31958
rect 27730 31144 28298 31958
rect 28466 31144 29034 31958
rect 29202 31144 29770 31958
rect 29938 31144 30506 31958
rect 30674 31144 31242 31958
rect 31410 31144 31978 31958
rect 32146 31144 32714 31958
rect 32882 31144 33450 31958
rect 33618 31144 34186 31958
rect 34354 31144 34922 31958
rect 35090 31144 35658 31958
rect 35826 31144 36394 31958
rect 36562 31144 37130 31958
rect 37298 31144 37866 31958
rect 38034 31144 38602 31958
rect 38770 31144 39338 31958
rect 39506 31144 40074 31958
rect 40242 31144 40810 31958
rect 40978 31144 41546 31958
rect 41714 31144 42282 31958
rect 42450 31144 43018 31958
rect 43186 31144 43754 31958
rect 43922 31144 44490 31958
rect 44658 31144 45226 31958
rect 45394 31144 45962 31958
rect 46130 31144 46698 31958
rect 46866 31144 47434 31958
rect 47602 31144 48170 31958
rect 48338 31144 48906 31958
rect 49074 31144 49642 31958
rect 49810 31144 50378 31958
rect 50546 31144 51114 31958
rect 51282 31144 51850 31958
rect 52018 31144 52586 31958
rect 52754 31144 53322 31958
rect 53490 31144 54058 31958
rect 54226 31144 54794 31958
rect 54962 31144 55530 31958
rect 55698 31144 56266 31958
rect 56434 31144 57002 31958
rect 57170 31144 57738 31958
rect 57906 31144 58474 31958
rect 58642 31144 59210 31958
rect 59378 31144 59946 31958
rect 60114 31144 60682 31958
rect 60850 31144 61418 31958
rect 61586 31144 62154 31958
rect 62322 31144 62890 31958
rect 63058 31144 63626 31958
rect 63794 31144 64362 31958
rect 64530 31144 65098 31958
rect 65266 31144 65834 31958
rect 66002 31144 66570 31958
rect 66738 31144 67306 31958
rect 67474 31144 68042 31958
rect 68210 31144 68778 31958
rect 68946 31144 69514 31958
rect 69682 31144 70250 31958
rect 70418 31144 70986 31958
rect 71154 31144 71722 31958
rect 71890 31144 72458 31958
rect 72626 31144 73194 31958
rect 73362 31144 73930 31958
rect 74098 31144 74666 31958
rect 74834 31144 75402 31958
rect 75570 31144 76138 31958
rect 76306 31144 76874 31958
rect 77042 31144 77610 31958
rect 77778 31144 78346 31958
rect 78514 31144 79082 31958
rect 79250 31144 79818 31958
rect 79986 31144 80554 31958
rect 80722 31144 81290 31958
rect 81458 31144 82026 31958
rect 82194 31144 82762 31958
rect 82930 31144 83498 31958
rect 83666 31144 84234 31958
rect 84402 31144 84970 31958
rect 85138 31144 85706 31958
rect 85874 31144 86442 31958
rect 86610 31144 87178 31958
rect 87346 31144 87914 31958
rect 88082 31144 88650 31958
rect 88818 31144 89386 31958
rect 89554 31144 90122 31958
rect 90290 31144 90858 31958
rect 91026 31144 91594 31958
rect 91762 31144 92330 31958
rect 92498 31144 93066 31958
rect 93234 31144 93802 31958
rect 93970 31144 94538 31958
rect 94706 31144 95274 31958
rect 95442 31144 96010 31958
rect 96178 31144 96746 31958
rect 96914 31144 97482 31958
rect 97650 31144 98218 31958
rect 98386 31144 98954 31958
rect 99122 31144 99690 31958
rect 99858 31144 100426 31958
rect 100594 31144 101162 31958
rect 101330 31144 101898 31958
rect 102066 31144 102634 31958
rect 102802 31144 103370 31958
rect 103538 31144 104106 31958
rect 104274 31144 104842 31958
rect 105010 31144 105578 31958
rect 105746 31144 106314 31958
rect 106482 31144 107050 31958
rect 107218 31144 107786 31958
rect 107954 31144 108522 31958
rect 108690 31144 109258 31958
rect 109426 31144 109994 31958
rect 110162 31144 110730 31958
rect 110898 31144 111466 31958
rect 111634 31144 112202 31958
rect 112370 31144 112938 31958
rect 113106 31144 113674 31958
rect 113842 31144 114410 31958
rect 114578 31144 115146 31958
rect 115314 31144 115882 31958
rect 116050 31144 116618 31958
rect 116786 31144 117354 31958
rect 117522 31144 118090 31958
rect 118258 31144 118826 31958
rect 118994 31144 119562 31958
rect 119730 31144 120298 31958
rect 120466 31144 121034 31958
rect 121202 31144 121770 31958
rect 121938 31144 122506 31958
rect 122674 31144 123242 31958
rect 123410 31144 123978 31958
rect 124146 31144 124714 31958
rect 124882 31144 125450 31958
rect 125618 31144 126186 31958
rect 126354 31144 126922 31958
rect 127090 31144 127658 31958
rect 127826 31144 128394 31958
rect 128562 31144 129130 31958
rect 129298 31144 129866 31958
rect 130034 31144 130602 31958
rect 130770 31144 131338 31958
rect 131506 31144 132074 31958
rect 132242 31144 132810 31958
rect 132978 31144 133546 31958
rect 133714 31144 134282 31958
rect 134450 31144 135018 31958
rect 135186 31144 135754 31958
rect 135922 31144 136490 31958
rect 136658 31144 137226 31958
rect 137394 31144 137962 31958
rect 138130 31144 138698 31958
rect 138866 31144 139434 31958
rect 139602 31144 140170 31958
rect 140338 31144 140906 31958
rect 141074 31144 141642 31958
rect 141810 31144 142378 31958
rect 142546 31144 143114 31958
rect 143282 31144 143850 31958
rect 144018 31144 144586 31958
rect 144754 31144 145322 31958
rect 145490 31144 146058 31958
rect 146226 31144 146794 31958
rect 146962 31144 147530 31958
rect 147698 31144 148266 31958
rect 148434 31144 149002 31958
rect 149170 31144 149738 31958
rect 149906 31144 150474 31958
rect 150642 31144 151210 31958
rect 151378 31144 151946 31958
rect 152114 31144 152682 31958
rect 152850 31144 153418 31958
rect 153586 31144 154154 31958
rect 154322 31144 154890 31958
rect 155058 31144 155626 31958
rect 155794 31144 156362 31958
rect 156530 31144 157098 31958
rect 157266 31144 157834 31958
rect 158002 31144 158570 31958
rect 158738 31144 159306 31958
rect 159474 31144 160042 31958
rect 160210 31144 160778 31958
rect 160946 31144 161514 31958
rect 161682 31144 162250 31958
rect 162418 31144 162986 31958
rect 163154 31144 163722 31958
rect 163890 31144 164458 31958
rect 164626 31144 165194 31958
rect 165362 31144 165930 31958
rect 166098 31144 166666 31958
rect 166834 31144 167402 31958
rect 167570 31144 168138 31958
rect 168306 31144 168874 31958
rect 169042 31144 169610 31958
rect 169778 31144 170346 31958
rect 170514 31144 171082 31958
rect 171250 31144 171818 31958
rect 171986 31144 172554 31958
rect 172722 31144 173290 31958
rect 173458 31144 174026 31958
rect 174194 31144 174762 31958
rect 174930 31144 175498 31958
rect 175666 31144 176234 31958
rect 176402 31144 176970 31958
rect 177138 31144 177706 31958
rect 177874 31144 178442 31958
rect 178610 31144 179178 31958
rect 179346 31144 179914 31958
rect 180082 31144 180650 31958
rect 180818 31144 181386 31958
rect 181554 31144 182122 31958
rect 182290 31144 182858 31958
rect 183026 31144 183594 31958
rect 183762 31144 184330 31958
rect 184498 31144 185066 31958
rect 185234 31144 185802 31958
rect 185970 31144 186538 31958
rect 186706 31144 187274 31958
rect 187442 31144 188010 31958
rect 188178 31144 188746 31958
rect 188914 31144 189482 31958
rect 189650 31144 190218 31958
rect 190386 31144 190954 31958
rect 191122 31144 191690 31958
rect 191858 31144 192426 31958
rect 192594 31144 193162 31958
rect 193330 31144 193898 31958
rect 194066 31144 194634 31958
rect 194802 31144 195370 31958
rect 195538 31144 196106 31958
rect 196274 31144 196842 31958
rect 197010 31144 197578 31958
rect 197746 31144 198314 31958
rect 198482 31144 199050 31958
rect 199218 31144 199786 31958
rect 199954 31144 200522 31958
rect 200690 31144 201258 31958
rect 201426 31144 201994 31958
rect 202162 31144 202730 31958
rect 202898 31144 203466 31958
rect 203634 31144 204202 31958
rect 204370 31144 204938 31958
rect 205106 31144 205674 31958
rect 205842 31144 206410 31958
rect 206578 31144 207146 31958
rect 207314 31144 207882 31958
rect 208050 31144 208618 31958
rect 208786 31144 209354 31958
rect 209522 31144 210090 31958
rect 210258 31144 210826 31958
rect 210994 31144 211562 31958
rect 211730 31144 212298 31958
rect 212466 31144 213034 31958
rect 213202 31144 213770 31958
rect 213938 31144 214506 31958
rect 214674 31144 215242 31958
rect 215410 31144 215978 31958
rect 216146 31144 216714 31958
rect 216882 31144 217450 31958
rect 217618 31144 218186 31958
rect 218354 31144 218922 31958
rect 219090 31144 219658 31958
rect 219826 31144 220394 31958
rect 220562 31144 221130 31958
rect 221298 31144 221866 31958
rect 222034 31144 222602 31958
rect 222770 31144 223338 31958
rect 223506 31144 224074 31958
rect 224242 31144 224810 31958
rect 224978 31144 225546 31958
rect 225714 31144 226282 31958
rect 226450 31144 227018 31958
rect 227186 31144 227754 31958
rect 227922 31144 228490 31958
rect 228658 31144 229226 31958
rect 229394 31144 229962 31958
rect 230130 31144 230698 31958
rect 230866 31144 231434 31958
rect 231602 31144 232170 31958
rect 232338 31144 232906 31958
rect 233074 31144 233642 31958
rect 233810 31144 234378 31958
rect 234546 31144 235114 31958
rect 235282 31144 235850 31958
rect 236018 31144 236586 31958
rect 236754 31144 237322 31958
rect 237490 31144 238058 31958
rect 238226 31144 238794 31958
rect 238962 31144 239530 31958
rect 239698 31144 240266 31958
rect 240434 31144 241002 31958
rect 241170 31144 241738 31958
rect 241906 31144 242474 31958
rect 242642 31144 243210 31958
rect 243378 31144 243946 31958
rect 244114 31144 244682 31958
rect 244850 31144 245418 31958
rect 245586 31144 246154 31958
rect 246322 31144 246890 31958
rect 247058 31144 247626 31958
rect 247794 31144 248362 31958
rect 248530 31144 249098 31958
rect 249266 31144 249834 31958
rect 250002 31144 250570 31958
rect 250738 31144 251306 31958
rect 251474 31144 252042 31958
rect 252210 31144 252778 31958
rect 252946 31144 253514 31958
rect 253682 31144 254250 31958
rect 254418 31144 254986 31958
rect 255154 31144 255722 31958
rect 255890 31144 256458 31958
rect 256626 31144 257194 31958
rect 257362 31144 257930 31958
rect 258098 31144 258666 31958
rect 258834 31144 259402 31958
rect 259570 31144 260138 31958
rect 260306 31144 260874 31958
rect 261042 31144 261610 31958
rect 261778 31144 262346 31958
rect 262514 31144 263082 31958
rect 263250 31144 263818 31958
rect 263986 31144 264554 31958
rect 264722 31144 265290 31958
rect 265458 31144 266026 31958
rect 266194 31144 266762 31958
rect 266930 31144 267498 31958
rect 267666 31144 268234 31958
rect 268402 31144 268970 31958
rect 269138 31144 269706 31958
rect 269874 31144 270442 31958
rect 270610 31144 271178 31958
rect 271346 31144 271914 31958
rect 272082 31144 272650 31958
rect 272818 31144 273386 31958
rect 273554 31144 274122 31958
rect 274290 31144 274858 31958
rect 275026 31144 275594 31958
rect 275762 31144 276330 31958
rect 276498 31144 277066 31958
rect 277234 31144 277802 31958
rect 277970 31144 278538 31958
rect 278706 31144 279274 31958
rect 279442 31144 280010 31958
rect 280178 31144 280746 31958
rect 280914 31144 281482 31958
rect 281650 31144 282218 31958
rect 282386 31144 282954 31958
rect 283122 31144 283690 31958
rect 283858 31144 284426 31958
rect 284594 31144 285162 31958
rect 285330 31144 285898 31958
rect 286066 31144 286634 31958
rect 286802 31144 287370 31958
rect 287538 31144 288106 31958
rect 288274 31144 288842 31958
rect 289010 31144 289578 31958
rect 289746 31144 290314 31958
rect 290482 31144 291050 31958
rect 291218 31144 291786 31958
rect 291954 31144 292522 31958
rect 292690 31144 293258 31958
rect 293426 31144 293994 31958
rect 294162 31144 294730 31958
rect 294898 31144 295466 31958
rect 295634 31144 296202 31958
rect 296370 31144 296938 31958
rect 297106 31144 297674 31958
rect 297842 31144 298410 31958
rect 298578 31144 299146 31958
rect 299314 31144 299882 31958
rect 300050 31144 300618 31958
rect 300786 31144 301354 31958
rect 301522 31144 302090 31958
rect 302258 31144 302826 31958
rect 302994 31144 303562 31958
rect 303730 31144 304298 31958
rect 304466 31144 305034 31958
rect 305202 31144 305770 31958
rect 305938 31144 306506 31958
rect 306674 31144 307242 31958
rect 307410 31144 307978 31958
rect 308146 31144 308714 31958
rect 308882 31144 309450 31958
rect 309618 31144 310186 31958
rect 310354 31144 310922 31958
rect 311090 31144 311658 31958
rect 311826 31144 312394 31958
rect 312562 31144 313130 31958
rect 313298 31144 313866 31958
rect 314034 31144 314602 31958
rect 314770 31144 315338 31958
rect 315506 31144 316074 31958
rect 316242 31144 316810 31958
rect 316978 31144 317546 31958
rect 317714 31144 318282 31958
rect 318450 31144 319018 31958
rect 319186 31144 319754 31958
rect 319922 31144 320490 31958
rect 320658 31144 321226 31958
rect 321394 31144 321962 31958
rect 322130 31144 322698 31958
rect 322866 31144 323434 31958
rect 323602 31144 324170 31958
rect 324338 31144 324906 31958
rect 325074 31144 325642 31958
rect 325810 31144 326378 31958
rect 326546 31144 327114 31958
rect 327282 31144 327850 31958
rect 328018 31144 328586 31958
rect 328754 31144 329322 31958
rect 329490 31144 330058 31958
rect 330226 31144 330794 31958
rect 330962 31144 331530 31958
rect 331698 31144 332266 31958
rect 332434 31144 333002 31958
rect 333170 31144 333738 31958
rect 333906 31144 334474 31958
rect 334642 31144 335210 31958
rect 335378 31144 335946 31958
rect 336114 31144 336682 31958
rect 336850 31144 337418 31958
rect 337586 31144 338154 31958
rect 338322 31144 338890 31958
rect 339058 31144 339626 31958
rect 339794 31144 340362 31958
rect 340530 31144 341098 31958
rect 341266 31144 341834 31958
rect 342002 31144 342570 31958
rect 342738 31144 343306 31958
rect 343474 31144 344042 31958
rect 344210 31144 344778 31958
rect 344946 31144 345514 31958
rect 345682 31144 346250 31958
rect 346418 31144 346986 31958
rect 347154 31144 347722 31958
rect 347890 31144 348458 31958
rect 348626 31144 349194 31958
rect 349362 31144 349930 31958
rect 350098 31144 350666 31958
rect 350834 31144 351402 31958
rect 351570 31144 352138 31958
rect 352306 31144 352874 31958
rect 353042 31144 353610 31958
rect 353778 31144 354346 31958
rect 354514 31144 355082 31958
rect 355250 31144 355818 31958
rect 355986 31144 356554 31958
rect 356722 31144 357290 31958
rect 357458 31144 358026 31958
rect 358194 31144 358762 31958
rect 358930 31144 359498 31958
rect 359666 31144 360234 31958
rect 360402 31144 360970 31958
rect 361138 31144 361706 31958
rect 361874 31144 362442 31958
rect 362610 31144 363178 31958
rect 363346 31144 363914 31958
rect 364082 31144 364650 31958
rect 364818 31144 365386 31958
rect 365554 31144 366122 31958
rect 366290 31144 366858 31958
rect 367026 31144 367594 31958
rect 367762 31144 368330 31958
rect 368498 31144 369066 31958
rect 369234 31144 369802 31958
rect 369970 31144 370538 31958
rect 370706 31144 371274 31958
rect 371442 31144 378378 31958
rect 5036 856 378378 31144
rect 5036 2 19834 856
rect 20002 2 20386 856
rect 20554 2 20938 856
rect 21106 2 21490 856
rect 21658 2 22042 856
rect 22210 2 22594 856
rect 22762 2 23146 856
rect 23314 2 23698 856
rect 23866 2 24250 856
rect 24418 2 24802 856
rect 24970 2 25354 856
rect 25522 2 25906 856
rect 26074 2 26458 856
rect 26626 2 27010 856
rect 27178 2 27562 856
rect 27730 2 28114 856
rect 28282 2 28666 856
rect 28834 2 29218 856
rect 29386 2 29770 856
rect 29938 2 30322 856
rect 30490 2 30874 856
rect 31042 2 31426 856
rect 31594 2 31978 856
rect 32146 2 32530 856
rect 32698 2 33082 856
rect 33250 2 33634 856
rect 33802 2 34186 856
rect 34354 2 34738 856
rect 34906 2 35290 856
rect 35458 2 35842 856
rect 36010 2 36394 856
rect 36562 2 36946 856
rect 37114 2 37498 856
rect 37666 2 38050 856
rect 38218 2 38602 856
rect 38770 2 39154 856
rect 39322 2 39706 856
rect 39874 2 40258 856
rect 40426 2 40810 856
rect 40978 2 41362 856
rect 41530 2 41914 856
rect 42082 2 42466 856
rect 42634 2 43018 856
rect 43186 2 43570 856
rect 43738 2 44122 856
rect 44290 2 44674 856
rect 44842 2 45226 856
rect 45394 2 45778 856
rect 45946 2 46330 856
rect 46498 2 46882 856
rect 47050 2 47434 856
rect 47602 2 47986 856
rect 48154 2 48538 856
rect 48706 2 49090 856
rect 49258 2 49642 856
rect 49810 2 50194 856
rect 50362 2 50746 856
rect 50914 2 51298 856
rect 51466 2 51850 856
rect 52018 2 52402 856
rect 52570 2 52954 856
rect 53122 2 53506 856
rect 53674 2 54058 856
rect 54226 2 54610 856
rect 54778 2 55162 856
rect 55330 2 55714 856
rect 55882 2 56266 856
rect 56434 2 56818 856
rect 56986 2 57370 856
rect 57538 2 57922 856
rect 58090 2 58474 856
rect 58642 2 59026 856
rect 59194 2 59578 856
rect 59746 2 60130 856
rect 60298 2 60682 856
rect 60850 2 61234 856
rect 61402 2 61786 856
rect 61954 2 62338 856
rect 62506 2 62890 856
rect 63058 2 63442 856
rect 63610 2 63994 856
rect 64162 2 64546 856
rect 64714 2 65098 856
rect 65266 2 65650 856
rect 65818 2 66202 856
rect 66370 2 66754 856
rect 66922 2 67306 856
rect 67474 2 67858 856
rect 68026 2 68410 856
rect 68578 2 68962 856
rect 69130 2 69514 856
rect 69682 2 70066 856
rect 70234 2 70618 856
rect 70786 2 71170 856
rect 71338 2 71722 856
rect 71890 2 72274 856
rect 72442 2 72826 856
rect 72994 2 73378 856
rect 73546 2 73930 856
rect 74098 2 74482 856
rect 74650 2 75034 856
rect 75202 2 75586 856
rect 75754 2 76138 856
rect 76306 2 76690 856
rect 76858 2 77242 856
rect 77410 2 77794 856
rect 77962 2 78346 856
rect 78514 2 78898 856
rect 79066 2 79450 856
rect 79618 2 80002 856
rect 80170 2 80554 856
rect 80722 2 81106 856
rect 81274 2 81658 856
rect 81826 2 82210 856
rect 82378 2 82762 856
rect 82930 2 83314 856
rect 83482 2 83866 856
rect 84034 2 84418 856
rect 84586 2 84970 856
rect 85138 2 85522 856
rect 85690 2 86074 856
rect 86242 2 86626 856
rect 86794 2 87178 856
rect 87346 2 87730 856
rect 87898 2 88282 856
rect 88450 2 88834 856
rect 89002 2 89386 856
rect 89554 2 89938 856
rect 90106 2 90490 856
rect 90658 2 91042 856
rect 91210 2 91594 856
rect 91762 2 92146 856
rect 92314 2 92698 856
rect 92866 2 93250 856
rect 93418 2 93802 856
rect 93970 2 94354 856
rect 94522 2 94906 856
rect 95074 2 95458 856
rect 95626 2 96010 856
rect 96178 2 96562 856
rect 96730 2 97114 856
rect 97282 2 97666 856
rect 97834 2 98218 856
rect 98386 2 98770 856
rect 98938 2 99322 856
rect 99490 2 99874 856
rect 100042 2 100426 856
rect 100594 2 100978 856
rect 101146 2 101530 856
rect 101698 2 102082 856
rect 102250 2 102634 856
rect 102802 2 103186 856
rect 103354 2 103738 856
rect 103906 2 104290 856
rect 104458 2 104842 856
rect 105010 2 105394 856
rect 105562 2 105946 856
rect 106114 2 106498 856
rect 106666 2 107050 856
rect 107218 2 107602 856
rect 107770 2 108154 856
rect 108322 2 108706 856
rect 108874 2 109258 856
rect 109426 2 109810 856
rect 109978 2 110362 856
rect 110530 2 110914 856
rect 111082 2 111466 856
rect 111634 2 112018 856
rect 112186 2 112570 856
rect 112738 2 113122 856
rect 113290 2 113674 856
rect 113842 2 114226 856
rect 114394 2 114778 856
rect 114946 2 115330 856
rect 115498 2 115882 856
rect 116050 2 116434 856
rect 116602 2 116986 856
rect 117154 2 117538 856
rect 117706 2 118090 856
rect 118258 2 118642 856
rect 118810 2 119194 856
rect 119362 2 119746 856
rect 119914 2 120298 856
rect 120466 2 120850 856
rect 121018 2 121402 856
rect 121570 2 121954 856
rect 122122 2 122506 856
rect 122674 2 123058 856
rect 123226 2 123610 856
rect 123778 2 124162 856
rect 124330 2 124714 856
rect 124882 2 125266 856
rect 125434 2 125818 856
rect 125986 2 126370 856
rect 126538 2 126922 856
rect 127090 2 127474 856
rect 127642 2 128026 856
rect 128194 2 128578 856
rect 128746 2 129130 856
rect 129298 2 129682 856
rect 129850 2 130234 856
rect 130402 2 130786 856
rect 130954 2 131338 856
rect 131506 2 131890 856
rect 132058 2 132442 856
rect 132610 2 132994 856
rect 133162 2 133546 856
rect 133714 2 134098 856
rect 134266 2 134650 856
rect 134818 2 135202 856
rect 135370 2 135754 856
rect 135922 2 136306 856
rect 136474 2 136858 856
rect 137026 2 137410 856
rect 137578 2 137962 856
rect 138130 2 138514 856
rect 138682 2 139066 856
rect 139234 2 139618 856
rect 139786 2 140170 856
rect 140338 2 140722 856
rect 140890 2 141274 856
rect 141442 2 141826 856
rect 141994 2 142378 856
rect 142546 2 142930 856
rect 143098 2 143482 856
rect 143650 2 144034 856
rect 144202 2 144586 856
rect 144754 2 145138 856
rect 145306 2 145690 856
rect 145858 2 146242 856
rect 146410 2 146794 856
rect 146962 2 147346 856
rect 147514 2 147898 856
rect 148066 2 148450 856
rect 148618 2 149002 856
rect 149170 2 149554 856
rect 149722 2 150106 856
rect 150274 2 150658 856
rect 150826 2 151210 856
rect 151378 2 151762 856
rect 151930 2 152314 856
rect 152482 2 152866 856
rect 153034 2 153418 856
rect 153586 2 153970 856
rect 154138 2 154522 856
rect 154690 2 155074 856
rect 155242 2 155626 856
rect 155794 2 156178 856
rect 156346 2 156730 856
rect 156898 2 157282 856
rect 157450 2 157834 856
rect 158002 2 158386 856
rect 158554 2 158938 856
rect 159106 2 159490 856
rect 159658 2 160042 856
rect 160210 2 160594 856
rect 160762 2 161146 856
rect 161314 2 161698 856
rect 161866 2 162250 856
rect 162418 2 162802 856
rect 162970 2 163354 856
rect 163522 2 163906 856
rect 164074 2 164458 856
rect 164626 2 165010 856
rect 165178 2 165562 856
rect 165730 2 166114 856
rect 166282 2 166666 856
rect 166834 2 167218 856
rect 167386 2 167770 856
rect 167938 2 168322 856
rect 168490 2 168874 856
rect 169042 2 169426 856
rect 169594 2 169978 856
rect 170146 2 170530 856
rect 170698 2 171082 856
rect 171250 2 171634 856
rect 171802 2 172186 856
rect 172354 2 172738 856
rect 172906 2 173290 856
rect 173458 2 173842 856
rect 174010 2 174394 856
rect 174562 2 174946 856
rect 175114 2 175498 856
rect 175666 2 176050 856
rect 176218 2 176602 856
rect 176770 2 177154 856
rect 177322 2 177706 856
rect 177874 2 178258 856
rect 178426 2 178810 856
rect 178978 2 179362 856
rect 179530 2 179914 856
rect 180082 2 180466 856
rect 180634 2 181018 856
rect 181186 2 181570 856
rect 181738 2 182122 856
rect 182290 2 182674 856
rect 182842 2 183226 856
rect 183394 2 183778 856
rect 183946 2 184330 856
rect 184498 2 184882 856
rect 185050 2 185434 856
rect 185602 2 185986 856
rect 186154 2 186538 856
rect 186706 2 187090 856
rect 187258 2 187642 856
rect 187810 2 188194 856
rect 188362 2 188746 856
rect 188914 2 189298 856
rect 189466 2 189850 856
rect 190018 2 190402 856
rect 190570 2 190954 856
rect 191122 2 191506 856
rect 191674 2 192058 856
rect 192226 2 192610 856
rect 192778 2 193162 856
rect 193330 2 193714 856
rect 193882 2 194266 856
rect 194434 2 194818 856
rect 194986 2 195370 856
rect 195538 2 195922 856
rect 196090 2 196474 856
rect 196642 2 197026 856
rect 197194 2 197578 856
rect 197746 2 198130 856
rect 198298 2 198682 856
rect 198850 2 199234 856
rect 199402 2 199786 856
rect 199954 2 200338 856
rect 200506 2 200890 856
rect 201058 2 201442 856
rect 201610 2 201994 856
rect 202162 2 202546 856
rect 202714 2 203098 856
rect 203266 2 203650 856
rect 203818 2 204202 856
rect 204370 2 204754 856
rect 204922 2 205306 856
rect 205474 2 205858 856
rect 206026 2 206410 856
rect 206578 2 206962 856
rect 207130 2 207514 856
rect 207682 2 208066 856
rect 208234 2 208618 856
rect 208786 2 209170 856
rect 209338 2 209722 856
rect 209890 2 210274 856
rect 210442 2 210826 856
rect 210994 2 211378 856
rect 211546 2 211930 856
rect 212098 2 212482 856
rect 212650 2 213034 856
rect 213202 2 213586 856
rect 213754 2 214138 856
rect 214306 2 214690 856
rect 214858 2 215242 856
rect 215410 2 215794 856
rect 215962 2 216346 856
rect 216514 2 216898 856
rect 217066 2 217450 856
rect 217618 2 218002 856
rect 218170 2 218554 856
rect 218722 2 219106 856
rect 219274 2 219658 856
rect 219826 2 220210 856
rect 220378 2 220762 856
rect 220930 2 221314 856
rect 221482 2 221866 856
rect 222034 2 222418 856
rect 222586 2 222970 856
rect 223138 2 223522 856
rect 223690 2 224074 856
rect 224242 2 224626 856
rect 224794 2 225178 856
rect 225346 2 225730 856
rect 225898 2 226282 856
rect 226450 2 226834 856
rect 227002 2 227386 856
rect 227554 2 227938 856
rect 228106 2 228490 856
rect 228658 2 229042 856
rect 229210 2 229594 856
rect 229762 2 230146 856
rect 230314 2 230698 856
rect 230866 2 231250 856
rect 231418 2 231802 856
rect 231970 2 232354 856
rect 232522 2 232906 856
rect 233074 2 233458 856
rect 233626 2 234010 856
rect 234178 2 234562 856
rect 234730 2 235114 856
rect 235282 2 235666 856
rect 235834 2 236218 856
rect 236386 2 236770 856
rect 236938 2 237322 856
rect 237490 2 237874 856
rect 238042 2 238426 856
rect 238594 2 238978 856
rect 239146 2 239530 856
rect 239698 2 240082 856
rect 240250 2 240634 856
rect 240802 2 241186 856
rect 241354 2 241738 856
rect 241906 2 242290 856
rect 242458 2 242842 856
rect 243010 2 243394 856
rect 243562 2 243946 856
rect 244114 2 244498 856
rect 244666 2 245050 856
rect 245218 2 245602 856
rect 245770 2 246154 856
rect 246322 2 246706 856
rect 246874 2 247258 856
rect 247426 2 247810 856
rect 247978 2 248362 856
rect 248530 2 248914 856
rect 249082 2 249466 856
rect 249634 2 250018 856
rect 250186 2 250570 856
rect 250738 2 251122 856
rect 251290 2 251674 856
rect 251842 2 252226 856
rect 252394 2 252778 856
rect 252946 2 253330 856
rect 253498 2 253882 856
rect 254050 2 254434 856
rect 254602 2 254986 856
rect 255154 2 255538 856
rect 255706 2 256090 856
rect 256258 2 256642 856
rect 256810 2 257194 856
rect 257362 2 257746 856
rect 257914 2 258298 856
rect 258466 2 258850 856
rect 259018 2 259402 856
rect 259570 2 259954 856
rect 260122 2 260506 856
rect 260674 2 261058 856
rect 261226 2 261610 856
rect 261778 2 262162 856
rect 262330 2 262714 856
rect 262882 2 263266 856
rect 263434 2 263818 856
rect 263986 2 264370 856
rect 264538 2 264922 856
rect 265090 2 265474 856
rect 265642 2 266026 856
rect 266194 2 266578 856
rect 266746 2 267130 856
rect 267298 2 267682 856
rect 267850 2 268234 856
rect 268402 2 268786 856
rect 268954 2 269338 856
rect 269506 2 269890 856
rect 270058 2 270442 856
rect 270610 2 270994 856
rect 271162 2 271546 856
rect 271714 2 272098 856
rect 272266 2 272650 856
rect 272818 2 273202 856
rect 273370 2 273754 856
rect 273922 2 274306 856
rect 274474 2 274858 856
rect 275026 2 275410 856
rect 275578 2 275962 856
rect 276130 2 276514 856
rect 276682 2 277066 856
rect 277234 2 277618 856
rect 277786 2 278170 856
rect 278338 2 278722 856
rect 278890 2 279274 856
rect 279442 2 279826 856
rect 279994 2 280378 856
rect 280546 2 280930 856
rect 281098 2 281482 856
rect 281650 2 282034 856
rect 282202 2 282586 856
rect 282754 2 283138 856
rect 283306 2 283690 856
rect 283858 2 284242 856
rect 284410 2 284794 856
rect 284962 2 285346 856
rect 285514 2 285898 856
rect 286066 2 286450 856
rect 286618 2 287002 856
rect 287170 2 287554 856
rect 287722 2 288106 856
rect 288274 2 288658 856
rect 288826 2 289210 856
rect 289378 2 289762 856
rect 289930 2 290314 856
rect 290482 2 290866 856
rect 291034 2 291418 856
rect 291586 2 291970 856
rect 292138 2 292522 856
rect 292690 2 293074 856
rect 293242 2 293626 856
rect 293794 2 294178 856
rect 294346 2 294730 856
rect 294898 2 295282 856
rect 295450 2 295834 856
rect 296002 2 296386 856
rect 296554 2 296938 856
rect 297106 2 297490 856
rect 297658 2 298042 856
rect 298210 2 298594 856
rect 298762 2 299146 856
rect 299314 2 299698 856
rect 299866 2 300250 856
rect 300418 2 300802 856
rect 300970 2 301354 856
rect 301522 2 301906 856
rect 302074 2 302458 856
rect 302626 2 303010 856
rect 303178 2 303562 856
rect 303730 2 304114 856
rect 304282 2 304666 856
rect 304834 2 305218 856
rect 305386 2 305770 856
rect 305938 2 306322 856
rect 306490 2 306874 856
rect 307042 2 307426 856
rect 307594 2 307978 856
rect 308146 2 308530 856
rect 308698 2 309082 856
rect 309250 2 309634 856
rect 309802 2 310186 856
rect 310354 2 310738 856
rect 310906 2 311290 856
rect 311458 2 311842 856
rect 312010 2 312394 856
rect 312562 2 312946 856
rect 313114 2 313498 856
rect 313666 2 314050 856
rect 314218 2 314602 856
rect 314770 2 315154 856
rect 315322 2 315706 856
rect 315874 2 316258 856
rect 316426 2 316810 856
rect 316978 2 317362 856
rect 317530 2 317914 856
rect 318082 2 318466 856
rect 318634 2 319018 856
rect 319186 2 319570 856
rect 319738 2 320122 856
rect 320290 2 320674 856
rect 320842 2 321226 856
rect 321394 2 321778 856
rect 321946 2 322330 856
rect 322498 2 322882 856
rect 323050 2 323434 856
rect 323602 2 323986 856
rect 324154 2 324538 856
rect 324706 2 325090 856
rect 325258 2 325642 856
rect 325810 2 326194 856
rect 326362 2 326746 856
rect 326914 2 327298 856
rect 327466 2 327850 856
rect 328018 2 328402 856
rect 328570 2 328954 856
rect 329122 2 329506 856
rect 329674 2 330058 856
rect 330226 2 330610 856
rect 330778 2 331162 856
rect 331330 2 331714 856
rect 331882 2 332266 856
rect 332434 2 332818 856
rect 332986 2 333370 856
rect 333538 2 333922 856
rect 334090 2 334474 856
rect 334642 2 335026 856
rect 335194 2 335578 856
rect 335746 2 336130 856
rect 336298 2 336682 856
rect 336850 2 337234 856
rect 337402 2 337786 856
rect 337954 2 338338 856
rect 338506 2 338890 856
rect 339058 2 339442 856
rect 339610 2 339994 856
rect 340162 2 340546 856
rect 340714 2 341098 856
rect 341266 2 341650 856
rect 341818 2 342202 856
rect 342370 2 342754 856
rect 342922 2 343306 856
rect 343474 2 343858 856
rect 344026 2 344410 856
rect 344578 2 344962 856
rect 345130 2 345514 856
rect 345682 2 346066 856
rect 346234 2 346618 856
rect 346786 2 347170 856
rect 347338 2 347722 856
rect 347890 2 348274 856
rect 348442 2 348826 856
rect 348994 2 349378 856
rect 349546 2 349930 856
rect 350098 2 350482 856
rect 350650 2 351034 856
rect 351202 2 351586 856
rect 351754 2 352138 856
rect 352306 2 352690 856
rect 352858 2 353242 856
rect 353410 2 353794 856
rect 353962 2 354346 856
rect 354514 2 354898 856
rect 355066 2 355450 856
rect 355618 2 356002 856
rect 356170 2 356554 856
rect 356722 2 357106 856
rect 357274 2 357658 856
rect 357826 2 358210 856
rect 358378 2 358762 856
rect 358930 2 359314 856
rect 359482 2 359866 856
rect 360034 2 378378 856
<< metal3 >>
rect 379200 30608 380400 30728
rect 379200 28160 380400 28280
rect 379200 25712 380400 25832
rect 379200 23264 380400 23384
rect 379200 20816 380400 20936
rect 379200 18368 380400 18488
rect 379200 15920 380400 16040
rect 379200 13472 380400 13592
rect 379200 11024 380400 11144
rect 379200 8576 380400 8696
rect 379200 6128 380400 6248
rect 379200 3680 380400 3800
rect 379200 1232 380400 1352
<< obsm3 >>
rect 5026 30808 379200 31925
rect 5026 30528 379120 30808
rect 5026 28360 379200 30528
rect 5026 28080 379120 28360
rect 5026 25912 379200 28080
rect 5026 25632 379120 25912
rect 5026 23464 379200 25632
rect 5026 23184 379120 23464
rect 5026 21016 379200 23184
rect 5026 20736 379120 21016
rect 5026 18568 379200 20736
rect 5026 18288 379120 18568
rect 5026 16120 379200 18288
rect 5026 15840 379120 16120
rect 5026 13672 379200 15840
rect 5026 13392 379120 13672
rect 5026 11224 379200 13392
rect 5026 10944 379120 11224
rect 5026 8776 379200 10944
rect 5026 8496 379120 8776
rect 5026 6328 379200 8496
rect 5026 6048 379120 6328
rect 5026 3880 379200 6048
rect 5026 3600 379120 3880
rect 5026 1432 379200 3600
rect 5026 1152 379120 1432
rect 5026 35 379200 1152
<< metal4 >>
rect 5014 1040 5194 30512
rect 12394 1040 12574 30512
rect 20064 1040 20244 30512
rect 27444 1040 27624 30512
rect 35114 1040 35294 30512
rect 42494 1040 42674 30512
rect 50164 1040 50344 30512
rect 57544 1040 57724 30512
rect 65214 1040 65394 30512
rect 66854 1040 67034 30512
rect 71034 1040 71214 30512
rect 72594 1040 72774 30512
rect 76854 1040 77034 30512
rect 80264 1040 80444 30512
rect 81034 1040 81214 30512
rect 87644 1040 87824 30512
rect 95314 1040 95494 30512
rect 102694 1040 102874 30512
rect 110364 1040 110544 30512
rect 117744 1040 117924 30512
rect 125414 1040 125594 30512
rect 132794 1040 132974 30512
rect 140464 1040 140644 30512
rect 141284 1040 141464 30512
rect 147844 1040 148024 30512
rect 148664 1040 148844 30512
rect 155514 1040 155694 30512
rect 156334 1040 156514 30512
rect 162894 1040 163074 30512
rect 163714 1040 163894 30512
rect 170564 1040 170744 30512
rect 171384 1040 171564 30512
rect 177944 1040 178124 30512
rect 178764 1040 178944 30512
rect 185614 1040 185794 30512
rect 186434 1040 186614 30512
rect 192994 1040 193174 30512
rect 193814 1040 193994 30512
rect 200664 1040 200844 30512
rect 208044 1040 208224 30512
rect 215714 1040 215894 30512
rect 223094 1040 223274 30512
rect 230764 1040 230944 30512
rect 238144 1040 238324 30512
rect 245814 1040 245994 30512
rect 253194 1040 253374 30512
rect 255814 1040 255994 30512
rect 256614 1040 256794 30512
rect 260864 1040 261044 30512
rect 263194 1040 263374 30512
rect 263994 1040 264174 30512
rect 268244 1040 268424 30512
rect 270864 1040 271044 30512
rect 271664 1040 271844 30512
rect 275914 1040 276094 30512
rect 278244 1040 278424 30512
rect 279044 1040 279224 30512
rect 283294 1040 283474 30512
rect 290964 1040 291144 30512
rect 298344 1040 298524 30512
rect 306014 1040 306194 30512
rect 313394 1040 313574 30512
rect 321064 1040 321244 30512
rect 328444 1040 328624 30512
rect 336114 1040 336294 30512
rect 343494 1040 343674 30512
rect 351164 1040 351344 30512
rect 358544 1040 358724 30512
rect 366214 1040 366394 30512
rect 373594 1040 373774 30512
<< obsm4 >>
rect 57835 960 65134 29205
rect 65474 960 66774 29205
rect 67114 960 70954 29205
rect 71294 960 72514 29205
rect 72854 960 76774 29205
rect 77114 960 80184 29205
rect 80524 960 80954 29205
rect 81294 960 87564 29205
rect 87904 960 95234 29205
rect 95574 960 102614 29205
rect 102954 960 110284 29205
rect 110624 960 117664 29205
rect 118004 960 125334 29205
rect 125674 960 132714 29205
rect 133054 960 140384 29205
rect 140724 960 141204 29205
rect 141544 960 147764 29205
rect 148104 960 148584 29205
rect 148924 960 155434 29205
rect 155774 960 156254 29205
rect 156594 960 162814 29205
rect 163154 960 163634 29205
rect 163974 960 170484 29205
rect 170824 960 171304 29205
rect 171644 960 177864 29205
rect 178204 960 178684 29205
rect 179024 960 185534 29205
rect 185874 960 186354 29205
rect 186694 960 192914 29205
rect 193254 960 193734 29205
rect 194074 960 200584 29205
rect 200924 960 207964 29205
rect 208304 960 215634 29205
rect 215974 960 223014 29205
rect 223354 960 230684 29205
rect 231024 960 238064 29205
rect 238404 960 245734 29205
rect 246074 960 253114 29205
rect 253454 960 255734 29205
rect 256074 960 256534 29205
rect 256874 960 260784 29205
rect 261124 960 263114 29205
rect 263454 960 263914 29205
rect 264254 960 268164 29205
rect 268504 960 270784 29205
rect 271124 960 271584 29205
rect 271924 960 275834 29205
rect 276174 960 278164 29205
rect 278504 960 278964 29205
rect 279304 960 283214 29205
rect 283554 960 290884 29205
rect 291224 960 298264 29205
rect 298604 960 305934 29205
rect 306274 960 313314 29205
rect 313654 960 320984 29205
rect 321324 960 328364 29205
rect 328704 960 336034 29205
rect 336374 960 338317 29205
rect 57835 35 338317 960
<< labels >>
rlabel metal3 s 379200 1232 380400 1352 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s 379200 3680 380400 3800 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s 379200 6128 380400 6248 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 86498 31200 86554 32400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 307298 31200 307354 32400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 309506 31200 309562 32400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 311714 31200 311770 32400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 313922 31200 313978 32400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 316130 31200 316186 32400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 318338 31200 318394 32400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 320546 31200 320602 32400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 322754 31200 322810 32400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 324962 31200 325018 32400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 327170 31200 327226 32400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 108578 31200 108634 32400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 329378 31200 329434 32400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 331586 31200 331642 32400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 333794 31200 333850 32400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 336002 31200 336058 32400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 338210 31200 338266 32400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 340418 31200 340474 32400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 342626 31200 342682 32400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 344834 31200 344890 32400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 347042 31200 347098 32400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 349250 31200 349306 32400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 110786 31200 110842 32400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 351458 31200 351514 32400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 353666 31200 353722 32400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 355874 31200 355930 32400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 358082 31200 358138 32400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 360290 31200 360346 32400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 362498 31200 362554 32400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 364706 31200 364762 32400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 366914 31200 366970 32400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 112994 31200 113050 32400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 115202 31200 115258 32400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 117410 31200 117466 32400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 119618 31200 119674 32400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 121826 31200 121882 32400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 124034 31200 124090 32400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 126242 31200 126298 32400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 128450 31200 128506 32400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 88706 31200 88762 32400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 130658 31200 130714 32400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 132866 31200 132922 32400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 135074 31200 135130 32400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 137282 31200 137338 32400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 139490 31200 139546 32400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 141698 31200 141754 32400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 143906 31200 143962 32400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 146114 31200 146170 32400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 148322 31200 148378 32400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 150530 31200 150586 32400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 90914 31200 90970 32400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 152738 31200 152794 32400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 154946 31200 155002 32400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 157154 31200 157210 32400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 159362 31200 159418 32400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 161570 31200 161626 32400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 163778 31200 163834 32400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 165986 31200 166042 32400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 168194 31200 168250 32400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 170402 31200 170458 32400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 172610 31200 172666 32400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 93122 31200 93178 32400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 174818 31200 174874 32400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 177026 31200 177082 32400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 179234 31200 179290 32400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 181442 31200 181498 32400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 183650 31200 183706 32400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 185858 31200 185914 32400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 188066 31200 188122 32400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 190274 31200 190330 32400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 192482 31200 192538 32400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 194690 31200 194746 32400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 95330 31200 95386 32400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 196898 31200 196954 32400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 199106 31200 199162 32400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 201314 31200 201370 32400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 203522 31200 203578 32400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 205730 31200 205786 32400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 207938 31200 207994 32400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 210146 31200 210202 32400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 212354 31200 212410 32400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 214562 31200 214618 32400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 216770 31200 216826 32400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 97538 31200 97594 32400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 218978 31200 219034 32400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 221186 31200 221242 32400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 223394 31200 223450 32400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 225602 31200 225658 32400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 227810 31200 227866 32400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 230018 31200 230074 32400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 232226 31200 232282 32400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 234434 31200 234490 32400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 236642 31200 236698 32400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 238850 31200 238906 32400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 99746 31200 99802 32400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 241058 31200 241114 32400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 243266 31200 243322 32400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 245474 31200 245530 32400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 247682 31200 247738 32400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 249890 31200 249946 32400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 252098 31200 252154 32400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 254306 31200 254362 32400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 256514 31200 256570 32400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 258722 31200 258778 32400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 260930 31200 260986 32400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 101954 31200 102010 32400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 263138 31200 263194 32400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 265346 31200 265402 32400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 267554 31200 267610 32400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 269762 31200 269818 32400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 271970 31200 272026 32400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 274178 31200 274234 32400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 276386 31200 276442 32400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 278594 31200 278650 32400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 280802 31200 280858 32400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 283010 31200 283066 32400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 104162 31200 104218 32400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 285218 31200 285274 32400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 287426 31200 287482 32400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 289634 31200 289690 32400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 291842 31200 291898 32400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 294050 31200 294106 32400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 296258 31200 296314 32400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 298466 31200 298522 32400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 300674 31200 300730 32400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 302882 31200 302938 32400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 305090 31200 305146 32400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 106370 31200 106426 32400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 19890 -400 19946 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 240690 -400 240746 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 242898 -400 242954 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 245106 -400 245162 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 247314 -400 247370 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 249522 -400 249578 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 251730 -400 251786 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 253938 -400 253994 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 256146 -400 256202 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 258354 -400 258410 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 260562 -400 260618 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 41970 -400 42026 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 262770 -400 262826 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 264978 -400 265034 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 267186 -400 267242 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 269394 -400 269450 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 271602 -400 271658 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 273810 -400 273866 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 276018 -400 276074 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 278226 -400 278282 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 280434 -400 280490 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 282642 -400 282698 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 44178 -400 44234 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 284850 -400 284906 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 287058 -400 287114 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 289266 -400 289322 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 291474 -400 291530 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 293682 -400 293738 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 295890 -400 295946 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 298098 -400 298154 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 300306 -400 300362 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 46386 -400 46442 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 48594 -400 48650 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 50802 -400 50858 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 53010 -400 53066 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 55218 -400 55274 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 57426 -400 57482 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 59634 -400 59690 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 61842 -400 61898 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 22098 -400 22154 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 64050 -400 64106 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 66258 -400 66314 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 68466 -400 68522 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 70674 -400 70730 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 72882 -400 72938 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 75090 -400 75146 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 77298 -400 77354 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 79506 -400 79562 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 81714 -400 81770 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 83922 -400 83978 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 24306 -400 24362 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 86130 -400 86186 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 88338 -400 88394 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 90546 -400 90602 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 92754 -400 92810 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 94962 -400 95018 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 97170 -400 97226 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 99378 -400 99434 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 101586 -400 101642 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 103794 -400 103850 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 106002 -400 106058 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 26514 -400 26570 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 108210 -400 108266 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 110418 -400 110474 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 112626 -400 112682 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 114834 -400 114890 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 117042 -400 117098 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 119250 -400 119306 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 121458 -400 121514 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 123666 -400 123722 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 125874 -400 125930 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 128082 -400 128138 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 28722 -400 28778 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 130290 -400 130346 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 132498 -400 132554 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 134706 -400 134762 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 136914 -400 136970 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 139122 -400 139178 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 141330 -400 141386 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 143538 -400 143594 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 145746 -400 145802 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 147954 -400 148010 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 150162 -400 150218 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 30930 -400 30986 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 152370 -400 152426 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 154578 -400 154634 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 156786 -400 156842 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 158994 -400 159050 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 161202 -400 161258 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 163410 -400 163466 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 165618 -400 165674 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 167826 -400 167882 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 170034 -400 170090 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 172242 -400 172298 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 33138 -400 33194 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 174450 -400 174506 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 176658 -400 176714 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 178866 -400 178922 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 181074 -400 181130 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 183282 -400 183338 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 185490 -400 185546 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 187698 -400 187754 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 189906 -400 189962 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 192114 -400 192170 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 194322 -400 194378 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 35346 -400 35402 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 196530 -400 196586 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 198738 -400 198794 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 200946 -400 201002 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 203154 -400 203210 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 205362 -400 205418 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 207570 -400 207626 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 209778 -400 209834 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 211986 -400 212042 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 214194 -400 214250 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 216402 -400 216458 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 37554 -400 37610 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 218610 -400 218666 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 220818 -400 220874 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 223026 -400 223082 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 225234 -400 225290 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 227442 -400 227498 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 229650 -400 229706 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 231858 -400 231914 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 234066 -400 234122 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 236274 -400 236330 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 238482 -400 238538 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 39762 -400 39818 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 87234 31200 87290 32400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 308034 31200 308090 32400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 310242 31200 310298 32400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 312450 31200 312506 32400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 314658 31200 314714 32400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 316866 31200 316922 32400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 319074 31200 319130 32400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 321282 31200 321338 32400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 323490 31200 323546 32400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 325698 31200 325754 32400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 327906 31200 327962 32400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 109314 31200 109370 32400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 330114 31200 330170 32400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 332322 31200 332378 32400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 334530 31200 334586 32400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 336738 31200 336794 32400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 338946 31200 339002 32400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 341154 31200 341210 32400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 343362 31200 343418 32400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 345570 31200 345626 32400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 347778 31200 347834 32400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 349986 31200 350042 32400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 111522 31200 111578 32400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 352194 31200 352250 32400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 354402 31200 354458 32400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 356610 31200 356666 32400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 358818 31200 358874 32400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 361026 31200 361082 32400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 363234 31200 363290 32400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 365442 31200 365498 32400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 367650 31200 367706 32400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 113730 31200 113786 32400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 115938 31200 115994 32400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 118146 31200 118202 32400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 120354 31200 120410 32400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 122562 31200 122618 32400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 124770 31200 124826 32400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 126978 31200 127034 32400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 129186 31200 129242 32400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 89442 31200 89498 32400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 131394 31200 131450 32400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 133602 31200 133658 32400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 135810 31200 135866 32400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 138018 31200 138074 32400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 140226 31200 140282 32400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 142434 31200 142490 32400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 144642 31200 144698 32400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 146850 31200 146906 32400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 149058 31200 149114 32400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 151266 31200 151322 32400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 91650 31200 91706 32400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 153474 31200 153530 32400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 155682 31200 155738 32400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 157890 31200 157946 32400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 160098 31200 160154 32400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 162306 31200 162362 32400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 164514 31200 164570 32400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 166722 31200 166778 32400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 168930 31200 168986 32400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 171138 31200 171194 32400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 173346 31200 173402 32400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 93858 31200 93914 32400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 175554 31200 175610 32400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 177762 31200 177818 32400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 179970 31200 180026 32400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 182178 31200 182234 32400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 184386 31200 184442 32400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 186594 31200 186650 32400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 188802 31200 188858 32400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 191010 31200 191066 32400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 193218 31200 193274 32400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 195426 31200 195482 32400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 96066 31200 96122 32400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 197634 31200 197690 32400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 199842 31200 199898 32400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 202050 31200 202106 32400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 204258 31200 204314 32400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 206466 31200 206522 32400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 208674 31200 208730 32400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 210882 31200 210938 32400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 213090 31200 213146 32400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 215298 31200 215354 32400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 217506 31200 217562 32400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 98274 31200 98330 32400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 219714 31200 219770 32400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 221922 31200 221978 32400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 224130 31200 224186 32400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 226338 31200 226394 32400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 228546 31200 228602 32400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 230754 31200 230810 32400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 232962 31200 233018 32400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 235170 31200 235226 32400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 237378 31200 237434 32400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 239586 31200 239642 32400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 100482 31200 100538 32400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 241794 31200 241850 32400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 244002 31200 244058 32400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 246210 31200 246266 32400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 248418 31200 248474 32400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 250626 31200 250682 32400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 252834 31200 252890 32400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 255042 31200 255098 32400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 257250 31200 257306 32400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 259458 31200 259514 32400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 261666 31200 261722 32400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 102690 31200 102746 32400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 263874 31200 263930 32400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 266082 31200 266138 32400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 268290 31200 268346 32400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 270498 31200 270554 32400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 272706 31200 272762 32400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 274914 31200 274970 32400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 277122 31200 277178 32400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 279330 31200 279386 32400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 281538 31200 281594 32400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 283746 31200 283802 32400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 104898 31200 104954 32400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 285954 31200 286010 32400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 288162 31200 288218 32400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 290370 31200 290426 32400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 292578 31200 292634 32400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 294786 31200 294842 32400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 296994 31200 297050 32400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 299202 31200 299258 32400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 301410 31200 301466 32400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 303618 31200 303674 32400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 305826 31200 305882 32400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 107106 31200 107162 32400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 20442 -400 20498 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 241242 -400 241298 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 243450 -400 243506 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 245658 -400 245714 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 247866 -400 247922 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 250074 -400 250130 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 252282 -400 252338 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 254490 -400 254546 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 256698 -400 256754 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 258906 -400 258962 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 261114 -400 261170 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 42522 -400 42578 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 263322 -400 263378 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 265530 -400 265586 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 267738 -400 267794 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 269946 -400 270002 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 272154 -400 272210 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 274362 -400 274418 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 276570 -400 276626 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 278778 -400 278834 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 280986 -400 281042 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 283194 -400 283250 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 44730 -400 44786 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 285402 -400 285458 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 287610 -400 287666 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 289818 -400 289874 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 292026 -400 292082 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 294234 -400 294290 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 296442 -400 296498 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 298650 -400 298706 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 300858 -400 300914 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 46938 -400 46994 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 49146 -400 49202 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 51354 -400 51410 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 53562 -400 53618 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 55770 -400 55826 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 57978 -400 58034 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 60186 -400 60242 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 62394 -400 62450 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 22650 -400 22706 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 64602 -400 64658 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 66810 -400 66866 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 69018 -400 69074 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 71226 -400 71282 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 73434 -400 73490 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 75642 -400 75698 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 77850 -400 77906 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 80058 -400 80114 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 82266 -400 82322 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 84474 -400 84530 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 24858 -400 24914 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 86682 -400 86738 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 88890 -400 88946 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 91098 -400 91154 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 93306 -400 93362 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 95514 -400 95570 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 97722 -400 97778 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 99930 -400 99986 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 102138 -400 102194 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 104346 -400 104402 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 106554 -400 106610 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 27066 -400 27122 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 108762 -400 108818 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 110970 -400 111026 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 113178 -400 113234 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 115386 -400 115442 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 117594 -400 117650 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 119802 -400 119858 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 122010 -400 122066 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 124218 -400 124274 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 126426 -400 126482 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 128634 -400 128690 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 29274 -400 29330 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 130842 -400 130898 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 133050 -400 133106 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 135258 -400 135314 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 137466 -400 137522 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 139674 -400 139730 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 141882 -400 141938 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 144090 -400 144146 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 146298 -400 146354 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 148506 -400 148562 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 150714 -400 150770 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 31482 -400 31538 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 152922 -400 152978 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 155130 -400 155186 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 157338 -400 157394 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 159546 -400 159602 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 161754 -400 161810 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 163962 -400 164018 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 166170 -400 166226 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 168378 -400 168434 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 170586 -400 170642 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 172794 -400 172850 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 33690 -400 33746 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 175002 -400 175058 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 177210 -400 177266 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 179418 -400 179474 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 181626 -400 181682 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 183834 -400 183890 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 186042 -400 186098 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 188250 -400 188306 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 190458 -400 190514 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 192666 -400 192722 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 194874 -400 194930 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 35898 -400 35954 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 197082 -400 197138 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 199290 -400 199346 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 201498 -400 201554 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 203706 -400 203762 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 205914 -400 205970 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 208122 -400 208178 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 210330 -400 210386 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 212538 -400 212594 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 214746 -400 214802 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 216954 -400 217010 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 38106 -400 38162 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 219162 -400 219218 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 221370 -400 221426 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 223578 -400 223634 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 225786 -400 225842 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 227994 -400 228050 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 230202 -400 230258 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 232410 -400 232466 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 234618 -400 234674 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 236826 -400 236882 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 239034 -400 239090 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 40314 -400 40370 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 20994 -400 21050 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 241794 -400 241850 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 244002 -400 244058 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 246210 -400 246266 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 248418 -400 248474 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 250626 -400 250682 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 252834 -400 252890 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 255042 -400 255098 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 257250 -400 257306 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 259458 -400 259514 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 261666 -400 261722 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 43074 -400 43130 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 263874 -400 263930 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 266082 -400 266138 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 268290 -400 268346 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 270498 -400 270554 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 272706 -400 272762 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 274914 -400 274970 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 277122 -400 277178 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 279330 -400 279386 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 281538 -400 281594 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 283746 -400 283802 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 45282 -400 45338 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 285954 -400 286010 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 288162 -400 288218 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 290370 -400 290426 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 292578 -400 292634 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 294786 -400 294842 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 296994 -400 297050 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 299202 -400 299258 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 301410 -400 301466 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 47490 -400 47546 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 49698 -400 49754 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 51906 -400 51962 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 54114 -400 54170 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 56322 -400 56378 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 58530 -400 58586 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 60738 -400 60794 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 62946 -400 63002 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 23202 -400 23258 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 65154 -400 65210 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 67362 -400 67418 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 69570 -400 69626 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 71778 -400 71834 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 73986 -400 74042 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 76194 -400 76250 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 78402 -400 78458 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 80610 -400 80666 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 82818 -400 82874 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 85026 -400 85082 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 25410 -400 25466 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 87234 -400 87290 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 89442 -400 89498 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 91650 -400 91706 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 93858 -400 93914 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 96066 -400 96122 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 100482 -400 100538 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 102690 -400 102746 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 104898 -400 104954 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 107106 -400 107162 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 27618 -400 27674 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 109314 -400 109370 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 111522 -400 111578 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 113730 -400 113786 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 115938 -400 115994 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 118146 -400 118202 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 120354 -400 120410 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 122562 -400 122618 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 124770 -400 124826 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 126978 -400 127034 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 129186 -400 129242 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 29826 -400 29882 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 131394 -400 131450 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 133602 -400 133658 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 135810 -400 135866 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 138018 -400 138074 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 140226 -400 140282 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 142434 -400 142490 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 144642 -400 144698 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 146850 -400 146906 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 149058 -400 149114 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 151266 -400 151322 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 32034 -400 32090 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 153474 -400 153530 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 155682 -400 155738 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 157890 -400 157946 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 160098 -400 160154 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 162306 -400 162362 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 164514 -400 164570 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 166722 -400 166778 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 168930 -400 168986 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 171138 -400 171194 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 173346 -400 173402 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 34242 -400 34298 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 175554 -400 175610 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 177762 -400 177818 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 179970 -400 180026 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 182178 -400 182234 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 184386 -400 184442 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 186594 -400 186650 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 188802 -400 188858 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 191010 -400 191066 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 193218 -400 193274 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 195426 -400 195482 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 36450 -400 36506 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 197634 -400 197690 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 199842 -400 199898 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 202050 -400 202106 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 204258 -400 204314 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 206466 -400 206522 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 208674 -400 208730 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 210882 -400 210938 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 213090 -400 213146 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 215298 -400 215354 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 217506 -400 217562 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 38658 -400 38714 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 219714 -400 219770 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 221922 -400 221978 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 224130 -400 224186 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 226338 -400 226394 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 228546 -400 228602 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 230754 -400 230810 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 232962 -400 233018 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 235170 -400 235226 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 237378 -400 237434 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 239586 -400 239642 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 40866 -400 40922 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 87970 31200 88026 32400 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 308770 31200 308826 32400 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 310978 31200 311034 32400 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 313186 31200 313242 32400 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 315394 31200 315450 32400 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 317602 31200 317658 32400 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 319810 31200 319866 32400 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 322018 31200 322074 32400 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 324226 31200 324282 32400 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 326434 31200 326490 32400 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 328642 31200 328698 32400 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 110050 31200 110106 32400 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 330850 31200 330906 32400 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 333058 31200 333114 32400 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 335266 31200 335322 32400 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 337474 31200 337530 32400 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 339682 31200 339738 32400 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 341890 31200 341946 32400 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 344098 31200 344154 32400 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 346306 31200 346362 32400 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 348514 31200 348570 32400 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 350722 31200 350778 32400 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 112258 31200 112314 32400 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 352930 31200 352986 32400 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 355138 31200 355194 32400 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 357346 31200 357402 32400 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 359554 31200 359610 32400 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 361762 31200 361818 32400 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 363970 31200 364026 32400 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 366178 31200 366234 32400 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 368386 31200 368442 32400 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 114466 31200 114522 32400 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 116674 31200 116730 32400 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 118882 31200 118938 32400 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 121090 31200 121146 32400 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 123298 31200 123354 32400 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 125506 31200 125562 32400 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 127714 31200 127770 32400 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 129922 31200 129978 32400 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 90178 31200 90234 32400 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 132130 31200 132186 32400 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 134338 31200 134394 32400 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 136546 31200 136602 32400 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 138754 31200 138810 32400 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 140962 31200 141018 32400 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 143170 31200 143226 32400 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 145378 31200 145434 32400 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 147586 31200 147642 32400 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 149794 31200 149850 32400 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 152002 31200 152058 32400 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 92386 31200 92442 32400 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 154210 31200 154266 32400 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 156418 31200 156474 32400 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 158626 31200 158682 32400 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 160834 31200 160890 32400 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 163042 31200 163098 32400 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 165250 31200 165306 32400 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 167458 31200 167514 32400 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 169666 31200 169722 32400 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 171874 31200 171930 32400 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 174082 31200 174138 32400 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 94594 31200 94650 32400 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 176290 31200 176346 32400 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 178498 31200 178554 32400 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 180706 31200 180762 32400 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 182914 31200 182970 32400 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 185122 31200 185178 32400 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 187330 31200 187386 32400 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 189538 31200 189594 32400 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 191746 31200 191802 32400 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 193954 31200 194010 32400 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 196162 31200 196218 32400 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 96802 31200 96858 32400 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 198370 31200 198426 32400 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 200578 31200 200634 32400 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 202786 31200 202842 32400 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 204994 31200 205050 32400 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 207202 31200 207258 32400 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 209410 31200 209466 32400 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 211618 31200 211674 32400 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 213826 31200 213882 32400 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 216034 31200 216090 32400 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 218242 31200 218298 32400 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 99010 31200 99066 32400 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 220450 31200 220506 32400 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 222658 31200 222714 32400 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 224866 31200 224922 32400 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 227074 31200 227130 32400 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 229282 31200 229338 32400 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 231490 31200 231546 32400 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 233698 31200 233754 32400 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 235906 31200 235962 32400 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 238114 31200 238170 32400 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 240322 31200 240378 32400 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 101218 31200 101274 32400 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 242530 31200 242586 32400 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 244738 31200 244794 32400 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 246946 31200 247002 32400 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 249154 31200 249210 32400 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 251362 31200 251418 32400 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 253570 31200 253626 32400 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 255778 31200 255834 32400 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 257986 31200 258042 32400 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 260194 31200 260250 32400 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 262402 31200 262458 32400 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 103426 31200 103482 32400 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 264610 31200 264666 32400 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 266818 31200 266874 32400 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 269026 31200 269082 32400 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 271234 31200 271290 32400 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 273442 31200 273498 32400 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 275650 31200 275706 32400 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 277858 31200 277914 32400 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 280066 31200 280122 32400 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 282274 31200 282330 32400 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 284482 31200 284538 32400 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 105634 31200 105690 32400 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 286690 31200 286746 32400 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 288898 31200 288954 32400 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 291106 31200 291162 32400 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 293314 31200 293370 32400 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 295522 31200 295578 32400 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 297730 31200 297786 32400 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 299938 31200 299994 32400 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 302146 31200 302202 32400 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 304354 31200 304410 32400 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 306562 31200 306618 32400 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 107842 31200 107898 32400 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 21546 -400 21602 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 242346 -400 242402 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 244554 -400 244610 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 246762 -400 246818 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 248970 -400 249026 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 251178 -400 251234 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 253386 -400 253442 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 255594 -400 255650 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 257802 -400 257858 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 260010 -400 260066 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 262218 -400 262274 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 43626 -400 43682 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 264426 -400 264482 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 266634 -400 266690 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 268842 -400 268898 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 271050 -400 271106 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 273258 -400 273314 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 275466 -400 275522 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 277674 -400 277730 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 279882 -400 279938 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 282090 -400 282146 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 284298 -400 284354 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 45834 -400 45890 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 286506 -400 286562 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 288714 -400 288770 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 290922 -400 290978 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 293130 -400 293186 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 295338 -400 295394 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 297546 -400 297602 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 299754 -400 299810 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 301962 -400 302018 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 48042 -400 48098 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 50250 -400 50306 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 52458 -400 52514 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 54666 -400 54722 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 56874 -400 56930 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 59082 -400 59138 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 61290 -400 61346 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 63498 -400 63554 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 23754 -400 23810 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 65706 -400 65762 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 67914 -400 67970 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 70122 -400 70178 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 72330 -400 72386 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 74538 -400 74594 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 76746 -400 76802 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 78954 -400 79010 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 81162 -400 81218 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 83370 -400 83426 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 85578 -400 85634 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 25962 -400 26018 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 87786 -400 87842 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 89994 -400 90050 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 92202 -400 92258 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 94410 -400 94466 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 96618 -400 96674 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 98826 -400 98882 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 101034 -400 101090 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 103242 -400 103298 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 105450 -400 105506 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 107658 -400 107714 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 28170 -400 28226 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 109866 -400 109922 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 112074 -400 112130 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 114282 -400 114338 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 116490 -400 116546 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 118698 -400 118754 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 120906 -400 120962 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 123114 -400 123170 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 125322 -400 125378 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 127530 -400 127586 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 129738 -400 129794 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 30378 -400 30434 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 131946 -400 132002 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 134154 -400 134210 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 136362 -400 136418 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 138570 -400 138626 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 140778 -400 140834 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 142986 -400 143042 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 145194 -400 145250 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 147402 -400 147458 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 149610 -400 149666 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 151818 -400 151874 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 32586 -400 32642 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 154026 -400 154082 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 156234 -400 156290 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 158442 -400 158498 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 160650 -400 160706 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 162858 -400 162914 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 165066 -400 165122 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 167274 -400 167330 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 169482 -400 169538 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 171690 -400 171746 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 173898 -400 173954 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 34794 -400 34850 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 176106 -400 176162 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 178314 -400 178370 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 180522 -400 180578 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 182730 -400 182786 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 184938 -400 184994 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 187146 -400 187202 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 189354 -400 189410 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 191562 -400 191618 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 193770 -400 193826 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 195978 -400 196034 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 37002 -400 37058 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 198186 -400 198242 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 200394 -400 200450 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 202602 -400 202658 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 204810 -400 204866 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 207018 -400 207074 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 209226 -400 209282 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 211434 -400 211490 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 213642 -400 213698 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 215850 -400 215906 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 218058 -400 218114 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 39210 -400 39266 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 220266 -400 220322 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 222474 -400 222530 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 224682 -400 224738 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 226890 -400 226946 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 229098 -400 229154 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 231306 -400 231362 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 233514 -400 233570 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 235722 -400 235778 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 237930 -400 237986 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 240138 -400 240194 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 41418 -400 41474 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal2 s 302514 -400 302570 800 6 mprj_ack_i_core
port 900 nsew signal output
rlabel metal2 s 9954 31200 10010 32400 6 mprj_ack_i_user
port 901 nsew signal input
rlabel metal2 s 304722 -400 304778 800 6 mprj_adr_o_core[0]
port 902 nsew signal input
rlabel metal2 s 323490 -400 323546 800 6 mprj_adr_o_core[10]
port 903 nsew signal input
rlabel metal2 s 325146 -400 325202 800 6 mprj_adr_o_core[11]
port 904 nsew signal input
rlabel metal2 s 326802 -400 326858 800 6 mprj_adr_o_core[12]
port 905 nsew signal input
rlabel metal2 s 328458 -400 328514 800 6 mprj_adr_o_core[13]
port 906 nsew signal input
rlabel metal2 s 330114 -400 330170 800 6 mprj_adr_o_core[14]
port 907 nsew signal input
rlabel metal2 s 331770 -400 331826 800 6 mprj_adr_o_core[15]
port 908 nsew signal input
rlabel metal2 s 333426 -400 333482 800 6 mprj_adr_o_core[16]
port 909 nsew signal input
rlabel metal2 s 335082 -400 335138 800 6 mprj_adr_o_core[17]
port 910 nsew signal input
rlabel metal2 s 336738 -400 336794 800 6 mprj_adr_o_core[18]
port 911 nsew signal input
rlabel metal2 s 338394 -400 338450 800 6 mprj_adr_o_core[19]
port 912 nsew signal input
rlabel metal2 s 306930 -400 306986 800 6 mprj_adr_o_core[1]
port 913 nsew signal input
rlabel metal2 s 340050 -400 340106 800 6 mprj_adr_o_core[20]
port 914 nsew signal input
rlabel metal2 s 341706 -400 341762 800 6 mprj_adr_o_core[21]
port 915 nsew signal input
rlabel metal2 s 343362 -400 343418 800 6 mprj_adr_o_core[22]
port 916 nsew signal input
rlabel metal2 s 345018 -400 345074 800 6 mprj_adr_o_core[23]
port 917 nsew signal input
rlabel metal2 s 346674 -400 346730 800 6 mprj_adr_o_core[24]
port 918 nsew signal input
rlabel metal2 s 348330 -400 348386 800 6 mprj_adr_o_core[25]
port 919 nsew signal input
rlabel metal2 s 349986 -400 350042 800 6 mprj_adr_o_core[26]
port 920 nsew signal input
rlabel metal2 s 351642 -400 351698 800 6 mprj_adr_o_core[27]
port 921 nsew signal input
rlabel metal2 s 353298 -400 353354 800 6 mprj_adr_o_core[28]
port 922 nsew signal input
rlabel metal2 s 354954 -400 355010 800 6 mprj_adr_o_core[29]
port 923 nsew signal input
rlabel metal2 s 309138 -400 309194 800 6 mprj_adr_o_core[2]
port 924 nsew signal input
rlabel metal2 s 356610 -400 356666 800 6 mprj_adr_o_core[30]
port 925 nsew signal input
rlabel metal2 s 358266 -400 358322 800 6 mprj_adr_o_core[31]
port 926 nsew signal input
rlabel metal2 s 311346 -400 311402 800 6 mprj_adr_o_core[3]
port 927 nsew signal input
rlabel metal2 s 313554 -400 313610 800 6 mprj_adr_o_core[4]
port 928 nsew signal input
rlabel metal2 s 315210 -400 315266 800 6 mprj_adr_o_core[5]
port 929 nsew signal input
rlabel metal2 s 316866 -400 316922 800 6 mprj_adr_o_core[6]
port 930 nsew signal input
rlabel metal2 s 318522 -400 318578 800 6 mprj_adr_o_core[7]
port 931 nsew signal input
rlabel metal2 s 320178 -400 320234 800 6 mprj_adr_o_core[8]
port 932 nsew signal input
rlabel metal2 s 321834 -400 321890 800 6 mprj_adr_o_core[9]
port 933 nsew signal input
rlabel metal2 s 12898 31200 12954 32400 6 mprj_adr_o_user[0]
port 934 nsew signal output
rlabel metal2 s 37922 31200 37978 32400 6 mprj_adr_o_user[10]
port 935 nsew signal output
rlabel metal2 s 40130 31200 40186 32400 6 mprj_adr_o_user[11]
port 936 nsew signal output
rlabel metal2 s 42338 31200 42394 32400 6 mprj_adr_o_user[12]
port 937 nsew signal output
rlabel metal2 s 44546 31200 44602 32400 6 mprj_adr_o_user[13]
port 938 nsew signal output
rlabel metal2 s 46754 31200 46810 32400 6 mprj_adr_o_user[14]
port 939 nsew signal output
rlabel metal2 s 48962 31200 49018 32400 6 mprj_adr_o_user[15]
port 940 nsew signal output
rlabel metal2 s 51170 31200 51226 32400 6 mprj_adr_o_user[16]
port 941 nsew signal output
rlabel metal2 s 53378 31200 53434 32400 6 mprj_adr_o_user[17]
port 942 nsew signal output
rlabel metal2 s 55586 31200 55642 32400 6 mprj_adr_o_user[18]
port 943 nsew signal output
rlabel metal2 s 57794 31200 57850 32400 6 mprj_adr_o_user[19]
port 944 nsew signal output
rlabel metal2 s 15842 31200 15898 32400 6 mprj_adr_o_user[1]
port 945 nsew signal output
rlabel metal2 s 60002 31200 60058 32400 6 mprj_adr_o_user[20]
port 946 nsew signal output
rlabel metal2 s 62210 31200 62266 32400 6 mprj_adr_o_user[21]
port 947 nsew signal output
rlabel metal2 s 64418 31200 64474 32400 6 mprj_adr_o_user[22]
port 948 nsew signal output
rlabel metal2 s 66626 31200 66682 32400 6 mprj_adr_o_user[23]
port 949 nsew signal output
rlabel metal2 s 68834 31200 68890 32400 6 mprj_adr_o_user[24]
port 950 nsew signal output
rlabel metal2 s 71042 31200 71098 32400 6 mprj_adr_o_user[25]
port 951 nsew signal output
rlabel metal2 s 73250 31200 73306 32400 6 mprj_adr_o_user[26]
port 952 nsew signal output
rlabel metal2 s 75458 31200 75514 32400 6 mprj_adr_o_user[27]
port 953 nsew signal output
rlabel metal2 s 77666 31200 77722 32400 6 mprj_adr_o_user[28]
port 954 nsew signal output
rlabel metal2 s 79874 31200 79930 32400 6 mprj_adr_o_user[29]
port 955 nsew signal output
rlabel metal2 s 18786 31200 18842 32400 6 mprj_adr_o_user[2]
port 956 nsew signal output
rlabel metal2 s 82082 31200 82138 32400 6 mprj_adr_o_user[30]
port 957 nsew signal output
rlabel metal2 s 84290 31200 84346 32400 6 mprj_adr_o_user[31]
port 958 nsew signal output
rlabel metal2 s 21730 31200 21786 32400 6 mprj_adr_o_user[3]
port 959 nsew signal output
rlabel metal2 s 24674 31200 24730 32400 6 mprj_adr_o_user[4]
port 960 nsew signal output
rlabel metal2 s 26882 31200 26938 32400 6 mprj_adr_o_user[5]
port 961 nsew signal output
rlabel metal2 s 29090 31200 29146 32400 6 mprj_adr_o_user[6]
port 962 nsew signal output
rlabel metal2 s 31298 31200 31354 32400 6 mprj_adr_o_user[7]
port 963 nsew signal output
rlabel metal2 s 33506 31200 33562 32400 6 mprj_adr_o_user[8]
port 964 nsew signal output
rlabel metal2 s 35714 31200 35770 32400 6 mprj_adr_o_user[9]
port 965 nsew signal output
rlabel metal2 s 303066 -400 303122 800 6 mprj_cyc_o_core
port 966 nsew signal input
rlabel metal2 s 10690 31200 10746 32400 6 mprj_cyc_o_user
port 967 nsew signal output
rlabel metal2 s 305274 -400 305330 800 6 mprj_dat_i_core[0]
port 968 nsew signal output
rlabel metal2 s 324042 -400 324098 800 6 mprj_dat_i_core[10]
port 969 nsew signal output
rlabel metal2 s 325698 -400 325754 800 6 mprj_dat_i_core[11]
port 970 nsew signal output
rlabel metal2 s 327354 -400 327410 800 6 mprj_dat_i_core[12]
port 971 nsew signal output
rlabel metal2 s 329010 -400 329066 800 6 mprj_dat_i_core[13]
port 972 nsew signal output
rlabel metal2 s 330666 -400 330722 800 6 mprj_dat_i_core[14]
port 973 nsew signal output
rlabel metal2 s 332322 -400 332378 800 6 mprj_dat_i_core[15]
port 974 nsew signal output
rlabel metal2 s 333978 -400 334034 800 6 mprj_dat_i_core[16]
port 975 nsew signal output
rlabel metal2 s 335634 -400 335690 800 6 mprj_dat_i_core[17]
port 976 nsew signal output
rlabel metal2 s 337290 -400 337346 800 6 mprj_dat_i_core[18]
port 977 nsew signal output
rlabel metal2 s 338946 -400 339002 800 6 mprj_dat_i_core[19]
port 978 nsew signal output
rlabel metal2 s 307482 -400 307538 800 6 mprj_dat_i_core[1]
port 979 nsew signal output
rlabel metal2 s 340602 -400 340658 800 6 mprj_dat_i_core[20]
port 980 nsew signal output
rlabel metal2 s 342258 -400 342314 800 6 mprj_dat_i_core[21]
port 981 nsew signal output
rlabel metal2 s 343914 -400 343970 800 6 mprj_dat_i_core[22]
port 982 nsew signal output
rlabel metal2 s 345570 -400 345626 800 6 mprj_dat_i_core[23]
port 983 nsew signal output
rlabel metal2 s 347226 -400 347282 800 6 mprj_dat_i_core[24]
port 984 nsew signal output
rlabel metal2 s 348882 -400 348938 800 6 mprj_dat_i_core[25]
port 985 nsew signal output
rlabel metal2 s 350538 -400 350594 800 6 mprj_dat_i_core[26]
port 986 nsew signal output
rlabel metal2 s 352194 -400 352250 800 6 mprj_dat_i_core[27]
port 987 nsew signal output
rlabel metal2 s 353850 -400 353906 800 6 mprj_dat_i_core[28]
port 988 nsew signal output
rlabel metal2 s 355506 -400 355562 800 6 mprj_dat_i_core[29]
port 989 nsew signal output
rlabel metal2 s 309690 -400 309746 800 6 mprj_dat_i_core[2]
port 990 nsew signal output
rlabel metal2 s 357162 -400 357218 800 6 mprj_dat_i_core[30]
port 991 nsew signal output
rlabel metal2 s 358818 -400 358874 800 6 mprj_dat_i_core[31]
port 992 nsew signal output
rlabel metal2 s 311898 -400 311954 800 6 mprj_dat_i_core[3]
port 993 nsew signal output
rlabel metal2 s 314106 -400 314162 800 6 mprj_dat_i_core[4]
port 994 nsew signal output
rlabel metal2 s 315762 -400 315818 800 6 mprj_dat_i_core[5]
port 995 nsew signal output
rlabel metal2 s 317418 -400 317474 800 6 mprj_dat_i_core[6]
port 996 nsew signal output
rlabel metal2 s 319074 -400 319130 800 6 mprj_dat_i_core[7]
port 997 nsew signal output
rlabel metal2 s 320730 -400 320786 800 6 mprj_dat_i_core[8]
port 998 nsew signal output
rlabel metal2 s 322386 -400 322442 800 6 mprj_dat_i_core[9]
port 999 nsew signal output
rlabel metal2 s 13634 31200 13690 32400 6 mprj_dat_i_user[0]
port 1000 nsew signal input
rlabel metal2 s 38658 31200 38714 32400 6 mprj_dat_i_user[10]
port 1001 nsew signal input
rlabel metal2 s 40866 31200 40922 32400 6 mprj_dat_i_user[11]
port 1002 nsew signal input
rlabel metal2 s 43074 31200 43130 32400 6 mprj_dat_i_user[12]
port 1003 nsew signal input
rlabel metal2 s 45282 31200 45338 32400 6 mprj_dat_i_user[13]
port 1004 nsew signal input
rlabel metal2 s 47490 31200 47546 32400 6 mprj_dat_i_user[14]
port 1005 nsew signal input
rlabel metal2 s 49698 31200 49754 32400 6 mprj_dat_i_user[15]
port 1006 nsew signal input
rlabel metal2 s 51906 31200 51962 32400 6 mprj_dat_i_user[16]
port 1007 nsew signal input
rlabel metal2 s 54114 31200 54170 32400 6 mprj_dat_i_user[17]
port 1008 nsew signal input
rlabel metal2 s 56322 31200 56378 32400 6 mprj_dat_i_user[18]
port 1009 nsew signal input
rlabel metal2 s 58530 31200 58586 32400 6 mprj_dat_i_user[19]
port 1010 nsew signal input
rlabel metal2 s 16578 31200 16634 32400 6 mprj_dat_i_user[1]
port 1011 nsew signal input
rlabel metal2 s 60738 31200 60794 32400 6 mprj_dat_i_user[20]
port 1012 nsew signal input
rlabel metal2 s 62946 31200 63002 32400 6 mprj_dat_i_user[21]
port 1013 nsew signal input
rlabel metal2 s 65154 31200 65210 32400 6 mprj_dat_i_user[22]
port 1014 nsew signal input
rlabel metal2 s 67362 31200 67418 32400 6 mprj_dat_i_user[23]
port 1015 nsew signal input
rlabel metal2 s 69570 31200 69626 32400 6 mprj_dat_i_user[24]
port 1016 nsew signal input
rlabel metal2 s 71778 31200 71834 32400 6 mprj_dat_i_user[25]
port 1017 nsew signal input
rlabel metal2 s 73986 31200 74042 32400 6 mprj_dat_i_user[26]
port 1018 nsew signal input
rlabel metal2 s 76194 31200 76250 32400 6 mprj_dat_i_user[27]
port 1019 nsew signal input
rlabel metal2 s 78402 31200 78458 32400 6 mprj_dat_i_user[28]
port 1020 nsew signal input
rlabel metal2 s 80610 31200 80666 32400 6 mprj_dat_i_user[29]
port 1021 nsew signal input
rlabel metal2 s 19522 31200 19578 32400 6 mprj_dat_i_user[2]
port 1022 nsew signal input
rlabel metal2 s 82818 31200 82874 32400 6 mprj_dat_i_user[30]
port 1023 nsew signal input
rlabel metal2 s 85026 31200 85082 32400 6 mprj_dat_i_user[31]
port 1024 nsew signal input
rlabel metal2 s 22466 31200 22522 32400 6 mprj_dat_i_user[3]
port 1025 nsew signal input
rlabel metal2 s 25410 31200 25466 32400 6 mprj_dat_i_user[4]
port 1026 nsew signal input
rlabel metal2 s 27618 31200 27674 32400 6 mprj_dat_i_user[5]
port 1027 nsew signal input
rlabel metal2 s 29826 31200 29882 32400 6 mprj_dat_i_user[6]
port 1028 nsew signal input
rlabel metal2 s 32034 31200 32090 32400 6 mprj_dat_i_user[7]
port 1029 nsew signal input
rlabel metal2 s 34242 31200 34298 32400 6 mprj_dat_i_user[8]
port 1030 nsew signal input
rlabel metal2 s 36450 31200 36506 32400 6 mprj_dat_i_user[9]
port 1031 nsew signal input
rlabel metal2 s 305826 -400 305882 800 6 mprj_dat_o_core[0]
port 1032 nsew signal input
rlabel metal2 s 324594 -400 324650 800 6 mprj_dat_o_core[10]
port 1033 nsew signal input
rlabel metal2 s 326250 -400 326306 800 6 mprj_dat_o_core[11]
port 1034 nsew signal input
rlabel metal2 s 327906 -400 327962 800 6 mprj_dat_o_core[12]
port 1035 nsew signal input
rlabel metal2 s 329562 -400 329618 800 6 mprj_dat_o_core[13]
port 1036 nsew signal input
rlabel metal2 s 331218 -400 331274 800 6 mprj_dat_o_core[14]
port 1037 nsew signal input
rlabel metal2 s 332874 -400 332930 800 6 mprj_dat_o_core[15]
port 1038 nsew signal input
rlabel metal2 s 334530 -400 334586 800 6 mprj_dat_o_core[16]
port 1039 nsew signal input
rlabel metal2 s 336186 -400 336242 800 6 mprj_dat_o_core[17]
port 1040 nsew signal input
rlabel metal2 s 337842 -400 337898 800 6 mprj_dat_o_core[18]
port 1041 nsew signal input
rlabel metal2 s 339498 -400 339554 800 6 mprj_dat_o_core[19]
port 1042 nsew signal input
rlabel metal2 s 308034 -400 308090 800 6 mprj_dat_o_core[1]
port 1043 nsew signal input
rlabel metal2 s 341154 -400 341210 800 6 mprj_dat_o_core[20]
port 1044 nsew signal input
rlabel metal2 s 342810 -400 342866 800 6 mprj_dat_o_core[21]
port 1045 nsew signal input
rlabel metal2 s 344466 -400 344522 800 6 mprj_dat_o_core[22]
port 1046 nsew signal input
rlabel metal2 s 346122 -400 346178 800 6 mprj_dat_o_core[23]
port 1047 nsew signal input
rlabel metal2 s 347778 -400 347834 800 6 mprj_dat_o_core[24]
port 1048 nsew signal input
rlabel metal2 s 349434 -400 349490 800 6 mprj_dat_o_core[25]
port 1049 nsew signal input
rlabel metal2 s 351090 -400 351146 800 6 mprj_dat_o_core[26]
port 1050 nsew signal input
rlabel metal2 s 352746 -400 352802 800 6 mprj_dat_o_core[27]
port 1051 nsew signal input
rlabel metal2 s 354402 -400 354458 800 6 mprj_dat_o_core[28]
port 1052 nsew signal input
rlabel metal2 s 356058 -400 356114 800 6 mprj_dat_o_core[29]
port 1053 nsew signal input
rlabel metal2 s 310242 -400 310298 800 6 mprj_dat_o_core[2]
port 1054 nsew signal input
rlabel metal2 s 357714 -400 357770 800 6 mprj_dat_o_core[30]
port 1055 nsew signal input
rlabel metal2 s 359370 -400 359426 800 6 mprj_dat_o_core[31]
port 1056 nsew signal input
rlabel metal2 s 312450 -400 312506 800 6 mprj_dat_o_core[3]
port 1057 nsew signal input
rlabel metal2 s 314658 -400 314714 800 6 mprj_dat_o_core[4]
port 1058 nsew signal input
rlabel metal2 s 316314 -400 316370 800 6 mprj_dat_o_core[5]
port 1059 nsew signal input
rlabel metal2 s 317970 -400 318026 800 6 mprj_dat_o_core[6]
port 1060 nsew signal input
rlabel metal2 s 319626 -400 319682 800 6 mprj_dat_o_core[7]
port 1061 nsew signal input
rlabel metal2 s 321282 -400 321338 800 6 mprj_dat_o_core[8]
port 1062 nsew signal input
rlabel metal2 s 322938 -400 322994 800 6 mprj_dat_o_core[9]
port 1063 nsew signal input
rlabel metal2 s 14370 31200 14426 32400 6 mprj_dat_o_user[0]
port 1064 nsew signal output
rlabel metal2 s 39394 31200 39450 32400 6 mprj_dat_o_user[10]
port 1065 nsew signal output
rlabel metal2 s 41602 31200 41658 32400 6 mprj_dat_o_user[11]
port 1066 nsew signal output
rlabel metal2 s 43810 31200 43866 32400 6 mprj_dat_o_user[12]
port 1067 nsew signal output
rlabel metal2 s 46018 31200 46074 32400 6 mprj_dat_o_user[13]
port 1068 nsew signal output
rlabel metal2 s 48226 31200 48282 32400 6 mprj_dat_o_user[14]
port 1069 nsew signal output
rlabel metal2 s 50434 31200 50490 32400 6 mprj_dat_o_user[15]
port 1070 nsew signal output
rlabel metal2 s 52642 31200 52698 32400 6 mprj_dat_o_user[16]
port 1071 nsew signal output
rlabel metal2 s 54850 31200 54906 32400 6 mprj_dat_o_user[17]
port 1072 nsew signal output
rlabel metal2 s 57058 31200 57114 32400 6 mprj_dat_o_user[18]
port 1073 nsew signal output
rlabel metal2 s 59266 31200 59322 32400 6 mprj_dat_o_user[19]
port 1074 nsew signal output
rlabel metal2 s 17314 31200 17370 32400 6 mprj_dat_o_user[1]
port 1075 nsew signal output
rlabel metal2 s 61474 31200 61530 32400 6 mprj_dat_o_user[20]
port 1076 nsew signal output
rlabel metal2 s 63682 31200 63738 32400 6 mprj_dat_o_user[21]
port 1077 nsew signal output
rlabel metal2 s 65890 31200 65946 32400 6 mprj_dat_o_user[22]
port 1078 nsew signal output
rlabel metal2 s 68098 31200 68154 32400 6 mprj_dat_o_user[23]
port 1079 nsew signal output
rlabel metal2 s 70306 31200 70362 32400 6 mprj_dat_o_user[24]
port 1080 nsew signal output
rlabel metal2 s 72514 31200 72570 32400 6 mprj_dat_o_user[25]
port 1081 nsew signal output
rlabel metal2 s 74722 31200 74778 32400 6 mprj_dat_o_user[26]
port 1082 nsew signal output
rlabel metal2 s 76930 31200 76986 32400 6 mprj_dat_o_user[27]
port 1083 nsew signal output
rlabel metal2 s 79138 31200 79194 32400 6 mprj_dat_o_user[28]
port 1084 nsew signal output
rlabel metal2 s 81346 31200 81402 32400 6 mprj_dat_o_user[29]
port 1085 nsew signal output
rlabel metal2 s 20258 31200 20314 32400 6 mprj_dat_o_user[2]
port 1086 nsew signal output
rlabel metal2 s 83554 31200 83610 32400 6 mprj_dat_o_user[30]
port 1087 nsew signal output
rlabel metal2 s 85762 31200 85818 32400 6 mprj_dat_o_user[31]
port 1088 nsew signal output
rlabel metal2 s 23202 31200 23258 32400 6 mprj_dat_o_user[3]
port 1089 nsew signal output
rlabel metal2 s 26146 31200 26202 32400 6 mprj_dat_o_user[4]
port 1090 nsew signal output
rlabel metal2 s 28354 31200 28410 32400 6 mprj_dat_o_user[5]
port 1091 nsew signal output
rlabel metal2 s 30562 31200 30618 32400 6 mprj_dat_o_user[6]
port 1092 nsew signal output
rlabel metal2 s 32770 31200 32826 32400 6 mprj_dat_o_user[7]
port 1093 nsew signal output
rlabel metal2 s 34978 31200 35034 32400 6 mprj_dat_o_user[8]
port 1094 nsew signal output
rlabel metal2 s 37186 31200 37242 32400 6 mprj_dat_o_user[9]
port 1095 nsew signal output
rlabel metal2 s 359922 -400 359978 800 6 mprj_iena_wb
port 1096 nsew signal input
rlabel metal2 s 306378 -400 306434 800 6 mprj_sel_o_core[0]
port 1097 nsew signal input
rlabel metal2 s 308586 -400 308642 800 6 mprj_sel_o_core[1]
port 1098 nsew signal input
rlabel metal2 s 310794 -400 310850 800 6 mprj_sel_o_core[2]
port 1099 nsew signal input
rlabel metal2 s 313002 -400 313058 800 6 mprj_sel_o_core[3]
port 1100 nsew signal input
rlabel metal2 s 15106 31200 15162 32400 6 mprj_sel_o_user[0]
port 1101 nsew signal output
rlabel metal2 s 18050 31200 18106 32400 6 mprj_sel_o_user[1]
port 1102 nsew signal output
rlabel metal2 s 20994 31200 21050 32400 6 mprj_sel_o_user[2]
port 1103 nsew signal output
rlabel metal2 s 23938 31200 23994 32400 6 mprj_sel_o_user[3]
port 1104 nsew signal output
rlabel metal2 s 303618 -400 303674 800 6 mprj_stb_o_core
port 1105 nsew signal input
rlabel metal2 s 11426 31200 11482 32400 6 mprj_stb_o_user
port 1106 nsew signal output
rlabel metal2 s 304170 -400 304226 800 6 mprj_we_o_core
port 1107 nsew signal input
rlabel metal2 s 12162 31200 12218 32400 6 mprj_we_o_user
port 1108 nsew signal output
rlabel metal3 s 379200 8576 380400 8696 6 user1_vcc_powergood
port 1109 nsew signal output
rlabel metal3 s 379200 11024 380400 11144 6 user1_vdd_powergood
port 1110 nsew signal output
rlabel metal3 s 379200 13472 380400 13592 6 user2_vcc_powergood
port 1111 nsew signal output
rlabel metal3 s 379200 15920 380400 16040 6 user2_vdd_powergood
port 1112 nsew signal output
rlabel metal2 s 8482 31200 8538 32400 6 user_clock
port 1113 nsew signal output
rlabel metal2 s 369122 31200 369178 32400 6 user_clock2
port 1114 nsew signal output
rlabel metal3 s 379200 18368 380400 18488 6 user_irq[0]
port 1115 nsew signal output
rlabel metal3 s 379200 20816 380400 20936 6 user_irq[1]
port 1116 nsew signal output
rlabel metal3 s 379200 23264 380400 23384 6 user_irq[2]
port 1117 nsew signal output
rlabel metal2 s 369858 31200 369914 32400 6 user_irq_core[0]
port 1118 nsew signal input
rlabel metal2 s 370594 31200 370650 32400 6 user_irq_core[1]
port 1119 nsew signal input
rlabel metal2 s 371330 31200 371386 32400 6 user_irq_core[2]
port 1120 nsew signal input
rlabel metal3 s 379200 25712 380400 25832 6 user_irq_ena[0]
port 1121 nsew signal input
rlabel metal3 s 379200 28160 380400 28280 6 user_irq_ena[1]
port 1122 nsew signal input
rlabel metal3 s 379200 30608 380400 30728 6 user_irq_ena[2]
port 1123 nsew signal input
rlabel metal2 s 9218 31200 9274 32400 6 user_reset
port 1124 nsew signal output
rlabel metal4 s 5014 1040 5194 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 20064 1040 20244 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 35114 1040 35294 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 50164 1040 50344 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 65214 1040 65394 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 80264 1040 80444 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 95314 1040 95494 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 110364 1040 110544 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 125414 1040 125594 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 140464 1040 140644 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 155514 1040 155694 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 170564 1040 170744 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 185614 1040 185794 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 200664 1040 200844 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 215714 1040 215894 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 230764 1040 230944 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 245814 1040 245994 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 260864 1040 261044 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 275914 1040 276094 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 290964 1040 291144 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 306014 1040 306194 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 321064 1040 321244 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 336114 1040 336294 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 351164 1040 351344 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 366214 1040 366394 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 141284 1040 141464 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 156334 1040 156514 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 171384 1040 171564 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 186434 1040 186614 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 66854 1040 67034 30512 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 76854 1040 77034 30512 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 255814 1040 255994 30512 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 270864 1040 271044 30512 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 256614 1040 256794 30512 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 271664 1040 271844 30512 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 263194 1040 263374 30512 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 278244 1040 278424 30512 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 263994 1040 264174 30512 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 279044 1040 279224 30512 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 12394 1040 12574 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 27444 1040 27624 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 42494 1040 42674 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 57544 1040 57724 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 72594 1040 72774 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 87644 1040 87824 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 102694 1040 102874 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 117744 1040 117924 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 132794 1040 132974 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 147844 1040 148024 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 162894 1040 163074 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 177944 1040 178124 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 192994 1040 193174 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 208044 1040 208224 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 223094 1040 223274 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 238144 1040 238324 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 253194 1040 253374 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 268244 1040 268424 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 283294 1040 283474 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 298344 1040 298524 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 313394 1040 313574 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 328444 1040 328624 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 343494 1040 343674 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 358544 1040 358724 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 373594 1040 373774 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 148664 1040 148844 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 163714 1040 163894 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 178764 1040 178944 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 193814 1040 193994 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 71034 1040 71214 30512 6 vssd2
port 1134 nsew ground bidirectional
rlabel metal4 s 81034 1040 81214 30512 6 vssd2
port 1134 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 380000 32000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23108758
string GDS_FILE /openlane/designs/mgmt_protect/runs/THE_ONLY_RUN_2/results/signoff/mgmt_protect.magic.gds
string GDS_START 687408
<< end >>

