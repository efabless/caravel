magic
tech sky130A
magscale 1 2
timestamp 1636130125
<< locali >>
rect 2697 8823 2731 8993
rect 765 6851 799 7361
rect 6193 5763 6227 5865
rect 2697 2091 2731 5049
rect 2789 3451 2823 5049
rect 2881 2839 2915 5117
rect 4629 3383 4663 3485
rect 2789 1547 2823 2329
rect 9965 1751 9999 2601
<< viali >>
rect 1501 11305 1535 11339
rect 2881 11305 2915 11339
rect 3157 11305 3191 11339
rect 4261 11305 4295 11339
rect 5457 11305 5491 11339
rect 5917 11305 5951 11339
rect 6285 11305 6319 11339
rect 6561 11305 6595 11339
rect 7389 11305 7423 11339
rect 7665 11305 7699 11339
rect 7849 11305 7883 11339
rect 8401 11305 8435 11339
rect 8769 11305 8803 11339
rect 1869 11237 1903 11271
rect 3433 11237 3467 11271
rect 3801 11237 3835 11271
rect 7021 11237 7055 11271
rect 9413 11237 9447 11271
rect 1317 11101 1351 11135
rect 1593 11101 1627 11135
rect 2053 11101 2087 11135
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 3249 11101 3283 11135
rect 3617 11101 3651 11135
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 5089 11101 5123 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7573 11101 7607 11135
rect 8125 11101 8159 11135
rect 8585 11101 8619 11135
rect 8953 11101 8987 11135
rect 9321 11101 9355 11135
rect 4445 11033 4479 11067
rect 1777 10965 1811 10999
rect 2329 10965 2363 10999
rect 2605 10965 2639 10999
rect 3893 10965 3927 10999
rect 4813 10965 4847 10999
rect 4905 10965 4939 10999
rect 9137 10965 9171 10999
rect 1685 10761 1719 10795
rect 1961 10761 1995 10795
rect 2329 10761 2363 10795
rect 2789 10761 2823 10795
rect 8953 10761 8987 10795
rect 5641 10693 5675 10727
rect 5825 10693 5859 10727
rect 8585 10693 8619 10727
rect 1225 10625 1259 10659
rect 1501 10625 1535 10659
rect 1777 10625 1811 10659
rect 2053 10625 2087 10659
rect 2513 10625 2547 10659
rect 2605 10625 2639 10659
rect 3341 10625 3375 10659
rect 3525 10625 3559 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 6009 10625 6043 10659
rect 6561 10625 6595 10659
rect 8033 10625 8067 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 6193 10557 6227 10591
rect 9413 10557 9447 10591
rect 1409 10489 1443 10523
rect 2881 10489 2915 10523
rect 8493 10489 8527 10523
rect 2237 10421 2271 10455
rect 3065 10421 3099 10455
rect 4905 10421 4939 10455
rect 5365 10421 5399 10455
rect 9045 10421 9079 10455
rect 1685 10217 1719 10251
rect 8125 10217 8159 10251
rect 9137 10217 9171 10251
rect 9413 10149 9447 10183
rect 3709 10081 3743 10115
rect 4077 10081 4111 10115
rect 6009 10081 6043 10115
rect 7849 10081 7883 10115
rect 1409 10013 1443 10047
rect 3433 10013 3467 10047
rect 5549 10013 5583 10047
rect 8401 10013 8435 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 3157 9945 3191 9979
rect 7573 9945 7607 9979
rect 1317 9877 1351 9911
rect 1593 9877 1627 9911
rect 6101 9877 6135 9911
rect 7941 9877 7975 9911
rect 8493 9877 8527 9911
rect 1777 9673 1811 9707
rect 2513 9673 2547 9707
rect 6837 9673 6871 9707
rect 1317 9605 1351 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 2697 9537 2731 9571
rect 4629 9537 4663 9571
rect 5641 9537 5675 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 7113 9537 7147 9571
rect 7665 9537 7699 9571
rect 9505 9537 9539 9571
rect 2789 9469 2823 9503
rect 3157 9469 3191 9503
rect 5089 9469 5123 9503
rect 7205 9469 7239 9503
rect 9137 9469 9171 9503
rect 2421 9401 2455 9435
rect 1593 9333 1627 9367
rect 2145 9333 2179 9367
rect 5273 9333 5307 9367
rect 5457 9333 5491 9367
rect 5825 9333 5859 9367
rect 7021 9333 7055 9367
rect 1501 9129 1535 9163
rect 2513 9129 2547 9163
rect 2973 9129 3007 9163
rect 3801 9129 3835 9163
rect 4813 9129 4847 9163
rect 9413 9129 9447 9163
rect 3617 9061 3651 9095
rect 2697 8993 2731 9027
rect 5365 8993 5399 9027
rect 1317 8925 1351 8959
rect 1593 8925 1627 8959
rect 1869 8925 1903 8959
rect 2145 8925 2179 8959
rect 2605 8925 2639 8959
rect 2789 8925 2823 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 5089 8925 5123 8959
rect 7389 8925 7423 8959
rect 8769 8925 8803 8959
rect 3249 8857 3283 8891
rect 3433 8857 3467 8891
rect 4905 8857 4939 8891
rect 5641 8857 5675 8891
rect 8125 8857 8159 8891
rect 1777 8789 1811 8823
rect 2053 8789 2087 8823
rect 2329 8789 2363 8823
rect 2697 8789 2731 8823
rect 3065 8789 3099 8823
rect 5273 8789 5307 8823
rect 7113 8789 7147 8823
rect 1501 8585 1535 8619
rect 5917 8585 5951 8619
rect 7205 8585 7239 8619
rect 1317 8449 1351 8483
rect 2203 8449 2237 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7665 8449 7699 8483
rect 9505 8449 9539 8483
rect 2329 8381 2363 8415
rect 4169 8381 4203 8415
rect 4445 8381 4479 8415
rect 9137 8381 9171 8415
rect 1593 8245 1627 8279
rect 2586 8245 2620 8279
rect 4077 8245 4111 8279
rect 6837 8245 6871 8279
rect 7113 8245 7147 8279
rect 1317 8041 1351 8075
rect 8217 8041 8251 8075
rect 5181 7905 5215 7939
rect 5549 7905 5583 7939
rect 1409 7837 1443 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 5089 7837 5123 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 8309 7837 8343 7871
rect 8769 7837 8803 7871
rect 3157 7769 3191 7803
rect 4445 7769 4479 7803
rect 1501 7701 1535 7735
rect 1685 7701 1719 7735
rect 4261 7701 4295 7735
rect 7481 7701 7515 7735
rect 8493 7701 8527 7735
rect 9413 7701 9447 7735
rect 8585 7497 8619 7531
rect 1409 7429 1443 7463
rect 1593 7429 1627 7463
rect 5641 7429 5675 7463
rect 5917 7429 5951 7463
rect 6193 7429 6227 7463
rect 7941 7429 7975 7463
rect 765 7361 799 7395
rect 1685 7361 1719 7395
rect 2605 7361 2639 7395
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 5733 7361 5767 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 9045 7361 9079 7395
rect 2329 7293 2363 7327
rect 2973 7293 3007 7327
rect 9137 7293 9171 7327
rect 9229 7293 9263 7327
rect 8401 7225 8435 7259
rect 4905 7157 4939 7191
rect 8677 7157 8711 7191
rect 1409 6953 1443 6987
rect 1942 6953 1976 6987
rect 5917 6953 5951 6987
rect 6732 6953 6766 6987
rect 765 6817 799 6851
rect 1674 6817 1708 6851
rect 3985 6817 4019 6851
rect 6469 6817 6503 6851
rect 8217 6817 8251 6851
rect 9321 6817 9355 6851
rect 1593 6749 1627 6783
rect 3617 6749 3651 6783
rect 5457 6749 5491 6783
rect 8309 6749 8343 6783
rect 6009 6681 6043 6715
rect 6193 6681 6227 6715
rect 3433 6613 3467 6647
rect 6377 6613 6411 6647
rect 8493 6613 8527 6647
rect 8769 6613 8803 6647
rect 9137 6613 9171 6647
rect 9229 6613 9263 6647
rect 1501 6409 1535 6443
rect 4905 6409 4939 6443
rect 5273 6409 5307 6443
rect 2697 6341 2731 6375
rect 1317 6273 1351 6307
rect 1593 6273 1627 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 4261 6273 4295 6307
rect 5089 6273 5123 6307
rect 6009 6273 6043 6307
rect 6653 6273 6687 6307
rect 8677 6273 8711 6307
rect 9229 6273 9263 6307
rect 2421 6205 2455 6239
rect 4169 6205 4203 6239
rect 6193 6205 6227 6239
rect 6837 6205 6871 6239
rect 7205 6205 7239 6239
rect 2145 6137 2179 6171
rect 1777 6069 1811 6103
rect 2053 6069 2087 6103
rect 5365 6069 5399 6103
rect 6377 6069 6411 6103
rect 9137 6069 9171 6103
rect 9413 6069 9447 6103
rect 1685 5865 1719 5899
rect 1961 5865 1995 5899
rect 2973 5865 3007 5899
rect 3617 5865 3651 5899
rect 3801 5865 3835 5899
rect 6193 5865 6227 5899
rect 6377 5865 6411 5899
rect 8769 5865 8803 5899
rect 1593 5797 1627 5831
rect 2697 5797 2731 5831
rect 4261 5729 4295 5763
rect 6193 5729 6227 5763
rect 8585 5729 8619 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 2145 5661 2179 5695
rect 2421 5661 2455 5695
rect 2881 5661 2915 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 6285 5661 6319 5695
rect 9413 5661 9447 5695
rect 4537 5593 4571 5627
rect 8309 5593 8343 5627
rect 2329 5525 2363 5559
rect 2605 5525 2639 5559
rect 6009 5525 6043 5559
rect 6745 5525 6779 5559
rect 6837 5525 6871 5559
rect 5089 5321 5123 5355
rect 3341 5185 3375 5219
rect 5273 5185 5307 5219
rect 6193 5185 6227 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 8861 5185 8895 5219
rect 2881 5117 2915 5151
rect 3617 5117 3651 5151
rect 5825 5117 5859 5151
rect 8125 5117 8159 5151
rect 8677 5117 8711 5151
rect 2697 5049 2731 5083
rect 2789 5049 2823 5083
rect 2789 3417 2823 3451
rect 8493 5049 8527 5083
rect 5365 4981 5399 5015
rect 5733 4981 5767 5015
rect 9321 4981 9355 5015
rect 3985 4777 4019 4811
rect 4537 4777 4571 4811
rect 8493 4777 8527 4811
rect 9413 4777 9447 4811
rect 4169 4641 4203 4675
rect 6285 4641 6319 4675
rect 8769 4641 8803 4675
rect 3617 4573 3651 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 8585 4573 8619 4607
rect 5917 4505 5951 4539
rect 6561 4505 6595 4539
rect 9045 4505 9079 4539
rect 3433 4437 3467 4471
rect 4813 4437 4847 4471
rect 4905 4437 4939 4471
rect 6101 4437 6135 4471
rect 8033 4437 8067 4471
rect 8125 4437 8159 4471
rect 8953 4437 8987 4471
rect 8677 4233 8711 4267
rect 3341 4097 3375 4131
rect 3985 4097 4019 4131
rect 5457 4097 5491 4131
rect 6009 4097 6043 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 7481 4097 7515 4131
rect 8585 4097 8619 4131
rect 9045 4097 9079 4131
rect 3617 4029 3651 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 3525 3961 3559 3995
rect 8125 3961 8159 3995
rect 5917 3893 5951 3927
rect 7389 3893 7423 3927
rect 8401 3893 8435 3927
rect 3525 3689 3559 3723
rect 3801 3689 3835 3723
rect 4537 3689 4571 3723
rect 4905 3689 4939 3723
rect 5089 3689 5123 3723
rect 6101 3689 6135 3723
rect 8861 3689 8895 3723
rect 9229 3689 9263 3723
rect 4077 3621 4111 3655
rect 4169 3553 4203 3587
rect 6929 3553 6963 3587
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 3893 3485 3927 3519
rect 4353 3485 4387 3519
rect 4629 3485 4663 3519
rect 4721 3485 4755 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 6561 3485 6595 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 4629 3349 4663 3383
rect 5549 3349 5583 3383
rect 5733 3349 5767 3383
rect 6469 3349 6503 3383
rect 8585 3349 8619 3383
rect 9413 3349 9447 3383
rect 9413 3145 9447 3179
rect 8677 3077 8711 3111
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4261 3009 4295 3043
rect 6101 3009 6135 3043
rect 7481 3009 7515 3043
rect 7573 3009 7607 3043
rect 8033 3009 8067 3043
rect 8309 3009 8343 3043
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 4629 2941 4663 2975
rect 8125 2941 8159 2975
rect 3525 2873 3559 2907
rect 4077 2873 4111 2907
rect 6837 2873 6871 2907
rect 2881 2805 2915 2839
rect 3801 2805 3835 2839
rect 6561 2805 6595 2839
rect 3525 2601 3559 2635
rect 3801 2601 3835 2635
rect 4077 2601 4111 2635
rect 4537 2601 4571 2635
rect 5089 2601 5123 2635
rect 5549 2601 5583 2635
rect 6101 2601 6135 2635
rect 7021 2601 7055 2635
rect 8125 2601 8159 2635
rect 8585 2601 8619 2635
rect 9045 2601 9079 2635
rect 9965 2601 9999 2635
rect 4169 2533 4203 2567
rect 4813 2533 4847 2567
rect 5825 2533 5859 2567
rect 6193 2533 6227 2567
rect 3341 2397 3375 2431
rect 3617 2397 3651 2431
rect 3893 2397 3927 2431
rect 4353 2393 4387 2427
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 5365 2397 5399 2431
rect 5917 2397 5951 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 6837 2397 6871 2431
rect 7297 2397 7331 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8309 2397 8343 2431
rect 8769 2397 8803 2431
rect 8861 2397 8895 2431
rect 9229 2397 9263 2431
rect 2697 2057 2731 2091
rect 2789 2329 2823 2363
rect 7113 2329 7147 2363
rect 7481 2329 7515 2363
rect 8401 2329 8435 2363
rect 5181 2261 5215 2295
rect 6469 2261 6503 2295
rect 7573 2261 7607 2295
rect 9413 2261 9447 2295
rect 3525 2057 3559 2091
rect 3801 2057 3835 2091
rect 4353 2057 4387 2091
rect 4905 2057 4939 2091
rect 6837 2057 6871 2091
rect 7849 2057 7883 2091
rect 8125 2057 8159 2091
rect 8309 2057 8343 2091
rect 8585 2057 8619 2091
rect 9413 2057 9447 2091
rect 4445 1989 4479 2023
rect 5089 1989 5123 2023
rect 3341 1921 3375 1955
rect 3617 1921 3651 1955
rect 4077 1921 4111 1955
rect 4169 1921 4203 1955
rect 6653 1921 6687 1955
rect 7665 1921 7699 1955
rect 7941 1921 7975 1955
rect 8493 1921 8527 1955
rect 8769 1921 8803 1955
rect 9045 1921 9079 1955
rect 9229 1921 9263 1955
rect 4721 1853 4755 1887
rect 5365 1853 5399 1887
rect 3893 1785 3927 1819
rect 8861 1785 8895 1819
rect 5181 1717 5215 1751
rect 9965 1717 9999 1751
rect 2789 1513 2823 1547
rect 9045 1513 9079 1547
rect 3525 1445 3559 1479
rect 4445 1445 4479 1479
rect 4629 1377 4663 1411
rect 9413 1377 9447 1411
rect 3341 1309 3375 1343
rect 3617 1309 3651 1343
rect 3893 1309 3927 1343
rect 4261 1309 4295 1343
rect 8125 1309 8159 1343
rect 8301 1309 8335 1343
rect 8677 1309 8711 1343
rect 8953 1309 8987 1343
rect 4169 1241 4203 1275
rect 3801 1173 3835 1207
rect 7941 1173 7975 1207
rect 8493 1173 8527 1207
rect 8861 1173 8895 1207
rect 9229 1173 9263 1207
<< metal1 >>
rect 2406 11908 2412 11960
rect 2464 11948 2470 11960
rect 8662 11948 8668 11960
rect 2464 11920 8668 11948
rect 2464 11908 2470 11920
rect 8662 11908 8668 11920
rect 8720 11908 8726 11960
rect 2958 11772 2964 11824
rect 3016 11812 3022 11824
rect 8294 11812 8300 11824
rect 3016 11784 8300 11812
rect 3016 11772 3022 11784
rect 8294 11772 8300 11784
rect 8352 11772 8358 11824
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 6914 11744 6920 11756
rect 1544 11716 6920 11744
rect 1544 11704 1550 11716
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 10410 11744 10416 11756
rect 8444 11716 10416 11744
rect 8444 11704 8450 11716
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 3418 11636 3424 11688
rect 3476 11676 3482 11688
rect 6086 11676 6092 11688
rect 3476 11648 6092 11676
rect 3476 11636 3482 11648
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 16666 11676 16672 11688
rect 6236 11648 16672 11676
rect 6236 11636 6242 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 1302 11568 1308 11620
rect 1360 11608 1366 11620
rect 6270 11608 6276 11620
rect 1360 11580 6276 11608
rect 1360 11568 1366 11580
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 9858 11608 9864 11620
rect 7432 11580 9864 11608
rect 7432 11568 7438 11580
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 7650 11540 7656 11552
rect 3568 11512 7656 11540
rect 3568 11500 3574 11512
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 9766 11540 9772 11552
rect 7800 11512 9772 11540
rect 7800 11500 7806 11512
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 5858 11450
rect 5910 11398 5922 11450
rect 5974 11398 8766 11450
rect 8818 11398 8830 11450
rect 8882 11398 8894 11450
rect 8946 11398 8958 11450
rect 9010 11398 9022 11450
rect 9074 11398 9844 11450
rect 920 11376 9844 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2958 11336 2964 11348
rect 2915 11308 2964 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 4249 11339 4307 11345
rect 3191 11308 4016 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3602 11268 3608 11280
rect 3467 11240 3608 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 1302 11132 1308 11144
rect 1263 11104 1308 11132
rect 1302 11092 1308 11104
rect 1360 11092 1366 11144
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 1872 11132 1900 11231
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 3789 11271 3847 11277
rect 3789 11237 3801 11271
rect 3835 11237 3847 11271
rect 3988 11268 4016 11308
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4614 11336 4620 11348
rect 4295 11308 4620 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4614 11296 4620 11308
rect 4672 11336 4678 11348
rect 5166 11336 5172 11348
rect 4672 11308 5172 11336
rect 4672 11296 4678 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5905 11339 5963 11345
rect 5905 11305 5917 11339
rect 5951 11336 5963 11339
rect 6178 11336 6184 11348
rect 5951 11308 6184 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6546 11336 6552 11348
rect 6328 11308 6373 11336
rect 6507 11308 6552 11336
rect 6328 11296 6334 11308
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7650 11336 7656 11348
rect 7611 11308 7656 11336
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8386 11336 8392 11348
rect 8347 11308 8392 11336
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8628 11308 8769 11336
rect 8628 11296 8634 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 3988 11240 4844 11268
rect 3789 11231 3847 11237
rect 3510 11200 3516 11212
rect 2700 11172 3516 11200
rect 2038 11132 2044 11144
rect 1627 11104 1900 11132
rect 1999 11104 2044 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 2406 11132 2412 11144
rect 2188 11104 2233 11132
rect 2367 11104 2412 11132
rect 2188 11092 2194 11104
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2700 11141 2728 11172
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 3804 11200 3832 11231
rect 4816 11200 4844 11240
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 6730 11268 6736 11280
rect 5592 11240 6736 11268
rect 5592 11228 5598 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7742 11268 7748 11280
rect 7055 11240 7748 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 8478 11228 8484 11280
rect 8536 11268 8542 11280
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 8536 11240 9413 11268
rect 8536 11228 8542 11240
rect 9401 11237 9413 11240
rect 9447 11268 9459 11271
rect 9447 11240 9628 11268
rect 9447 11237 9459 11240
rect 9401 11231 9459 11237
rect 9490 11200 9496 11212
rect 3804 11172 4752 11200
rect 4816 11172 9496 11200
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2685 11095 2743 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3418 11132 3424 11144
rect 3283 11104 3424 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3602 11132 3608 11144
rect 3563 11104 3608 11132
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 4614 11132 4620 11144
rect 4387 11104 4476 11132
rect 4575 11104 4620 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 934 11024 940 11076
rect 992 11064 998 11076
rect 1854 11064 1860 11076
rect 992 11036 1860 11064
rect 992 11024 998 11036
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 1946 11024 1952 11076
rect 2004 11064 2010 11076
rect 4448 11073 4476 11104
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4433 11067 4491 11073
rect 2004 11036 3924 11064
rect 2004 11024 2010 11036
rect 1762 10996 1768 11008
rect 1723 10968 1768 10996
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 2406 10996 2412 11008
rect 2363 10968 2412 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 2593 10999 2651 11005
rect 2593 10965 2605 10999
rect 2639 10996 2651 10999
rect 3510 10996 3516 11008
rect 2639 10968 3516 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3896 11005 3924 11036
rect 4433 11033 4445 11067
rect 4479 11064 4491 11067
rect 4522 11064 4528 11076
rect 4479 11036 4528 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 4724 11064 4752 11172
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 9600 11144 9628 11240
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5258 11132 5264 11144
rect 5123 11104 5264 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5626 11132 5632 11144
rect 5587 11104 5632 11132
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5776 11104 5821 11132
rect 5776 11092 5782 11104
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6420 11104 6745 11132
rect 6420 11092 6426 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7558 11132 7564 11144
rect 6880 11104 6925 11132
rect 7519 11104 7564 11132
rect 6880 11092 6886 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8444 11104 8585 11132
rect 8444 11092 8450 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 9122 11132 9128 11144
rect 8987 11104 9128 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9582 11132 9588 11144
rect 9355 11104 9588 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9214 11064 9220 11076
rect 4724 11036 9220 11064
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 3881 10999 3939 11005
rect 3881 10965 3893 10999
rect 3927 10965 3939 10999
rect 3881 10959 3939 10965
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4801 10999 4859 11005
rect 4801 10996 4813 10999
rect 4028 10968 4813 10996
rect 4028 10956 4034 10968
rect 4801 10965 4813 10968
rect 4847 10965 4859 10999
rect 4801 10959 4859 10965
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 4948 10968 4993 10996
rect 4948 10956 4954 10968
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 6822 10996 6828 11008
rect 5592 10968 6828 10996
rect 5592 10956 5598 10968
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 9122 10996 9128 11008
rect 9083 10968 9128 10996
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 920 10906 9844 10928
rect 920 10854 4116 10906
rect 4168 10854 4180 10906
rect 4232 10854 4244 10906
rect 4296 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 7216 10906
rect 7268 10854 7280 10906
rect 7332 10854 7344 10906
rect 7396 10854 7408 10906
rect 7460 10854 7472 10906
rect 7524 10854 9844 10906
rect 920 10832 9844 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1912 10764 1961 10792
rect 1912 10752 1918 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2188 10764 2329 10792
rect 2188 10752 2194 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 2317 10755 2375 10761
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 2958 10792 2964 10804
rect 2823 10764 2964 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3108 10764 8064 10792
rect 3108 10752 3114 10764
rect 1578 10724 1584 10736
rect 1228 10696 1584 10724
rect 1228 10665 1256 10696
rect 1578 10684 1584 10696
rect 1636 10684 1642 10736
rect 5629 10727 5687 10733
rect 5629 10724 5641 10727
rect 1780 10696 5641 10724
rect 1780 10665 1808 10696
rect 5629 10693 5641 10696
rect 5675 10693 5687 10727
rect 5629 10687 5687 10693
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 5859 10696 6132 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 1213 10659 1271 10665
rect 1213 10625 1225 10659
rect 1259 10625 1271 10659
rect 1213 10619 1271 10625
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 1118 10548 1124 10600
rect 1176 10588 1182 10600
rect 1504 10588 1532 10619
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 2004 10628 2053 10656
rect 2004 10616 2010 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2501 10659 2559 10665
rect 2501 10656 2513 10659
rect 2188 10628 2513 10656
rect 2188 10616 2194 10628
rect 2501 10625 2513 10628
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2958 10656 2964 10668
rect 2639 10628 2964 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 1176 10560 1532 10588
rect 1176 10548 1182 10560
rect 1394 10520 1400 10532
rect 1355 10492 1400 10520
rect 1394 10480 1400 10492
rect 1452 10480 1458 10532
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 2869 10523 2927 10529
rect 1636 10492 2820 10520
rect 1636 10480 1642 10492
rect 2222 10452 2228 10464
rect 2183 10424 2228 10452
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2792 10452 2820 10492
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3142 10520 3148 10532
rect 2915 10492 3148 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 3344 10520 3372 10619
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3476 10628 3525 10656
rect 3476 10616 3482 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4203 10628 4261 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4764 10628 4997 10656
rect 4764 10616 4770 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 5166 10656 5172 10668
rect 5127 10628 5172 10656
rect 4985 10619 5043 10625
rect 5166 10616 5172 10628
rect 5224 10656 5230 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5224 10628 6009 10656
rect 5224 10616 5230 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 6104 10656 6132 10696
rect 6914 10684 6920 10736
rect 6972 10684 6978 10736
rect 6362 10656 6368 10668
rect 6104 10628 6368 10656
rect 5997 10619 6055 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 8036 10665 8064 10764
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8720 10764 8953 10792
rect 8720 10752 8726 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 8168 10696 8585 10724
rect 8168 10684 8174 10696
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 8573 10687 8631 10693
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8021 10619 8079 10625
rect 8128 10628 8769 10656
rect 3804 10588 3832 10616
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 3804 10560 6193 10588
rect 6181 10557 6193 10560
rect 6227 10557 6239 10591
rect 8128 10588 8156 10628
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 6181 10551 6239 10557
rect 8036 10560 8156 10588
rect 3786 10520 3792 10532
rect 3344 10492 3792 10520
rect 3786 10480 3792 10492
rect 3844 10520 3850 10532
rect 4706 10520 4712 10532
rect 3844 10492 4712 10520
rect 3844 10480 3850 10492
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 8036 10520 8064 10560
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 9232 10588 9260 10619
rect 9398 10588 9404 10600
rect 8720 10560 9260 10588
rect 9359 10560 9404 10588
rect 8720 10548 8726 10560
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 7892 10492 8064 10520
rect 7892 10480 7898 10492
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 8481 10523 8539 10529
rect 8168 10492 8340 10520
rect 8168 10480 8174 10492
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2792 10424 3065 10452
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 3384 10424 4905 10452
rect 3384 10412 3390 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 4893 10415 4951 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 8202 10452 8208 10464
rect 6236 10424 8208 10452
rect 6236 10412 6242 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8312 10452 8340 10492
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 9582 10520 9588 10532
rect 8527 10492 9588 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8312 10424 9045 10452
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 9033 10415 9091 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 5858 10362
rect 5910 10310 5922 10362
rect 5974 10310 8766 10362
rect 8818 10310 8830 10362
rect 8882 10310 8894 10362
rect 8946 10310 8958 10362
rect 9010 10310 9022 10362
rect 9074 10310 9844 10362
rect 920 10288 9844 10310
rect 15194 10276 15200 10328
rect 15252 10316 15258 10328
rect 16574 10316 16580 10328
rect 15252 10288 16580 10316
rect 15252 10276 15258 10288
rect 16574 10276 16580 10288
rect 16632 10276 16638 10328
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1762 10248 1768 10260
rect 1719 10220 1768 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1762 10208 1768 10220
rect 1820 10248 1826 10260
rect 3418 10248 3424 10260
rect 1820 10220 3424 10248
rect 1820 10208 1826 10220
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 5644 10220 7788 10248
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 2464 10084 3709 10112
rect 2464 10072 2470 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4706 10112 4712 10124
rect 4111 10084 4712 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 1854 10044 1860 10056
rect 1636 10016 1860 10044
rect 1636 10004 1642 10016
rect 1854 10004 1860 10016
rect 1912 10044 1918 10056
rect 1912 10016 2070 10044
rect 1912 10004 1918 10016
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 5534 10044 5540 10056
rect 3476 10016 3521 10044
rect 5495 10016 5540 10044
rect 3476 10004 3482 10016
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 3145 9979 3203 9985
rect 3145 9945 3157 9979
rect 3191 9976 3203 9979
rect 3694 9976 3700 9988
rect 3191 9948 3700 9976
rect 3191 9945 3203 9948
rect 3145 9939 3203 9945
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 1302 9908 1308 9920
rect 1263 9880 1308 9908
rect 1302 9868 1308 9880
rect 1360 9868 1366 9920
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2222 9868 2228 9920
rect 2280 9908 2286 9920
rect 4448 9908 4476 9962
rect 2280 9880 4476 9908
rect 2280 9868 2286 9880
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5644 9908 5672 10220
rect 7760 10180 7788 10220
rect 7834 10208 7840 10260
rect 7892 10248 7898 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 7892 10220 8125 10248
rect 7892 10208 7898 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8260 10220 9137 10248
rect 8260 10208 8266 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 7760 10152 9413 10180
rect 9401 10149 9413 10152
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10112 6055 10115
rect 7466 10112 7472 10124
rect 6043 10084 7472 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7834 10112 7840 10124
rect 7747 10084 7840 10112
rect 7834 10072 7840 10084
rect 7892 10112 7898 10124
rect 7892 10084 9260 10112
rect 7892 10072 7898 10084
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6328 10016 6486 10044
rect 6328 10004 6334 10016
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 7984 10016 8401 10044
rect 7984 10004 7990 10016
rect 8389 10013 8401 10016
rect 8435 10044 8447 10047
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 8435 10016 8769 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8757 10013 8769 10016
rect 8803 10013 8815 10047
rect 8938 10044 8944 10056
rect 8899 10016 8944 10044
rect 8757 10007 8815 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9232 10053 9260 10084
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 6104 9976 6132 10004
rect 6104 9948 6316 9976
rect 6086 9908 6092 9920
rect 4672 9880 5672 9908
rect 6047 9880 6092 9908
rect 4672 9868 4678 9880
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6288 9908 6316 9948
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 7524 9948 7573 9976
rect 7524 9936 7530 9948
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 7561 9939 7619 9945
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 6288 9880 7941 9908
rect 7929 9877 7941 9880
rect 7975 9877 7987 9911
rect 8478 9908 8484 9920
rect 8439 9880 8484 9908
rect 7929 9871 7987 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 920 9818 9844 9840
rect 920 9766 4116 9818
rect 4168 9766 4180 9818
rect 4232 9766 4244 9818
rect 4296 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 7216 9818
rect 7268 9766 7280 9818
rect 7332 9766 7344 9818
rect 7396 9766 7408 9818
rect 7460 9766 7472 9818
rect 7524 9766 9844 9818
rect 920 9744 9844 9766
rect 1765 9707 1823 9713
rect 1765 9673 1777 9707
rect 1811 9704 1823 9707
rect 2130 9704 2136 9716
rect 1811 9676 2136 9704
rect 1811 9673 1823 9676
rect 1765 9667 1823 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 2501 9707 2559 9713
rect 2501 9673 2513 9707
rect 2547 9673 2559 9707
rect 2501 9667 2559 9673
rect 1302 9636 1308 9648
rect 1215 9608 1308 9636
rect 1302 9596 1308 9608
rect 1360 9636 1366 9648
rect 1360 9608 1716 9636
rect 1360 9596 1366 9608
rect 1688 9580 1716 9608
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 1084 9540 1409 9568
rect 1084 9528 1090 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1397 9531 1455 9537
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2516 9568 2544 9667
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 6086 9704 6092 9716
rect 3752 9676 6092 9704
rect 3752 9664 3758 9676
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6604 9676 6837 9704
rect 6604 9664 6610 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 8202 9704 8208 9716
rect 7760 9686 8208 9704
rect 6825 9667 6883 9673
rect 3510 9596 3516 9648
rect 3568 9596 3574 9648
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 5534 9636 5540 9648
rect 4948 9608 5540 9636
rect 4948 9596 4954 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5644 9608 7236 9636
rect 7742 9634 7748 9686
rect 7800 9676 8208 9686
rect 7800 9634 7806 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 22094 9704 22100 9716
rect 21416 9676 22100 9704
rect 21416 9664 21422 9676
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 8312 9622 8340 9664
rect 2271 9540 2544 9568
rect 2685 9571 2743 9577
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 2958 9568 2964 9580
rect 2731 9540 2964 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1964 9500 1992 9531
rect 2700 9500 2728 9531
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 5644 9577 5672 9608
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4488 9540 4629 9568
rect 4488 9528 4494 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5960 9540 6009 9568
rect 5960 9528 5966 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 6144 9540 6193 9568
rect 6144 9528 6150 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6328 9540 7113 9568
rect 6328 9528 6334 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 1360 9472 2728 9500
rect 2777 9503 2835 9509
rect 1360 9460 1366 9472
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3326 9500 3332 9512
rect 3191 9472 3332 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 2792 9432 2820 9463
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5718 9500 5724 9512
rect 5123 9472 5724 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 6822 9500 6828 9512
rect 5828 9472 6828 9500
rect 2455 9404 2820 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1946 9364 1952 9376
rect 1627 9336 1952 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 3602 9364 3608 9376
rect 2179 9336 3608 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5442 9364 5448 9376
rect 5403 9336 5448 9364
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5828 9373 5856 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7116 9432 7144 9531
rect 7208 9509 7236 9608
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 9490 9568 9496 9580
rect 9451 9540 9496 9568
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 9171 9472 9444 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 7116 9404 8248 9432
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6144 9336 7021 9364
rect 6144 9324 6150 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7650 9364 7656 9376
rect 7156 9336 7656 9364
rect 7156 9324 7162 9336
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8220 9364 8248 9404
rect 9416 9376 9444 9472
rect 8478 9364 8484 9376
rect 8220 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9398 9324 9404 9376
rect 9456 9324 9462 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 5858 9274
rect 5910 9222 5922 9274
rect 5974 9222 8766 9274
rect 8818 9222 8830 9274
rect 8882 9222 8894 9274
rect 8946 9222 8958 9274
rect 9010 9222 9022 9274
rect 9074 9222 9844 9274
rect 920 9200 9844 9222
rect 1486 9160 1492 9172
rect 1447 9132 1492 9160
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2501 9163 2559 9169
rect 2501 9160 2513 9163
rect 2096 9132 2513 9160
rect 2096 9120 2102 9132
rect 2501 9129 2513 9132
rect 2547 9129 2559 9163
rect 2501 9123 2559 9129
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3510 9160 3516 9172
rect 3007 9132 3516 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3694 9120 3700 9172
rect 3752 9160 3758 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3752 9132 3801 9160
rect 3752 9120 3758 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 3605 9095 3663 9101
rect 3605 9092 3617 9095
rect 1596 9064 3617 9092
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1596 8965 1624 9064
rect 3605 9061 3617 9064
rect 3651 9061 3663 9095
rect 3804 9092 3832 9123
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 4801 9163 4859 9169
rect 4801 9160 4813 9163
rect 4764 9132 4813 9160
rect 4764 9120 4770 9132
rect 4801 9129 4813 9132
rect 4847 9129 4859 9163
rect 4801 9123 4859 9129
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 9398 9160 9404 9172
rect 5316 9132 7972 9160
rect 9359 9132 9404 9160
rect 5316 9120 5322 9132
rect 3804 9064 5120 9092
rect 3605 9055 3663 9061
rect 4724 9036 4752 9064
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 2685 9027 2743 9033
rect 1728 8996 2636 9024
rect 1728 8984 1734 8996
rect 2608 8968 2636 8996
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 4430 9024 4436 9036
rect 2731 8996 4436 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4706 8984 4712 9036
rect 4764 8984 4770 9036
rect 1305 8959 1363 8965
rect 1305 8956 1317 8959
rect 900 8928 1317 8956
rect 900 8916 906 8928
rect 1305 8925 1317 8928
rect 1351 8925 1363 8959
rect 1305 8919 1363 8925
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1581 8919 1639 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 3142 8956 3148 8968
rect 2823 8928 3148 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3602 8956 3608 8968
rect 3252 8928 3608 8956
rect 2498 8888 2504 8900
rect 1780 8860 2504 8888
rect 1780 8829 1808 8860
rect 2498 8848 2504 8860
rect 2556 8848 2562 8900
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 3252 8897 3280 8928
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 5092 8965 5120 9064
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 6914 9024 6920 9036
rect 5399 8996 6920 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 6914 8984 6920 8996
rect 6972 9024 6978 9036
rect 7834 9024 7840 9036
rect 6972 8996 7840 9024
rect 6972 8984 6978 8996
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3712 8928 4077 8956
rect 3712 8900 3740 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7944 8956 7972 9132
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 7423 8928 8248 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 2924 8860 3249 8888
rect 2924 8848 2930 8860
rect 3237 8857 3249 8860
rect 3283 8857 3295 8891
rect 3237 8851 3295 8857
rect 3421 8891 3479 8897
rect 3421 8857 3433 8891
rect 3467 8888 3479 8891
rect 3694 8888 3700 8900
rect 3467 8860 3700 8888
rect 3467 8857 3479 8860
rect 3421 8851 3479 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4172 8888 4200 8919
rect 4890 8888 4896 8900
rect 4028 8860 4200 8888
rect 4851 8860 4896 8888
rect 4028 8848 4034 8860
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5902 8888 5908 8900
rect 5675 8860 5908 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6086 8848 6092 8900
rect 6144 8848 6150 8900
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 7064 8860 8125 8888
rect 7064 8848 7070 8860
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8220 8888 8248 8928
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8536 8928 8769 8956
rect 8536 8916 8542 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 9674 8888 9680 8900
rect 8220 8860 9680 8888
rect 8113 8851 8171 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8789 1823 8823
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 1765 8783 1823 8789
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2363 8792 2697 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 5166 8820 5172 8832
rect 3099 8792 5172 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5261 8823 5319 8829
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 6638 8820 6644 8832
rect 5307 8792 6644 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 8662 8820 8668 8832
rect 7892 8792 8668 8820
rect 7892 8780 7898 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 920 8730 9844 8752
rect 920 8678 4116 8730
rect 4168 8678 4180 8730
rect 4232 8678 4244 8730
rect 4296 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 7216 8730
rect 7268 8678 7280 8730
rect 7332 8678 7344 8730
rect 7396 8678 7408 8730
rect 7460 8678 7472 8730
rect 7524 8678 9844 8730
rect 920 8656 9844 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 1854 8616 1860 8628
rect 1535 8588 1860 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 3418 8616 3424 8628
rect 2424 8588 3424 8616
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 2424 8548 2452 8588
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 5718 8616 5724 8628
rect 3568 8588 5724 8616
rect 3568 8576 3574 8588
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5902 8616 5908 8628
rect 5863 8588 5908 8616
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7558 8616 7564 8628
rect 7239 8588 7564 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 9950 8616 9956 8628
rect 7760 8588 9956 8616
rect 2372 8520 2452 8548
rect 2372 8508 2378 8520
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 2924 8520 3082 8548
rect 2924 8508 2930 8520
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 4764 8520 4922 8548
rect 4764 8508 4770 8520
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 7760 8548 7788 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 6880 8520 7788 8548
rect 6880 8508 6886 8520
rect 8018 8508 8024 8560
rect 8076 8508 8082 8560
rect 1302 8480 1308 8492
rect 1263 8452 1308 8480
rect 1302 8440 1308 8452
rect 1360 8440 1366 8492
rect 2191 8483 2249 8489
rect 2191 8480 2203 8483
rect 1780 8452 2203 8480
rect 1780 8424 1808 8452
rect 2191 8449 2203 8452
rect 2237 8449 2249 8483
rect 2191 8443 2249 8449
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5960 8452 6193 8480
rect 5960 8440 5966 8452
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6696 8452 6929 8480
rect 6696 8440 6702 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 1762 8372 1768 8424
rect 1820 8372 1826 8424
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 3234 8412 3240 8424
rect 2648 8384 3240 8412
rect 2648 8372 2654 8384
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3660 8384 4169 8412
rect 3660 8372 3666 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4982 8412 4988 8424
rect 4479 8384 4988 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 7668 8412 7696 8443
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9272 8452 9505 8480
rect 9272 8440 9278 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 5776 8384 7696 8412
rect 5776 8372 5782 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8720 8384 9137 8412
rect 8720 8372 8726 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 1912 8316 2452 8344
rect 1912 8304 1918 8316
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8276 1639 8279
rect 1946 8276 1952 8288
rect 1627 8248 1952 8276
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2424 8276 2452 8316
rect 2574 8279 2632 8285
rect 2574 8276 2586 8279
rect 2424 8248 2586 8276
rect 2574 8245 2586 8248
rect 2620 8245 2632 8279
rect 2574 8239 2632 8245
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3970 8276 3976 8288
rect 3200 8248 3976 8276
rect 3200 8236 3206 8248
rect 3970 8236 3976 8248
rect 4028 8276 4034 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 4028 8248 4077 8276
rect 4028 8236 4034 8248
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4065 8239 4123 8245
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6052 8248 6837 8276
rect 6052 8236 6058 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 7064 8248 7113 8276
rect 7064 8236 7070 8248
rect 7101 8245 7113 8248
rect 7147 8245 7159 8279
rect 7101 8239 7159 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 5858 8186
rect 5910 8134 5922 8186
rect 5974 8134 8766 8186
rect 8818 8134 8830 8186
rect 8882 8134 8894 8186
rect 8946 8134 8958 8186
rect 9010 8134 9022 8186
rect 9074 8134 9844 8186
rect 920 8112 9844 8134
rect 1305 8075 1363 8081
rect 1305 8041 1317 8075
rect 1351 8072 1363 8075
rect 1670 8072 1676 8084
rect 1351 8044 1676 8072
rect 1351 8041 1363 8044
rect 1305 8035 1363 8041
rect 1412 7877 1440 8044
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 5166 8072 5172 8084
rect 3936 8044 5172 8072
rect 3936 8032 3942 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7834 8072 7840 8084
rect 7616 8044 7840 8072
rect 7616 8032 7622 8044
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8205 8075 8263 8081
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8478 8072 8484 8084
rect 8251 8044 8484 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9582 8072 9588 8084
rect 9272 8044 9588 8072
rect 9272 8032 9278 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 8110 8004 8116 8016
rect 6604 7976 8116 8004
rect 6604 7964 6610 7976
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 1636 7908 5181 7936
rect 1636 7896 1642 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 5994 7936 6000 7948
rect 5583 7908 6000 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 1544 7840 1992 7868
rect 1544 7828 1550 7840
rect 1026 7760 1032 7812
rect 1084 7800 1090 7812
rect 1504 7800 1532 7828
rect 1084 7772 1532 7800
rect 1964 7786 1992 7840
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3605 7871 3663 7877
rect 3476 7840 3521 7868
rect 3476 7828 3482 7840
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5626 7868 5632 7880
rect 5123 7840 5632 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 3142 7800 3148 7812
rect 3103 7772 3148 7800
rect 1084 7760 1090 7772
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 3620 7800 3648 7831
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7156 7840 7573 7868
rect 7156 7828 7162 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 3436 7772 3648 7800
rect 3436 7744 3464 7772
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 4433 7803 4491 7809
rect 4433 7800 4445 7803
rect 3936 7772 4445 7800
rect 3936 7760 3942 7772
rect 4433 7769 4445 7772
rect 4479 7769 4491 7803
rect 4433 7763 4491 7769
rect 5994 7760 6000 7812
rect 6052 7760 6058 7812
rect 8312 7800 8340 7831
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8536 7840 8769 7868
rect 8536 7828 8542 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 9490 7800 9496 7812
rect 6748 7772 8340 7800
rect 8496 7772 9496 7800
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 1673 7735 1731 7741
rect 1673 7732 1685 7735
rect 1636 7704 1685 7732
rect 1636 7692 1642 7704
rect 1673 7701 1685 7704
rect 1719 7732 1731 7735
rect 1762 7732 1768 7744
rect 1719 7704 1768 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 3418 7692 3424 7744
rect 3476 7692 3482 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4028 7704 4261 7732
rect 4028 7692 4034 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6454 7732 6460 7744
rect 5408 7704 6460 7732
rect 5408 7692 5414 7704
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 6748 7732 6776 7772
rect 6604 7704 6776 7732
rect 7469 7735 7527 7741
rect 6604 7692 6610 7704
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 7926 7732 7932 7744
rect 7515 7704 7932 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8496 7741 8524 7772
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 8481 7735 8539 7741
rect 8481 7701 8493 7735
rect 8527 7701 8539 7735
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 8481 7695 8539 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 920 7642 9844 7664
rect 920 7590 4116 7642
rect 4168 7590 4180 7642
rect 4232 7590 4244 7642
rect 4296 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 7216 7642
rect 7268 7590 7280 7642
rect 7332 7590 7344 7642
rect 7396 7590 7408 7642
rect 7460 7590 7472 7642
rect 7524 7590 9844 7642
rect 10686 7624 10692 7676
rect 10744 7664 10750 7676
rect 15194 7664 15200 7676
rect 10744 7636 15200 7664
rect 10744 7624 10750 7636
rect 15194 7624 15200 7636
rect 15252 7624 15258 7676
rect 20622 7664 20628 7676
rect 16546 7636 20628 7664
rect 920 7568 9844 7590
rect 11054 7556 11060 7608
rect 11112 7596 11118 7608
rect 16546 7596 16574 7636
rect 20622 7624 20628 7636
rect 20680 7624 20686 7676
rect 11112 7568 16574 7596
rect 11112 7556 11118 7568
rect 8573 7531 8631 7537
rect 1412 7500 5948 7528
rect 1412 7469 1440 7500
rect 1397 7463 1455 7469
rect 1397 7429 1409 7463
rect 1443 7429 1455 7463
rect 1397 7423 1455 7429
rect 1581 7463 1639 7469
rect 1581 7429 1593 7463
rect 1627 7460 1639 7463
rect 2314 7460 2320 7472
rect 1627 7432 2320 7460
rect 1627 7429 1639 7432
rect 1581 7423 1639 7429
rect 753 7395 811 7401
rect 753 7361 765 7395
rect 799 7392 811 7395
rect 1596 7392 1624 7423
rect 2314 7420 2320 7432
rect 2372 7420 2378 7472
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 5626 7460 5632 7472
rect 3292 7432 3358 7460
rect 5587 7432 5632 7460
rect 3292 7420 3298 7432
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 5920 7469 5948 7500
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 13814 7528 13820 7540
rect 8619 7500 13820 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 5951 7432 6193 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 6181 7429 6193 7432
rect 6227 7429 6239 7463
rect 6181 7423 6239 7429
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7460 7987 7463
rect 8588 7460 8616 7491
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 7975 7432 8616 7460
rect 7975 7429 7987 7432
rect 7929 7423 7987 7429
rect 799 7364 1624 7392
rect 1673 7395 1731 7401
rect 799 7361 811 7364
rect 753 7355 811 7361
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 1946 7392 1952 7404
rect 1719 7364 1952 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2096 7364 2605 7392
rect 2096 7352 2102 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4798 7392 4804 7404
rect 4479 7364 4804 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 6914 7392 6920 7404
rect 5767 7364 6920 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8021 7355 8079 7361
rect 8128 7364 8217 7392
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2363 7296 2973 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 8036 7324 8064 7355
rect 6236 7296 8064 7324
rect 6236 7284 6242 7296
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 2406 7256 2412 7268
rect 1820 7228 2412 7256
rect 1820 7216 1826 7228
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4798 7256 4804 7268
rect 4580 7228 4804 7256
rect 4580 7216 4586 7228
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 8128 7256 8156 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 9030 7392 9036 7404
rect 8991 7364 9036 7392
rect 8205 7355 8263 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8352 7296 9137 7324
rect 8352 7284 8358 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9272 7296 9317 7324
rect 9272 7284 9278 7296
rect 7248 7228 8156 7256
rect 8389 7259 8447 7265
rect 7248 7216 7254 7228
rect 8389 7225 8401 7259
rect 8435 7256 8447 7259
rect 9306 7256 9312 7268
rect 8435 7228 9312 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 750 7148 756 7200
rect 808 7188 814 7200
rect 3234 7188 3240 7200
rect 808 7160 3240 7188
rect 808 7148 814 7160
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 8018 7188 8024 7200
rect 4939 7160 8024 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8168 7160 8677 7188
rect 8168 7148 8174 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8665 7151 8723 7157
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 5858 7098
rect 5910 7046 5922 7098
rect 5974 7046 8766 7098
rect 8818 7046 8830 7098
rect 8882 7046 8894 7098
rect 8946 7046 8958 7098
rect 9010 7046 9022 7098
rect 9074 7046 9844 7098
rect 920 7024 9844 7046
rect 1302 6944 1308 6996
rect 1360 6984 1366 6996
rect 1397 6987 1455 6993
rect 1397 6984 1409 6987
rect 1360 6956 1409 6984
rect 1360 6944 1366 6956
rect 1397 6953 1409 6956
rect 1443 6953 1455 6987
rect 1397 6947 1455 6953
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 1930 6987 1988 6993
rect 1930 6984 1942 6987
rect 1636 6956 1942 6984
rect 1636 6944 1642 6956
rect 1930 6953 1942 6956
rect 1976 6953 1988 6987
rect 1930 6947 1988 6953
rect 5905 6987 5963 6993
rect 5905 6953 5917 6987
rect 5951 6984 5963 6987
rect 6546 6984 6552 6996
rect 5951 6956 6552 6984
rect 5951 6953 5963 6956
rect 5905 6947 5963 6953
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6720 6987 6778 6993
rect 6720 6953 6732 6987
rect 6766 6984 6778 6987
rect 7098 6984 7104 6996
rect 6766 6956 7104 6984
rect 6766 6953 6778 6956
rect 6720 6947 6778 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 5718 6876 5724 6928
rect 5776 6916 5782 6928
rect 6362 6916 6368 6928
rect 5776 6888 6368 6916
rect 5776 6876 5782 6888
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 8294 6876 8300 6928
rect 8352 6876 8358 6928
rect 753 6851 811 6857
rect 753 6817 765 6851
rect 799 6848 811 6851
rect 1662 6851 1720 6857
rect 1662 6848 1674 6851
rect 799 6820 1674 6848
rect 799 6817 811 6820
rect 753 6811 811 6817
rect 1662 6817 1674 6820
rect 1708 6817 1720 6851
rect 1662 6811 1720 6817
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 3973 6851 4031 6857
rect 2096 6820 3556 6848
rect 2096 6808 2102 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 1596 6706 1624 6743
rect 2038 6712 2044 6724
rect 1780 6706 2044 6712
rect 1596 6684 2044 6706
rect 1596 6678 1808 6684
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 1026 6604 1032 6656
rect 1084 6644 1090 6656
rect 2424 6644 2452 6698
rect 2590 6644 2596 6656
rect 1084 6616 2596 6644
rect 1084 6604 1090 6616
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3418 6644 3424 6656
rect 2740 6616 3424 6644
rect 2740 6604 2746 6616
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3528 6644 3556 6820
rect 3973 6817 3985 6851
rect 4019 6848 4031 6851
rect 4522 6848 4528 6860
rect 4019 6820 4528 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 6822 6848 6828 6860
rect 6503 6820 6828 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 8018 6808 8024 6860
rect 8076 6808 8082 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8312 6848 8340 6876
rect 8478 6848 8484 6860
rect 8251 6820 8484 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 5445 6783 5503 6789
rect 3660 6752 3705 6780
rect 3660 6740 3666 6752
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 8036 6780 8064 6808
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 5491 6752 6500 6780
rect 8036 6752 8309 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 4706 6672 4712 6724
rect 4764 6672 4770 6724
rect 5902 6672 5908 6724
rect 5960 6712 5966 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5960 6684 6009 6712
rect 5960 6672 5966 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6681 6239 6715
rect 6472 6712 6500 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 7006 6712 7012 6724
rect 6472 6684 7012 6712
rect 6181 6675 6239 6681
rect 5534 6644 5540 6656
rect 3528 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6196 6644 6224 6675
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7190 6672 7196 6724
rect 7248 6672 7254 6724
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8444 6684 8800 6712
rect 8444 6672 8450 6684
rect 5684 6616 6224 6644
rect 6365 6647 6423 6653
rect 5684 6604 5690 6616
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 7558 6644 7564 6656
rect 6411 6616 7564 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8478 6644 8484 6656
rect 8439 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8772 6653 8800 6684
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8904 6616 9137 6644
rect 8904 6604 8910 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9272 6616 9317 6644
rect 9272 6604 9278 6616
rect 920 6554 9844 6576
rect 920 6502 4116 6554
rect 4168 6502 4180 6554
rect 4232 6502 4244 6554
rect 4296 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 7216 6554
rect 7268 6502 7280 6554
rect 7332 6502 7344 6554
rect 7396 6502 7408 6554
rect 7460 6502 7472 6554
rect 7524 6502 9844 6554
rect 920 6480 9844 6502
rect 1302 6400 1308 6452
rect 1360 6400 1366 6452
rect 1489 6443 1547 6449
rect 1489 6409 1501 6443
rect 1535 6440 1547 6443
rect 1535 6412 4016 6440
rect 1535 6409 1547 6412
rect 1489 6403 1547 6409
rect 1320 6372 1348 6400
rect 2682 6372 2688 6384
rect 1320 6344 1624 6372
rect 2643 6344 2688 6372
rect 1302 6304 1308 6316
rect 1263 6276 1308 6304
rect 1302 6264 1308 6276
rect 1360 6264 1366 6316
rect 1596 6313 1624 6344
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 3142 6372 3148 6384
rect 2832 6344 3148 6372
rect 2832 6332 2838 6344
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 3988 6372 4016 6412
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4580 6412 4905 6440
rect 4580 6400 4586 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 4893 6403 4951 6409
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5994 6440 6000 6452
rect 5307 6412 6000 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7800 6412 9260 6440
rect 7800 6400 7806 6412
rect 4706 6372 4712 6384
rect 3988 6344 4712 6372
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 5902 6372 5908 6384
rect 4816 6344 5908 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2314 6304 2320 6316
rect 1903 6276 2176 6304
rect 2275 6276 2320 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2148 6177 2176 6276
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4028 6276 4261 6304
rect 4028 6264 4034 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 4816 6304 4844 6344
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 8628 6344 8708 6372
rect 8628 6332 8634 6344
rect 4488 6276 4844 6304
rect 5077 6307 5135 6313
rect 4488 6264 4494 6276
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5994 6304 6000 6316
rect 5123 6276 5534 6304
rect 5955 6276 6000 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 4157 6239 4215 6245
rect 2464 6208 2509 6236
rect 2464 6196 2470 6208
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4982 6236 4988 6248
rect 4203 6208 4988 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5506 6236 5534 6276
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6638 6304 6644 6316
rect 6328 6276 6644 6304
rect 6328 6264 6334 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 8680 6313 8708 6344
rect 9232 6313 9260 6412
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 5506 6208 6193 6236
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 7834 6236 7840 6248
rect 7239 6208 7840 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6137 2191 6171
rect 6840 6168 6868 6199
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 2133 6131 2191 6137
rect 3804 6140 6868 6168
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 1946 6100 1952 6112
rect 1811 6072 1952 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 3804 6100 3832 6140
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 2087 6072 3832 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4798 6100 4804 6112
rect 4028 6072 4804 6100
rect 4028 6060 4034 6072
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6100 5411 6103
rect 6178 6100 6184 6112
rect 5399 6072 6184 6100
rect 5399 6069 5411 6072
rect 5353 6063 5411 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 8864 6100 8892 6128
rect 7156 6072 8892 6100
rect 9125 6103 9183 6109
rect 7156 6060 7162 6072
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 9306 6100 9312 6112
rect 9171 6072 9312 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 16666 6100 16672 6112
rect 9447 6072 16672 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 5858 6010
rect 5910 5958 5922 6010
rect 5974 5958 8766 6010
rect 8818 5958 8830 6010
rect 8882 5958 8894 6010
rect 8946 5958 8958 6010
rect 9010 5958 9022 6010
rect 9074 5958 9844 6010
rect 920 5936 9844 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1673 5899 1731 5905
rect 1673 5896 1685 5899
rect 1452 5868 1685 5896
rect 1452 5856 1458 5868
rect 1673 5865 1685 5868
rect 1719 5865 1731 5899
rect 1673 5859 1731 5865
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 1949 5899 2007 5905
rect 1949 5896 1961 5899
rect 1912 5868 1961 5896
rect 1912 5856 1918 5868
rect 1949 5865 1961 5868
rect 1995 5865 2007 5899
rect 1949 5859 2007 5865
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2372 5868 2973 5896
rect 2372 5856 2378 5868
rect 1578 5828 1584 5840
rect 1539 5800 1584 5828
rect 1578 5788 1584 5800
rect 1636 5788 1642 5840
rect 2130 5788 2136 5840
rect 2188 5788 2194 5840
rect 2685 5831 2743 5837
rect 2685 5797 2697 5831
rect 2731 5797 2743 5831
rect 2685 5791 2743 5797
rect 2148 5760 2176 5788
rect 1412 5732 2176 5760
rect 1412 5701 1440 5732
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1544 5664 1869 5692
rect 1544 5652 1550 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 2004 5664 2145 5692
rect 2004 5652 2010 5664
rect 2133 5661 2145 5664
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 2700 5692 2728 5791
rect 2884 5701 2912 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3605 5899 3663 5905
rect 3605 5896 3617 5899
rect 3476 5868 3617 5896
rect 3476 5856 3482 5868
rect 3605 5865 3617 5868
rect 3651 5865 3663 5899
rect 3605 5859 3663 5865
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6362 5896 6368 5908
rect 6227 5868 6368 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 3142 5788 3148 5840
rect 3200 5828 3206 5840
rect 3804 5828 3832 5859
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 8570 5896 8576 5908
rect 7064 5868 8576 5896
rect 7064 5856 7070 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8720 5868 8769 5896
rect 8720 5856 8726 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 3200 5800 4384 5828
rect 3200 5788 3206 5800
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3660 5732 4261 5760
rect 3660 5720 3666 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4356 5760 4384 5800
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6638 5828 6644 5840
rect 5684 5800 6644 5828
rect 5684 5788 5690 5800
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 5166 5760 5172 5772
rect 4356 5732 5172 5760
rect 4249 5723 4307 5729
rect 5166 5720 5172 5732
rect 5224 5760 5230 5772
rect 5534 5760 5540 5772
rect 5224 5732 5540 5760
rect 5224 5720 5230 5732
rect 5534 5720 5540 5732
rect 5592 5760 5598 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5592 5732 6193 5760
rect 5592 5720 5598 5732
rect 6181 5729 6193 5732
rect 6227 5760 6239 5763
rect 6227 5732 6408 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 2455 5664 2728 5692
rect 2869 5695 2927 5701
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 2958 5692 2964 5704
rect 2915 5664 2964 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 3191 5664 3341 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 4065 5695 4123 5701
rect 3476 5664 3521 5692
rect 3476 5652 3482 5664
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 4065 5655 4123 5661
rect 1210 5584 1216 5636
rect 1268 5624 1274 5636
rect 3510 5624 3516 5636
rect 1268 5596 1900 5624
rect 1268 5584 1274 5596
rect 1872 5568 1900 5596
rect 2332 5596 3516 5624
rect 1854 5516 1860 5568
rect 1912 5516 1918 5568
rect 2332 5565 2360 5596
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 4080 5624 4108 5655
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6380 5692 6408 5732
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 6914 5760 6920 5772
rect 6604 5732 6920 5760
rect 6604 5720 6610 5732
rect 6914 5720 6920 5732
rect 6972 5760 6978 5772
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 6972 5732 8585 5760
rect 6972 5720 6978 5732
rect 8573 5729 8585 5732
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 7190 5692 7196 5704
rect 6380 5664 7196 5692
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 9398 5692 9404 5704
rect 9359 5664 9404 5692
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 4430 5624 4436 5636
rect 4080 5596 4436 5624
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5525 2375 5559
rect 2590 5556 2596 5568
rect 2551 5528 2596 5556
rect 2317 5519 2375 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 4080 5556 4108 5596
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5593 4583 5627
rect 4525 5587 4583 5593
rect 2924 5528 4108 5556
rect 4540 5556 4568 5587
rect 5166 5584 5172 5636
rect 5224 5584 5230 5636
rect 6362 5624 6368 5636
rect 5920 5596 6368 5624
rect 5920 5556 5948 5596
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 8294 5624 8300 5636
rect 6748 5596 7052 5624
rect 8255 5596 8300 5624
rect 4540 5528 5948 5556
rect 5997 5559 6055 5565
rect 2924 5516 2930 5528
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6454 5556 6460 5568
rect 6043 5528 6460 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 6748 5565 6776 5596
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7024 5556 7052 5596
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 9858 5556 9864 5568
rect 6880 5528 6925 5556
rect 7024 5528 9864 5556
rect 6880 5516 6886 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 920 5466 9844 5488
rect 920 5414 4116 5466
rect 4168 5414 4180 5466
rect 4232 5414 4244 5466
rect 4296 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 7216 5466
rect 7268 5414 7280 5466
rect 7332 5414 7344 5466
rect 7396 5414 7408 5466
rect 7460 5414 7472 5466
rect 7524 5414 9844 5466
rect 920 5392 9844 5414
rect 5074 5352 5080 5364
rect 5035 5324 5080 5352
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 9950 5352 9956 5364
rect 8168 5324 9956 5352
rect 8168 5312 8174 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 1118 5244 1124 5296
rect 1176 5284 1182 5296
rect 2498 5284 2504 5296
rect 1176 5256 2504 5284
rect 1176 5244 1182 5256
rect 2498 5244 2504 5256
rect 2556 5244 2562 5296
rect 3602 5284 3608 5296
rect 3344 5256 3608 5284
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 3344 5225 3372 5256
rect 3602 5244 3608 5256
rect 3660 5244 3666 5296
rect 6638 5244 6644 5296
rect 6696 5244 6702 5296
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 7800 5256 8892 5284
rect 7800 5244 7806 5256
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 2464 5188 3341 5216
rect 2464 5176 2470 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 5258 5216 5264 5228
rect 4738 5188 5120 5216
rect 5219 5188 5264 5216
rect 3329 5179 3387 5185
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3050 5148 3056 5160
rect 2915 5120 3056 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 4982 5148 4988 5160
rect 3651 5120 4988 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5092 5148 5120 5188
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 6178 5216 6184 5228
rect 6139 5188 6184 5216
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7156 5188 7665 5216
rect 7156 5176 7162 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7653 5179 7711 5185
rect 8128 5188 8309 5216
rect 5166 5148 5172 5160
rect 5092 5120 5172 5148
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 2685 5083 2743 5089
rect 2685 5080 2697 5083
rect 2372 5052 2697 5080
rect 2372 5040 2378 5052
rect 2685 5049 2697 5052
rect 2731 5049 2743 5083
rect 2685 5043 2743 5049
rect 2777 5083 2835 5089
rect 2777 5049 2789 5083
rect 2823 5080 2835 5083
rect 3326 5080 3332 5092
rect 2823 5052 3332 5080
rect 2823 5049 2835 5052
rect 2777 5043 2835 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 3418 5012 3424 5024
rect 3200 4984 3424 5012
rect 3200 4972 3206 4984
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 3602 4972 3608 5024
rect 3660 5012 3666 5024
rect 4890 5012 4896 5024
rect 3660 4984 4896 5012
rect 3660 4972 3666 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5092 5012 5120 5120
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 8128 5157 8156 5188
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 8478 5216 8484 5228
rect 8343 5188 8484 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8864 5225 8892 5256
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8444 5120 8677 5148
rect 8444 5108 8450 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 8527 5052 16574 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 16546 5024 16574 5052
rect 5353 5015 5411 5021
rect 5353 5012 5365 5015
rect 5040 4984 5365 5012
rect 5040 4972 5046 4984
rect 5353 4981 5365 4984
rect 5399 4981 5411 5015
rect 5353 4975 5411 4981
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6086 5012 6092 5024
rect 5767 4984 6092 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 9582 5012 9588 5024
rect 9355 4984 9588 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 16546 4984 16580 5024
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 3036 4922 9844 4944
rect 3036 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 5858 4922
rect 5910 4870 5922 4922
rect 5974 4870 8766 4922
rect 8818 4870 8830 4922
rect 8882 4870 8894 4922
rect 8946 4870 8958 4922
rect 9010 4870 9022 4922
rect 9074 4870 9844 4922
rect 3036 4848 9844 4870
rect 3973 4811 4031 4817
rect 3973 4777 3985 4811
rect 4019 4808 4031 4811
rect 4522 4808 4528 4820
rect 4019 4780 4528 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 8202 4808 8208 4820
rect 4764 4780 8208 4808
rect 4764 4768 4770 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8662 4808 8668 4820
rect 8527 4780 8668 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 3142 4740 3148 4752
rect 2832 4712 3148 4740
rect 2832 4700 2838 4712
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 5166 4740 5172 4752
rect 3712 4712 5172 4740
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 2774 4604 2780 4616
rect 1728 4576 2780 4604
rect 1728 4564 1734 4576
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3712 4613 3740 4712
rect 5166 4700 5172 4712
rect 5224 4700 5230 4752
rect 5276 4712 5948 4740
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4798 4672 4804 4684
rect 4203 4644 4804 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5276 4672 5304 4712
rect 5040 4644 5304 4672
rect 5368 4644 5764 4672
rect 5040 4632 5046 4644
rect 3605 4607 3663 4613
rect 3605 4604 3617 4607
rect 3016 4576 3617 4604
rect 3016 4564 3022 4576
rect 3605 4573 3617 4576
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4573 3755 4607
rect 3697 4567 3755 4573
rect 1026 4496 1032 4548
rect 1084 4536 1090 4548
rect 3620 4536 3648 4567
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4120 4576 4353 4604
rect 4120 4564 4126 4576
rect 4341 4573 4353 4576
rect 4387 4604 4399 4607
rect 5368 4604 5396 4644
rect 5534 4604 5540 4616
rect 4387 4576 5396 4604
rect 5495 4576 5540 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5736 4613 5764 4644
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 4522 4536 4528 4548
rect 1084 4508 3004 4536
rect 3620 4508 4528 4536
rect 1084 4496 1090 4508
rect 2976 4480 3004 4508
rect 4522 4496 4528 4508
rect 4580 4496 4586 4548
rect 5920 4545 5948 4712
rect 8570 4700 8576 4752
rect 8628 4740 8634 4752
rect 8628 4712 9260 4740
rect 8628 4700 8634 4712
rect 9232 4684 9260 4712
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6546 4672 6552 4684
rect 6319 4644 6552 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8202 4672 8208 4684
rect 8076 4644 8208 4672
rect 8076 4632 8082 4644
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 8757 4675 8815 4681
rect 8757 4672 8769 4675
rect 8260 4644 8769 4672
rect 8260 4632 8266 4644
rect 8757 4641 8769 4644
rect 8803 4641 8815 4675
rect 8757 4635 8815 4641
rect 9214 4632 9220 4684
rect 9272 4632 9278 4684
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9766 4604 9772 4616
rect 8619 4576 9772 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 5905 4539 5963 4545
rect 4816 4508 5580 4536
rect 2958 4428 2964 4480
rect 3016 4428 3022 4480
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 4816 4477 4844 4508
rect 5552 4480 5580 4508
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 5951 4508 6500 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 6472 4480 6500 4508
rect 6546 4496 6552 4548
rect 6604 4536 6610 4548
rect 6604 4508 6649 4536
rect 6604 4496 6610 4508
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 3384 4440 3433 4468
rect 3384 4428 3390 4440
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4437 4859 4471
rect 4801 4431 4859 4437
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 4982 4468 4988 4480
rect 4939 4440 4988 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5534 4428 5540 4480
rect 5592 4428 5598 4480
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6362 4468 6368 4480
rect 6135 4440 6368 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 7024 4468 7052 4522
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9033 4539 9091 4545
rect 9033 4536 9045 4539
rect 8904 4508 9045 4536
rect 8904 4496 8910 4508
rect 9033 4505 9045 4508
rect 9079 4505 9091 4539
rect 9033 4499 9091 4505
rect 6512 4440 7052 4468
rect 6512 4428 6518 4440
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7984 4440 8033 4468
rect 7984 4428 7990 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 8938 4468 8944 4480
rect 8168 4440 8213 4468
rect 8899 4440 8944 4468
rect 8168 4428 8174 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 3036 4378 9844 4400
rect 3036 4326 4116 4378
rect 4168 4326 4180 4378
rect 4232 4326 4244 4378
rect 4296 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 7216 4378
rect 7268 4326 7280 4378
rect 7332 4326 7344 4378
rect 7396 4326 7408 4378
rect 7460 4326 7472 4378
rect 7524 4326 9844 4378
rect 3036 4304 9844 4326
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 8110 4264 8116 4276
rect 6788 4236 8116 4264
rect 6788 4224 6794 4236
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 8665 4267 8723 4273
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 8938 4264 8944 4276
rect 8711 4236 8944 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 4430 4156 4436 4208
rect 4488 4156 4494 4208
rect 7742 4196 7748 4208
rect 7484 4168 7748 4196
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 4948 4100 5457 4128
rect 4948 4088 4954 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5994 4128 6000 4140
rect 5955 4100 6000 4128
rect 5445 4091 5503 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 7484 4137 7512 4168
rect 7742 4156 7748 4168
rect 7800 4196 7806 4208
rect 7926 4196 7932 4208
rect 7800 4168 7932 4196
rect 7800 4156 7806 4168
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8036 4168 9674 4196
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 6604 4100 6653 4128
rect 6604 4088 6610 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 8036 4128 8064 4168
rect 8570 4128 8576 4140
rect 7469 4091 7527 4097
rect 7576 4100 8064 4128
rect 8531 4100 8576 4128
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 3620 3992 3648 4023
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6748 4060 6776 4091
rect 6328 4032 6776 4060
rect 6328 4020 6334 4032
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7576 4060 7604 4100
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8720 4100 9045 4128
rect 8720 4088 8726 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 7248 4032 7604 4060
rect 7248 4020 7254 4032
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8846 4060 8852 4072
rect 7984 4032 8852 4060
rect 7984 4020 7990 4032
rect 8846 4020 8852 4032
rect 8904 4060 8910 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8904 4032 9137 4060
rect 8904 4020 8910 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9490 4060 9496 4072
rect 9355 4032 9496 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 3559 3964 3648 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 5626 3952 5632 4004
rect 5684 3952 5690 4004
rect 8113 3995 8171 4001
rect 8113 3961 8125 3995
rect 8159 3992 8171 3995
rect 9030 3992 9036 4004
rect 8159 3964 9036 3992
rect 8159 3961 8171 3964
rect 8113 3955 8171 3961
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9646 3992 9674 4168
rect 10042 3992 10048 4004
rect 9646 3964 10048 3992
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3602 3924 3608 3936
rect 3384 3896 3608 3924
rect 3384 3884 3390 3896
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 5644 3924 5672 3952
rect 4212 3896 5672 3924
rect 5905 3927 5963 3933
rect 4212 3884 4218 3896
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6454 3924 6460 3936
rect 5951 3896 6460 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 6972 3896 7389 3924
rect 6972 3884 6978 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 16574 3924 16580 3936
rect 8435 3896 16580 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 3036 3834 9844 3856
rect 3036 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 5858 3834
rect 5910 3782 5922 3834
rect 5974 3782 8766 3834
rect 8818 3782 8830 3834
rect 8882 3782 8894 3834
rect 8946 3782 8958 3834
rect 9010 3782 9022 3834
rect 9074 3782 9844 3834
rect 3036 3760 9844 3782
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3108 3692 3525 3720
rect 3108 3680 3114 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 3513 3683 3571 3689
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 4246 3720 4252 3732
rect 3835 3692 4252 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 4488 3692 4537 3720
rect 4488 3680 4494 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4890 3720 4896 3732
rect 4851 3692 4896 3720
rect 4525 3683 4583 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5074 3720 5080 3732
rect 5035 3692 5080 3720
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 5920 3692 6101 3720
rect 3602 3652 3608 3664
rect 3344 3624 3608 3652
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3344 3525 3372 3624
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 4062 3652 4068 3664
rect 4023 3624 4068 3652
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 5092 3652 5120 3680
rect 5920 3664 5948 3692
rect 6089 3689 6101 3692
rect 6135 3720 6147 3723
rect 6546 3720 6552 3732
rect 6135 3692 6552 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8628 3692 8861 3720
rect 8628 3680 8634 3692
rect 8849 3689 8861 3692
rect 8895 3689 8907 3723
rect 8849 3683 8907 3689
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9306 3720 9312 3732
rect 9263 3692 9312 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 4264 3624 5120 3652
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 3804 3556 4169 3584
rect 3804 3528 3832 3556
rect 4157 3553 4169 3556
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3292 3488 3341 3516
rect 3292 3476 3298 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3786 3516 3792 3528
rect 3651 3488 3792 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 4264 3516 4292 3624
rect 5902 3612 5908 3664
rect 5960 3612 5966 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8754 3652 8760 3664
rect 8260 3624 8760 3652
rect 8260 3612 8266 3624
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 4798 3584 4804 3596
rect 4356 3556 4804 3584
rect 4356 3525 4384 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5920 3584 5948 3612
rect 6914 3584 6920 3596
rect 5368 3556 5948 3584
rect 6875 3556 6920 3584
rect 3927 3488 4292 3516
rect 4341 3519 4399 3525
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4663 3488 4721 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4709 3479 4767 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5368 3525 5396 3556
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 9232 3584 9260 3683
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 8628 3556 9260 3584
rect 8628 3544 8634 3556
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5592 3488 5917 3516
rect 5592 3476 5598 3488
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 6546 3516 6552 3528
rect 6507 3488 6552 3516
rect 5997 3479 6055 3485
rect 2777 3451 2835 3457
rect 2777 3417 2789 3451
rect 2823 3448 2835 3451
rect 5074 3448 5080 3460
rect 2823 3420 5080 3448
rect 2823 3417 2835 3420
rect 2777 3411 2835 3417
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 5626 3408 5632 3460
rect 5684 3448 5690 3460
rect 6012 3448 6040 3479
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 7892 3488 8401 3516
rect 7892 3476 7898 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8536 3488 8953 3516
rect 8536 3476 8542 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 8202 3448 8208 3460
rect 5684 3420 6040 3448
rect 8050 3420 8208 3448
rect 5684 3408 5690 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 4617 3383 4675 3389
rect 4617 3349 4629 3383
rect 4663 3380 4675 3383
rect 5537 3383 5595 3389
rect 5537 3380 5549 3383
rect 4663 3352 5549 3380
rect 4663 3349 4675 3352
rect 4617 3343 4675 3349
rect 5537 3349 5549 3352
rect 5583 3349 5595 3383
rect 5718 3380 5724 3392
rect 5679 3352 5724 3380
rect 5537 3343 5595 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 8478 3380 8484 3392
rect 6503 3352 8484 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8662 3380 8668 3392
rect 8619 3352 8668 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 9364 3352 9413 3380
rect 9364 3340 9370 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 3036 3290 9844 3312
rect 3036 3238 4116 3290
rect 4168 3238 4180 3290
rect 4232 3238 4244 3290
rect 4296 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 7216 3290
rect 7268 3238 7280 3290
rect 7332 3238 7344 3290
rect 7396 3238 7408 3290
rect 7460 3238 7472 3290
rect 7524 3238 9844 3290
rect 3036 3216 9844 3238
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 3844 3148 7788 3176
rect 3844 3136 3850 3148
rect 5718 3068 5724 3120
rect 5776 3068 5782 3120
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 7282 3108 7288 3120
rect 5960 3080 7288 3108
rect 5960 3068 5966 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 3605 3003 3663 3009
rect 3620 2972 3648 3003
rect 3878 3000 3884 3012
rect 3936 3040 3942 3052
rect 4154 3040 4160 3052
rect 3936 3012 4160 3040
rect 3936 3000 3942 3012
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4430 3040 4436 3052
rect 4295 3012 4436 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6178 3040 6184 3052
rect 6135 3012 6184 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6880 3012 7481 3040
rect 6880 3000 6886 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7760 3040 7788 3148
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9088 3148 9413 3176
rect 9088 3136 9094 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 8665 3111 8723 3117
rect 7607 3012 7788 3040
rect 7852 3080 8156 3108
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 4617 2975 4675 2981
rect 3620 2944 4384 2972
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 3513 2907 3571 2913
rect 3513 2904 3525 2907
rect 2740 2876 3525 2904
rect 2740 2864 2746 2876
rect 3513 2873 3525 2876
rect 3559 2873 3571 2907
rect 3513 2867 3571 2873
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 3878 2904 3884 2916
rect 3660 2876 3884 2904
rect 3660 2864 3666 2876
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 4028 2876 4077 2904
rect 4028 2864 4034 2876
rect 4065 2873 4077 2876
rect 4111 2873 4123 2907
rect 4065 2867 4123 2873
rect 4356 2848 4384 2944
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4982 2972 4988 2984
rect 4663 2944 4988 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 6104 2944 6960 2972
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 3789 2839 3847 2845
rect 3789 2836 3801 2839
rect 2915 2808 3801 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 3789 2805 3801 2808
rect 3835 2805 3847 2839
rect 3789 2799 3847 2805
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 4798 2836 4804 2848
rect 4396 2808 4804 2836
rect 4396 2796 4402 2808
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5258 2836 5264 2848
rect 4948 2808 5264 2836
rect 4948 2796 4954 2808
rect 5258 2796 5264 2808
rect 5316 2836 5322 2848
rect 6104 2836 6132 2944
rect 6270 2864 6276 2916
rect 6328 2904 6334 2916
rect 6825 2907 6883 2913
rect 6825 2904 6837 2907
rect 6328 2876 6837 2904
rect 6328 2864 6334 2876
rect 6825 2873 6837 2876
rect 6871 2873 6883 2907
rect 6825 2867 6883 2873
rect 5316 2808 6132 2836
rect 6549 2839 6607 2845
rect 5316 2796 5322 2808
rect 6549 2805 6561 2839
rect 6595 2836 6607 2839
rect 6638 2836 6644 2848
rect 6595 2808 6644 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 6932 2836 6960 2944
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7650 2972 7656 2984
rect 7248 2944 7656 2972
rect 7248 2932 7254 2944
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7558 2904 7564 2916
rect 7064 2876 7564 2904
rect 7064 2864 7070 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 7852 2836 7880 3080
rect 8018 3040 8024 3052
rect 7979 3012 8024 3040
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8128 3040 8156 3080
rect 8665 3077 8677 3111
rect 8711 3108 8723 3111
rect 8938 3108 8944 3120
rect 8711 3080 8944 3108
rect 8711 3077 8723 3080
rect 8665 3071 8723 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8128 3012 8309 3040
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3040 8815 3043
rect 8846 3040 8852 3052
rect 8803 3012 8852 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2941 8171 2975
rect 8496 2972 8524 3003
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9214 3040 9220 3052
rect 9088 3012 9220 3040
rect 9088 3000 9094 3012
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 8662 2972 8668 2984
rect 8496 2944 8668 2972
rect 8113 2935 8171 2941
rect 8128 2848 8156 2935
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 6932 2808 7880 2836
rect 8110 2796 8116 2848
rect 8168 2796 8174 2848
rect 3036 2746 9844 2768
rect 3036 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 5858 2746
rect 5910 2694 5922 2746
rect 5974 2694 8766 2746
rect 8818 2694 8830 2746
rect 8882 2694 8894 2746
rect 8946 2694 8958 2746
rect 9010 2694 9022 2746
rect 9074 2694 9844 2746
rect 3036 2672 9844 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 3513 2635 3571 2641
rect 3513 2632 3525 2635
rect 3476 2604 3525 2632
rect 3476 2592 3482 2604
rect 3513 2601 3525 2604
rect 3559 2601 3571 2635
rect 3513 2595 3571 2601
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3660 2604 3801 2632
rect 3660 2592 3666 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 4062 2632 4068 2644
rect 4023 2604 4068 2632
rect 3789 2595 3847 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4890 2632 4896 2644
rect 4571 2604 4896 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5166 2632 5172 2644
rect 5123 2604 5172 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5994 2632 6000 2644
rect 5583 2604 6000 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6546 2632 6552 2644
rect 6135 2604 6552 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7098 2632 7104 2644
rect 7055 2604 7104 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7616 2604 8125 2632
rect 7616 2592 7622 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9214 2632 9220 2644
rect 9079 2604 9220 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 3326 2524 3332 2576
rect 3384 2564 3390 2576
rect 4157 2567 4215 2573
rect 4157 2564 4169 2567
rect 3384 2536 4169 2564
rect 3384 2524 3390 2536
rect 4157 2533 4169 2536
rect 4203 2533 4215 2567
rect 4157 2527 4215 2533
rect 4338 2524 4344 2576
rect 4396 2564 4402 2576
rect 4706 2564 4712 2576
rect 4396 2536 4712 2564
rect 4396 2524 4402 2536
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 5258 2564 5264 2576
rect 4847 2536 5264 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 5810 2564 5816 2576
rect 5771 2536 5816 2564
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 6178 2564 6184 2576
rect 6139 2536 6184 2564
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 6512 2536 7880 2564
rect 6512 2524 6518 2536
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 3786 2496 3792 2508
rect 2740 2468 3792 2496
rect 2740 2456 2746 2468
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 4488 2468 6684 2496
rect 4488 2456 4494 2468
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 2792 2400 3341 2428
rect 2792 2369 2820 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3476 2400 3617 2428
rect 3476 2388 3482 2400
rect 3605 2397 3617 2400
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 3927 2400 4016 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 2777 2363 2835 2369
rect 2777 2329 2789 2363
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 3602 2292 3608 2304
rect 3016 2264 3608 2292
rect 3016 2252 3022 2264
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 3988 2292 4016 2400
rect 4080 2422 4292 2428
rect 4341 2427 4399 2433
rect 4341 2422 4353 2427
rect 4080 2400 4353 2422
rect 4080 2372 4108 2400
rect 4264 2394 4353 2400
rect 4341 2393 4353 2394
rect 4387 2393 4399 2427
rect 4341 2387 4399 2393
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 4663 2400 4844 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 4062 2320 4068 2372
rect 4120 2320 4126 2372
rect 4816 2360 4844 2400
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5353 2431 5411 2437
rect 4948 2400 4993 2428
rect 4948 2388 4954 2400
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 5905 2431 5963 2437
rect 5399 2400 5856 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 5718 2360 5724 2372
rect 4816 2332 5724 2360
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 4982 2292 4988 2304
rect 3988 2264 4988 2292
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5534 2292 5540 2304
rect 5316 2264 5540 2292
rect 5316 2252 5322 2264
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 5828 2292 5856 2400
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 6362 2428 6368 2440
rect 6323 2400 6368 2428
rect 5905 2391 5963 2397
rect 5920 2360 5948 2391
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 6656 2437 6684 2468
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2397 6699 2431
rect 6822 2428 6828 2440
rect 6783 2400 6828 2428
rect 6641 2391 6699 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 5920 2332 6500 2360
rect 6086 2292 6092 2304
rect 5828 2264 6092 2292
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 6472 2301 6500 2332
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 7101 2363 7159 2369
rect 7101 2360 7113 2363
rect 6788 2332 7113 2360
rect 6788 2320 6794 2332
rect 7101 2329 7113 2332
rect 7147 2329 7159 2363
rect 7101 2323 7159 2329
rect 7469 2363 7527 2369
rect 7469 2329 7481 2363
rect 7515 2360 7527 2363
rect 7650 2360 7656 2372
rect 7515 2332 7656 2360
rect 7515 2329 7527 2332
rect 7469 2323 7527 2329
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 7852 2360 7880 2536
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 8588 2496 8616 2595
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 21358 2632 21364 2644
rect 9999 2604 21364 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 9122 2496 9128 2508
rect 8076 2468 8524 2496
rect 8588 2468 9128 2496
rect 8076 2456 8082 2468
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 8294 2428 8300 2440
rect 8255 2400 8300 2428
rect 7929 2391 7987 2397
rect 7760 2332 7880 2360
rect 7760 2304 7788 2332
rect 6457 2295 6515 2301
rect 6457 2261 6469 2295
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7561 2295 7619 2301
rect 7561 2292 7573 2295
rect 7064 2264 7573 2292
rect 7064 2252 7070 2264
rect 7561 2261 7573 2264
rect 7607 2261 7619 2295
rect 7561 2255 7619 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 7944 2292 7972 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8018 2320 8024 2372
rect 8076 2360 8082 2372
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 8076 2332 8401 2360
rect 8076 2320 8082 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8496 2360 8524 2468
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 8720 2400 8769 2428
rect 8720 2388 8726 2400
rect 8757 2397 8769 2400
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2397 8907 2431
rect 8849 2391 8907 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9766 2428 9772 2440
rect 9263 2400 9772 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 8864 2360 8892 2391
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 8496 2332 8892 2360
rect 8389 2323 8447 2329
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 16574 2360 16580 2372
rect 8996 2332 16580 2360
rect 8996 2320 9002 2332
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 9214 2292 9220 2304
rect 7944 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9401 2295 9459 2301
rect 9401 2261 9413 2295
rect 9447 2292 9459 2295
rect 16666 2292 16672 2304
rect 9447 2264 16672 2292
rect 9447 2261 9459 2264
rect 9401 2255 9459 2261
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 3036 2202 9844 2224
rect 3036 2150 4116 2202
rect 4168 2150 4180 2202
rect 4232 2150 4244 2202
rect 4296 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 7216 2202
rect 7268 2150 7280 2202
rect 7332 2150 7344 2202
rect 7396 2150 7408 2202
rect 7460 2150 7472 2202
rect 7524 2150 9844 2202
rect 3036 2128 9844 2150
rect 2685 2091 2743 2097
rect 2685 2057 2697 2091
rect 2731 2057 2743 2091
rect 2685 2051 2743 2057
rect 2700 2020 2728 2051
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 3513 2091 3571 2097
rect 3513 2088 3525 2091
rect 3200 2060 3525 2088
rect 3200 2048 3206 2060
rect 3513 2057 3525 2060
rect 3559 2057 3571 2091
rect 3786 2088 3792 2100
rect 3747 2060 3792 2088
rect 3513 2051 3571 2057
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 4341 2091 4399 2097
rect 4341 2057 4353 2091
rect 4387 2088 4399 2091
rect 4614 2088 4620 2100
rect 4387 2060 4620 2088
rect 4387 2057 4399 2060
rect 4341 2051 4399 2057
rect 4614 2048 4620 2060
rect 4672 2048 4678 2100
rect 4893 2091 4951 2097
rect 4893 2057 4905 2091
rect 4939 2088 4951 2091
rect 5350 2088 5356 2100
rect 4939 2060 5356 2088
rect 4939 2057 4951 2060
rect 4893 2051 4951 2057
rect 4433 2023 4491 2029
rect 2700 1992 4108 2020
rect 4080 1964 4108 1992
rect 4433 1989 4445 2023
rect 4479 2020 4491 2023
rect 4706 2020 4712 2032
rect 4479 1992 4712 2020
rect 4479 1989 4491 1992
rect 4433 1983 4491 1989
rect 4706 1980 4712 1992
rect 4764 1980 4770 2032
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 3329 1955 3387 1961
rect 3329 1952 3341 1955
rect 2740 1924 3341 1952
rect 2740 1912 2746 1924
rect 3329 1921 3341 1924
rect 3375 1921 3387 1955
rect 3602 1952 3608 1964
rect 3563 1924 3608 1952
rect 3329 1915 3387 1921
rect 3344 1884 3372 1915
rect 3602 1912 3608 1924
rect 3660 1912 3666 1964
rect 4062 1952 4068 1964
rect 3975 1924 4068 1952
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4157 1955 4215 1961
rect 4157 1921 4169 1955
rect 4203 1952 4215 1955
rect 4522 1952 4528 1964
rect 4203 1924 4528 1952
rect 4203 1921 4215 1924
rect 4157 1915 4215 1921
rect 4522 1912 4528 1924
rect 4580 1912 4586 1964
rect 4246 1884 4252 1896
rect 3344 1856 4252 1884
rect 4246 1844 4252 1856
rect 4304 1844 4310 1896
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1884 4767 1887
rect 4798 1884 4804 1896
rect 4755 1856 4804 1884
rect 4755 1853 4767 1856
rect 4709 1847 4767 1853
rect 4798 1844 4804 1856
rect 4856 1844 4862 1896
rect 3694 1776 3700 1828
rect 3752 1816 3758 1828
rect 3881 1819 3939 1825
rect 3881 1816 3893 1819
rect 3752 1788 3893 1816
rect 3752 1776 3758 1788
rect 3881 1785 3893 1788
rect 3927 1785 3939 1819
rect 3881 1779 3939 1785
rect 3970 1776 3976 1828
rect 4028 1816 4034 1828
rect 4908 1816 4936 2051
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 6825 2091 6883 2097
rect 6825 2057 6837 2091
rect 6871 2088 6883 2091
rect 7098 2088 7104 2100
rect 6871 2060 7104 2088
rect 6871 2057 6883 2060
rect 6825 2051 6883 2057
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 7834 2088 7840 2100
rect 7795 2060 7840 2088
rect 7834 2048 7840 2060
rect 7892 2048 7898 2100
rect 7926 2048 7932 2100
rect 7984 2088 7990 2100
rect 8113 2091 8171 2097
rect 8113 2088 8125 2091
rect 7984 2060 8125 2088
rect 7984 2048 7990 2060
rect 8113 2057 8125 2060
rect 8159 2057 8171 2091
rect 8113 2051 8171 2057
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 8297 2091 8355 2097
rect 8297 2088 8309 2091
rect 8260 2060 8309 2088
rect 8260 2048 8266 2060
rect 8297 2057 8309 2060
rect 8343 2057 8355 2091
rect 8297 2051 8355 2057
rect 8573 2091 8631 2097
rect 8573 2057 8585 2091
rect 8619 2088 8631 2091
rect 9030 2088 9036 2100
rect 8619 2060 9036 2088
rect 8619 2057 8631 2060
rect 8573 2051 8631 2057
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 9398 2088 9404 2100
rect 9359 2060 9404 2088
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 4982 1980 4988 2032
rect 5040 2020 5046 2032
rect 5077 2023 5135 2029
rect 5077 2020 5089 2023
rect 5040 1992 5089 2020
rect 5040 1980 5046 1992
rect 5077 1989 5089 1992
rect 5123 2020 5135 2023
rect 5442 2020 5448 2032
rect 5123 1992 5448 2020
rect 5123 1989 5135 1992
rect 5077 1983 5135 1989
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 5534 1980 5540 2032
rect 5592 2020 5598 2032
rect 6730 2020 6736 2032
rect 5592 1992 6736 2020
rect 5592 1980 5598 1992
rect 6730 1980 6736 1992
rect 6788 1980 6794 2032
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 9306 2020 9312 2032
rect 7616 1992 8800 2020
rect 7616 1980 7622 1992
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 6914 1952 6920 1964
rect 6687 1924 6920 1952
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 6914 1912 6920 1924
rect 6972 1912 6978 1964
rect 7650 1952 7656 1964
rect 7611 1924 7656 1952
rect 7650 1912 7656 1924
rect 7708 1912 7714 1964
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1952 7987 1955
rect 8018 1952 8024 1964
rect 7975 1924 8024 1952
rect 7975 1921 7987 1924
rect 7929 1915 7987 1921
rect 8018 1912 8024 1924
rect 8076 1912 8082 1964
rect 8478 1952 8484 1964
rect 8439 1924 8484 1952
rect 8478 1912 8484 1924
rect 8536 1912 8542 1964
rect 8772 1961 8800 1992
rect 9048 1992 9312 2020
rect 9048 1961 9076 1992
rect 9306 1980 9312 1992
rect 9364 1980 9370 2032
rect 8757 1955 8815 1961
rect 8757 1921 8769 1955
rect 8803 1921 8815 1955
rect 8757 1915 8815 1921
rect 9033 1955 9091 1961
rect 9033 1921 9045 1955
rect 9079 1921 9091 1955
rect 9033 1915 9091 1921
rect 9217 1955 9275 1961
rect 9217 1921 9229 1955
rect 9263 1921 9275 1955
rect 9217 1915 9275 1921
rect 5074 1844 5080 1896
rect 5132 1884 5138 1896
rect 5353 1887 5411 1893
rect 5353 1884 5365 1887
rect 5132 1856 5365 1884
rect 5132 1844 5138 1856
rect 5353 1853 5365 1856
rect 5399 1853 5411 1887
rect 5353 1847 5411 1853
rect 6730 1844 6736 1896
rect 6788 1884 6794 1896
rect 9232 1884 9260 1915
rect 6788 1856 9260 1884
rect 6788 1844 6794 1856
rect 4028 1788 4936 1816
rect 8849 1819 8907 1825
rect 4028 1776 4034 1788
rect 8849 1785 8861 1819
rect 8895 1816 8907 1819
rect 9490 1816 9496 1828
rect 8895 1788 9496 1816
rect 8895 1785 8907 1788
rect 8849 1779 8907 1785
rect 9490 1776 9496 1788
rect 9548 1776 9554 1828
rect 3602 1708 3608 1760
rect 3660 1748 3666 1760
rect 5169 1751 5227 1757
rect 5169 1748 5181 1751
rect 3660 1720 5181 1748
rect 3660 1708 3666 1720
rect 5169 1717 5181 1720
rect 5215 1717 5227 1751
rect 5169 1711 5227 1717
rect 5258 1708 5264 1760
rect 5316 1748 5322 1760
rect 9953 1751 10011 1757
rect 9953 1748 9965 1751
rect 5316 1720 9965 1748
rect 5316 1708 5322 1720
rect 9953 1717 9965 1720
rect 9999 1717 10011 1751
rect 9953 1711 10011 1717
rect 3036 1658 9844 1680
rect 3036 1606 5666 1658
rect 5718 1606 5730 1658
rect 5782 1606 5794 1658
rect 5846 1606 5858 1658
rect 5910 1606 5922 1658
rect 5974 1606 8766 1658
rect 8818 1606 8830 1658
rect 8882 1606 8894 1658
rect 8946 1606 8958 1658
rect 9010 1606 9022 1658
rect 9074 1606 9844 1658
rect 3036 1584 9844 1606
rect 2777 1547 2835 1553
rect 2777 1513 2789 1547
rect 2823 1544 2835 1547
rect 5166 1544 5172 1556
rect 2823 1516 5172 1544
rect 2823 1513 2835 1516
rect 2777 1507 2835 1513
rect 5166 1504 5172 1516
rect 5224 1544 5230 1556
rect 5224 1516 7052 1544
rect 5224 1504 5230 1516
rect 2866 1436 2872 1488
rect 2924 1476 2930 1488
rect 3513 1479 3571 1485
rect 3513 1476 3525 1479
rect 2924 1448 3525 1476
rect 2924 1436 2930 1448
rect 3513 1445 3525 1448
rect 3559 1445 3571 1479
rect 3513 1439 3571 1445
rect 4062 1436 4068 1488
rect 4120 1476 4126 1488
rect 4433 1479 4491 1485
rect 4433 1476 4445 1479
rect 4120 1448 4445 1476
rect 4120 1436 4126 1448
rect 4433 1445 4445 1448
rect 4479 1445 4491 1479
rect 7024 1476 7052 1516
rect 8110 1504 8116 1556
rect 8168 1544 8174 1556
rect 9033 1547 9091 1553
rect 9033 1544 9045 1547
rect 8168 1516 9045 1544
rect 8168 1504 8174 1516
rect 9033 1513 9045 1516
rect 9079 1513 9091 1547
rect 9033 1507 9091 1513
rect 10962 1476 10968 1488
rect 7024 1448 10968 1476
rect 4433 1439 4491 1445
rect 10962 1436 10968 1448
rect 11020 1436 11026 1488
rect 4617 1411 4675 1417
rect 4617 1408 4629 1411
rect 3528 1380 4629 1408
rect 3528 1352 3556 1380
rect 4617 1377 4629 1380
rect 4663 1377 4675 1411
rect 4617 1371 4675 1377
rect 8220 1380 8432 1408
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1340 3387 1343
rect 3510 1340 3516 1352
rect 3375 1312 3516 1340
rect 3375 1309 3387 1312
rect 3329 1303 3387 1309
rect 3510 1300 3516 1312
rect 3568 1300 3574 1352
rect 3602 1300 3608 1352
rect 3660 1340 3666 1352
rect 3878 1340 3884 1352
rect 3660 1312 3705 1340
rect 3839 1312 3884 1340
rect 3660 1300 3666 1312
rect 3878 1300 3884 1312
rect 3936 1300 3942 1352
rect 4246 1340 4252 1352
rect 4207 1312 4252 1340
rect 4246 1300 4252 1312
rect 4304 1300 4310 1352
rect 8113 1343 8171 1349
rect 8113 1309 8125 1343
rect 8159 1340 8171 1343
rect 8220 1340 8248 1380
rect 8159 1312 8248 1340
rect 8289 1343 8347 1349
rect 8159 1309 8171 1312
rect 8113 1303 8171 1309
rect 8289 1309 8301 1343
rect 8335 1309 8347 1343
rect 8404 1340 8432 1380
rect 8478 1368 8484 1420
rect 8536 1408 8542 1420
rect 9398 1408 9404 1420
rect 8536 1380 8800 1408
rect 9359 1380 9404 1408
rect 8536 1368 8542 1380
rect 8570 1340 8576 1352
rect 8404 1312 8576 1340
rect 8289 1303 8347 1309
rect 3418 1232 3424 1284
rect 3476 1272 3482 1284
rect 4157 1275 4215 1281
rect 4157 1272 4169 1275
rect 3476 1244 4169 1272
rect 3476 1232 3482 1244
rect 4157 1241 4169 1244
rect 4203 1272 4215 1275
rect 5258 1272 5264 1284
rect 4203 1244 5264 1272
rect 4203 1241 4215 1244
rect 4157 1235 4215 1241
rect 5258 1232 5264 1244
rect 5316 1232 5322 1284
rect 3786 1204 3792 1216
rect 3747 1176 3792 1204
rect 3786 1164 3792 1176
rect 3844 1164 3850 1216
rect 7926 1204 7932 1216
rect 7887 1176 7932 1204
rect 7926 1164 7932 1176
rect 7984 1204 7990 1216
rect 8312 1204 8340 1303
rect 8570 1300 8576 1312
rect 8628 1340 8634 1352
rect 8665 1343 8723 1349
rect 8665 1340 8677 1343
rect 8628 1312 8677 1340
rect 8628 1300 8634 1312
rect 8665 1309 8677 1312
rect 8711 1309 8723 1343
rect 8772 1340 8800 1380
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
rect 8941 1343 8999 1349
rect 8941 1340 8953 1343
rect 8772 1312 8953 1340
rect 8665 1303 8723 1309
rect 8941 1309 8953 1312
rect 8987 1309 8999 1343
rect 8941 1303 8999 1309
rect 7984 1176 8340 1204
rect 7984 1164 7990 1176
rect 8386 1164 8392 1216
rect 8444 1204 8450 1216
rect 8481 1207 8539 1213
rect 8481 1204 8493 1207
rect 8444 1176 8493 1204
rect 8444 1164 8450 1176
rect 8481 1173 8493 1176
rect 8527 1173 8539 1207
rect 8481 1167 8539 1173
rect 8662 1164 8668 1216
rect 8720 1204 8726 1216
rect 8849 1207 8907 1213
rect 8849 1204 8861 1207
rect 8720 1176 8861 1204
rect 8720 1164 8726 1176
rect 8849 1173 8861 1176
rect 8895 1173 8907 1207
rect 9214 1204 9220 1216
rect 9175 1176 9220 1204
rect 8849 1167 8907 1173
rect 9214 1164 9220 1176
rect 9272 1164 9278 1216
rect 3036 1114 9844 1136
rect 3036 1062 4116 1114
rect 4168 1062 4180 1114
rect 4232 1062 4244 1114
rect 4296 1062 4308 1114
rect 4360 1062 4372 1114
rect 4424 1062 7216 1114
rect 7268 1062 7280 1114
rect 7332 1062 7344 1114
rect 7396 1062 7408 1114
rect 7460 1062 7472 1114
rect 7524 1062 9844 1114
rect 3036 1040 9844 1062
rect 3786 960 3792 1012
rect 3844 1000 3850 1012
rect 10686 1000 10692 1012
rect 3844 972 10692 1000
rect 3844 960 3850 972
rect 10686 960 10692 972
rect 10744 960 10750 1012
rect 7926 892 7932 944
rect 7984 932 7990 944
rect 9674 932 9680 944
rect 7984 904 9680 932
rect 7984 892 7990 904
rect 9674 892 9680 904
rect 9732 892 9738 944
rect 8570 824 8576 876
rect 8628 864 8634 876
rect 16574 864 16580 876
rect 8628 836 16580 864
rect 8628 824 8634 836
rect 16574 824 16580 836
rect 16632 824 16638 876
<< via1 >>
rect 2412 11908 2464 11960
rect 8668 11908 8720 11960
rect 2964 11772 3016 11824
rect 8300 11772 8352 11824
rect 1492 11704 1544 11756
rect 6920 11704 6972 11756
rect 8392 11704 8444 11756
rect 10416 11704 10468 11756
rect 3424 11636 3476 11688
rect 6092 11636 6144 11688
rect 6184 11636 6236 11688
rect 16672 11636 16724 11688
rect 1308 11568 1360 11620
rect 6276 11568 6328 11620
rect 7380 11568 7432 11620
rect 9864 11568 9916 11620
rect 3516 11500 3568 11552
rect 7656 11500 7708 11552
rect 7748 11500 7800 11552
rect 9772 11500 9824 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 5858 11398 5910 11450
rect 5922 11398 5974 11450
rect 8766 11398 8818 11450
rect 8830 11398 8882 11450
rect 8894 11398 8946 11450
rect 8958 11398 9010 11450
rect 9022 11398 9074 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 2964 11296 3016 11348
rect 1308 11135 1360 11144
rect 1308 11101 1317 11135
rect 1317 11101 1351 11135
rect 1351 11101 1360 11135
rect 1308 11092 1360 11101
rect 3608 11228 3660 11280
rect 4620 11296 4672 11348
rect 5172 11296 5224 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 6184 11296 6236 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6552 11339 6604 11348
rect 6276 11296 6328 11305
rect 6552 11305 6561 11339
rect 6561 11305 6595 11339
rect 6595 11305 6604 11339
rect 6552 11296 6604 11305
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 8576 11296 8628 11348
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2412 11135 2464 11144
rect 2136 11092 2188 11101
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 3516 11160 3568 11212
rect 5540 11228 5592 11280
rect 6736 11228 6788 11280
rect 7748 11228 7800 11280
rect 8484 11228 8536 11280
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3424 11092 3476 11144
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 4620 11135 4672 11144
rect 940 11024 992 11076
rect 1860 11024 1912 11076
rect 1952 11024 2004 11076
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 2412 10956 2464 11008
rect 3516 10956 3568 11008
rect 4528 11024 4580 11076
rect 9496 11160 9548 11212
rect 5264 11092 5316 11144
rect 5632 11135 5684 11144
rect 5632 11101 5641 11135
rect 5641 11101 5675 11135
rect 5675 11101 5684 11135
rect 5632 11092 5684 11101
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6368 11092 6420 11144
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 7564 11135 7616 11144
rect 6828 11092 6880 11101
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8392 11092 8444 11144
rect 9128 11092 9180 11144
rect 9588 11092 9640 11144
rect 9220 11024 9272 11076
rect 3976 10956 4028 11008
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 5540 10956 5592 11008
rect 6828 10956 6880 11008
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 4116 10854 4168 10906
rect 4180 10854 4232 10906
rect 4244 10854 4296 10906
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 7216 10854 7268 10906
rect 7280 10854 7332 10906
rect 7344 10854 7396 10906
rect 7408 10854 7460 10906
rect 7472 10854 7524 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 1860 10752 1912 10804
rect 2136 10752 2188 10804
rect 2964 10752 3016 10804
rect 3056 10752 3108 10804
rect 1584 10684 1636 10736
rect 1124 10548 1176 10600
rect 1952 10616 2004 10668
rect 2136 10616 2188 10668
rect 2964 10616 3016 10668
rect 1400 10523 1452 10532
rect 1400 10489 1409 10523
rect 1409 10489 1443 10523
rect 1443 10489 1452 10523
rect 1400 10480 1452 10489
rect 1584 10480 1636 10532
rect 2228 10455 2280 10464
rect 2228 10421 2237 10455
rect 2237 10421 2271 10455
rect 2271 10421 2280 10455
rect 2228 10412 2280 10421
rect 3148 10480 3200 10532
rect 3424 10616 3476 10668
rect 3792 10616 3844 10668
rect 4712 10616 4764 10668
rect 5172 10659 5224 10668
rect 5172 10625 5181 10659
rect 5181 10625 5215 10659
rect 5215 10625 5224 10659
rect 5172 10616 5224 10625
rect 6920 10684 6972 10736
rect 6368 10616 6420 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 8668 10752 8720 10804
rect 8116 10684 8168 10736
rect 3792 10480 3844 10532
rect 4712 10480 4764 10532
rect 7840 10480 7892 10532
rect 8668 10548 8720 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 8116 10480 8168 10532
rect 3332 10412 3384 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 6184 10412 6236 10464
rect 8208 10412 8260 10464
rect 9588 10480 9640 10532
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 5858 10310 5910 10362
rect 5922 10310 5974 10362
rect 8766 10310 8818 10362
rect 8830 10310 8882 10362
rect 8894 10310 8946 10362
rect 8958 10310 9010 10362
rect 9022 10310 9074 10362
rect 15200 10276 15252 10328
rect 16580 10276 16632 10328
rect 1768 10208 1820 10260
rect 3424 10208 3476 10260
rect 2412 10072 2464 10124
rect 4712 10072 4764 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1584 10004 1636 10056
rect 1860 10004 1912 10056
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 5540 10047 5592 10056
rect 3424 10004 3476 10013
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 3700 9936 3752 9988
rect 1308 9911 1360 9920
rect 1308 9877 1317 9911
rect 1317 9877 1351 9911
rect 1351 9877 1360 9911
rect 1308 9868 1360 9877
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2228 9868 2280 9920
rect 4620 9868 4672 9920
rect 7840 10208 7892 10260
rect 8208 10208 8260 10260
rect 7472 10072 7524 10124
rect 7840 10115 7892 10124
rect 7840 10081 7849 10115
rect 7849 10081 7883 10115
rect 7883 10081 7892 10115
rect 7840 10072 7892 10081
rect 6092 10004 6144 10056
rect 6276 10004 6328 10056
rect 7932 10004 7984 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 7472 9936 7524 9988
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 4116 9766 4168 9818
rect 4180 9766 4232 9818
rect 4244 9766 4296 9818
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 7216 9766 7268 9818
rect 7280 9766 7332 9818
rect 7344 9766 7396 9818
rect 7408 9766 7460 9818
rect 7472 9766 7524 9818
rect 2136 9664 2188 9716
rect 1308 9639 1360 9648
rect 1308 9605 1317 9639
rect 1317 9605 1351 9639
rect 1351 9605 1360 9639
rect 1308 9596 1360 9605
rect 1032 9528 1084 9580
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 3700 9664 3752 9716
rect 6092 9664 6144 9716
rect 6552 9664 6604 9716
rect 3516 9596 3568 9648
rect 4896 9596 4948 9648
rect 5540 9596 5592 9648
rect 7748 9634 7800 9686
rect 8208 9664 8260 9716
rect 8300 9664 8352 9716
rect 21364 9664 21416 9716
rect 22100 9664 22152 9716
rect 1308 9460 1360 9512
rect 2964 9528 3016 9580
rect 4436 9528 4488 9580
rect 5908 9528 5960 9580
rect 6092 9528 6144 9580
rect 6276 9528 6328 9580
rect 3332 9460 3384 9512
rect 5724 9460 5776 9512
rect 1952 9324 2004 9376
rect 3608 9324 3660 9376
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 6828 9460 6880 9512
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 6092 9324 6144 9376
rect 7104 9324 7156 9376
rect 7656 9324 7708 9376
rect 8484 9324 8536 9376
rect 9404 9324 9456 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 5858 9222 5910 9274
rect 5922 9222 5974 9274
rect 8766 9222 8818 9274
rect 8830 9222 8882 9274
rect 8894 9222 8946 9274
rect 8958 9222 9010 9274
rect 9022 9222 9074 9274
rect 1492 9163 1544 9172
rect 1492 9129 1501 9163
rect 1501 9129 1535 9163
rect 1535 9129 1544 9163
rect 1492 9120 1544 9129
rect 2044 9120 2096 9172
rect 3516 9120 3568 9172
rect 3700 9120 3752 9172
rect 848 8916 900 8968
rect 4712 9120 4764 9172
rect 5264 9120 5316 9172
rect 9404 9163 9456 9172
rect 1676 8984 1728 9036
rect 4436 8984 4488 9036
rect 4712 8984 4764 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 3148 8916 3200 8968
rect 2504 8848 2556 8900
rect 2872 8848 2924 8900
rect 3608 8916 3660 8968
rect 6920 8984 6972 9036
rect 7840 8984 7892 9036
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 3700 8848 3752 8900
rect 3976 8848 4028 8900
rect 4896 8891 4948 8900
rect 4896 8857 4905 8891
rect 4905 8857 4939 8891
rect 4939 8857 4948 8891
rect 4896 8848 4948 8857
rect 5908 8848 5960 8900
rect 6092 8848 6144 8900
rect 7012 8848 7064 8900
rect 8484 8916 8536 8968
rect 9680 8848 9732 8900
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 5172 8780 5224 8832
rect 6644 8780 6696 8832
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 7840 8780 7892 8832
rect 8668 8780 8720 8832
rect 4116 8678 4168 8730
rect 4180 8678 4232 8730
rect 4244 8678 4296 8730
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 7216 8678 7268 8730
rect 7280 8678 7332 8730
rect 7344 8678 7396 8730
rect 7408 8678 7460 8730
rect 7472 8678 7524 8730
rect 1860 8576 1912 8628
rect 2320 8508 2372 8560
rect 3424 8576 3476 8628
rect 3516 8576 3568 8628
rect 5724 8576 5776 8628
rect 5908 8619 5960 8628
rect 5908 8585 5917 8619
rect 5917 8585 5951 8619
rect 5951 8585 5960 8619
rect 5908 8576 5960 8585
rect 7564 8576 7616 8628
rect 2872 8508 2924 8560
rect 4712 8508 4764 8560
rect 6828 8508 6880 8560
rect 9956 8576 10008 8628
rect 8024 8508 8076 8560
rect 1308 8483 1360 8492
rect 1308 8449 1317 8483
rect 1317 8449 1351 8483
rect 1351 8449 1360 8483
rect 1308 8440 1360 8449
rect 5908 8440 5960 8492
rect 6644 8440 6696 8492
rect 1768 8372 1820 8424
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 2596 8372 2648 8424
rect 3240 8372 3292 8424
rect 3608 8372 3660 8424
rect 4988 8372 5040 8424
rect 5724 8372 5776 8424
rect 9220 8440 9272 8492
rect 8668 8372 8720 8424
rect 1860 8304 1912 8356
rect 1952 8236 2004 8288
rect 3148 8236 3200 8288
rect 3976 8236 4028 8288
rect 6000 8236 6052 8288
rect 7012 8236 7064 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 5858 8134 5910 8186
rect 5922 8134 5974 8186
rect 8766 8134 8818 8186
rect 8830 8134 8882 8186
rect 8894 8134 8946 8186
rect 8958 8134 9010 8186
rect 9022 8134 9074 8186
rect 1676 8032 1728 8084
rect 3884 8032 3936 8084
rect 5172 8032 5224 8084
rect 7564 8032 7616 8084
rect 7840 8032 7892 8084
rect 8484 8032 8536 8084
rect 9220 8032 9272 8084
rect 9588 8032 9640 8084
rect 6552 7964 6604 8016
rect 8116 7964 8168 8016
rect 1584 7896 1636 7948
rect 6000 7896 6052 7948
rect 1492 7828 1544 7880
rect 1032 7760 1084 7812
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3148 7803 3200 7812
rect 3148 7769 3157 7803
rect 3157 7769 3191 7803
rect 3191 7769 3200 7803
rect 3148 7760 3200 7769
rect 5632 7828 5684 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7104 7828 7156 7880
rect 3884 7760 3936 7812
rect 6000 7760 6052 7812
rect 8484 7828 8536 7880
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 1584 7692 1636 7744
rect 1768 7692 1820 7744
rect 3424 7692 3476 7744
rect 3976 7692 4028 7744
rect 5356 7692 5408 7744
rect 6460 7692 6512 7744
rect 6552 7692 6604 7744
rect 7932 7692 7984 7744
rect 9496 7760 9548 7812
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 4116 7590 4168 7642
rect 4180 7590 4232 7642
rect 4244 7590 4296 7642
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 7216 7590 7268 7642
rect 7280 7590 7332 7642
rect 7344 7590 7396 7642
rect 7408 7590 7460 7642
rect 7472 7590 7524 7642
rect 10692 7624 10744 7676
rect 15200 7624 15252 7676
rect 11060 7556 11112 7608
rect 20628 7624 20680 7676
rect 2320 7420 2372 7472
rect 3240 7420 3292 7472
rect 5632 7463 5684 7472
rect 5632 7429 5641 7463
rect 5641 7429 5675 7463
rect 5675 7429 5684 7463
rect 5632 7420 5684 7429
rect 13820 7488 13872 7540
rect 1952 7352 2004 7404
rect 2044 7352 2096 7404
rect 4804 7352 4856 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 6920 7352 6972 7404
rect 6184 7284 6236 7336
rect 1768 7216 1820 7268
rect 2412 7216 2464 7268
rect 4528 7216 4580 7268
rect 4804 7216 4856 7268
rect 7196 7216 7248 7268
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 8300 7284 8352 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9312 7216 9364 7268
rect 756 7148 808 7200
rect 3240 7148 3292 7200
rect 8024 7148 8076 7200
rect 8116 7148 8168 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 5858 7046 5910 7098
rect 5922 7046 5974 7098
rect 8766 7046 8818 7098
rect 8830 7046 8882 7098
rect 8894 7046 8946 7098
rect 8958 7046 9010 7098
rect 9022 7046 9074 7098
rect 1308 6944 1360 6996
rect 1584 6944 1636 6996
rect 6552 6944 6604 6996
rect 7104 6944 7156 6996
rect 5724 6876 5776 6928
rect 6368 6876 6420 6928
rect 8300 6876 8352 6928
rect 2044 6808 2096 6860
rect 2044 6672 2096 6724
rect 1032 6604 1084 6656
rect 2596 6604 2648 6656
rect 2688 6604 2740 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4528 6808 4580 6860
rect 6828 6808 6880 6860
rect 8024 6808 8076 6860
rect 8484 6808 8536 6860
rect 9220 6808 9272 6860
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 4712 6672 4764 6724
rect 5908 6672 5960 6724
rect 5540 6604 5592 6656
rect 5632 6604 5684 6656
rect 7012 6672 7064 6724
rect 7196 6672 7248 6724
rect 8392 6672 8444 6724
rect 7564 6604 7616 6656
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 8852 6604 8904 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 4116 6502 4168 6554
rect 4180 6502 4232 6554
rect 4244 6502 4296 6554
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 7216 6502 7268 6554
rect 7280 6502 7332 6554
rect 7344 6502 7396 6554
rect 7408 6502 7460 6554
rect 7472 6502 7524 6554
rect 1308 6400 1360 6452
rect 2688 6375 2740 6384
rect 1308 6307 1360 6316
rect 1308 6273 1317 6307
rect 1317 6273 1351 6307
rect 1351 6273 1360 6307
rect 1308 6264 1360 6273
rect 2688 6341 2697 6375
rect 2697 6341 2731 6375
rect 2731 6341 2740 6375
rect 2688 6332 2740 6341
rect 2780 6332 2832 6384
rect 3148 6332 3200 6384
rect 4528 6400 4580 6452
rect 6000 6400 6052 6452
rect 7748 6400 7800 6452
rect 4712 6332 4764 6384
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3976 6264 4028 6316
rect 4436 6264 4488 6316
rect 5908 6332 5960 6384
rect 8116 6332 8168 6384
rect 8576 6332 8628 6384
rect 6000 6307 6052 6316
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 4988 6196 5040 6248
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6276 6264 6328 6316
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 7840 6196 7892 6248
rect 1952 6060 2004 6112
rect 8852 6128 8904 6180
rect 3976 6060 4028 6112
rect 4804 6060 4856 6112
rect 6184 6060 6236 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 7104 6060 7156 6112
rect 9312 6060 9364 6112
rect 16672 6060 16724 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 5858 5958 5910 6010
rect 5922 5958 5974 6010
rect 8766 5958 8818 6010
rect 8830 5958 8882 6010
rect 8894 5958 8946 6010
rect 8958 5958 9010 6010
rect 9022 5958 9074 6010
rect 1400 5856 1452 5908
rect 1860 5856 1912 5908
rect 2320 5856 2372 5908
rect 1584 5831 1636 5840
rect 1584 5797 1593 5831
rect 1593 5797 1627 5831
rect 1627 5797 1636 5831
rect 1584 5788 1636 5797
rect 2136 5788 2188 5840
rect 1492 5652 1544 5704
rect 1952 5652 2004 5704
rect 3424 5856 3476 5908
rect 6368 5899 6420 5908
rect 3148 5788 3200 5840
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 7012 5856 7064 5908
rect 8576 5856 8628 5908
rect 8668 5856 8720 5908
rect 3608 5720 3660 5772
rect 5632 5788 5684 5840
rect 6644 5788 6696 5840
rect 5172 5720 5224 5772
rect 5540 5720 5592 5772
rect 2964 5652 3016 5704
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 6276 5695 6328 5704
rect 1216 5584 1268 5636
rect 1860 5516 1912 5568
rect 3516 5584 3568 5636
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6552 5720 6604 5772
rect 6920 5720 6972 5772
rect 7196 5652 7248 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 2596 5559 2648 5568
rect 2596 5525 2605 5559
rect 2605 5525 2639 5559
rect 2639 5525 2648 5559
rect 2596 5516 2648 5525
rect 2872 5516 2924 5568
rect 4436 5584 4488 5636
rect 5172 5584 5224 5636
rect 6368 5584 6420 5636
rect 8300 5627 8352 5636
rect 6460 5516 6512 5568
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 8300 5593 8309 5627
rect 8309 5593 8343 5627
rect 8343 5593 8352 5627
rect 8300 5584 8352 5593
rect 6828 5516 6880 5525
rect 9864 5516 9916 5568
rect 4116 5414 4168 5466
rect 4180 5414 4232 5466
rect 4244 5414 4296 5466
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 7216 5414 7268 5466
rect 7280 5414 7332 5466
rect 7344 5414 7396 5466
rect 7408 5414 7460 5466
rect 7472 5414 7524 5466
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 8116 5312 8168 5364
rect 9956 5312 10008 5364
rect 1124 5244 1176 5296
rect 2504 5244 2556 5296
rect 2412 5176 2464 5228
rect 3608 5244 3660 5296
rect 6644 5244 6696 5296
rect 7748 5244 7800 5296
rect 5264 5219 5316 5228
rect 3056 5108 3108 5160
rect 4988 5108 5040 5160
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 7104 5176 7156 5228
rect 2320 5040 2372 5092
rect 3332 5040 3384 5092
rect 3148 4972 3200 5024
rect 3424 4972 3476 5024
rect 3608 4972 3660 5024
rect 4896 4972 4948 5024
rect 4988 4972 5040 5024
rect 5172 5108 5224 5160
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 8484 5176 8536 5228
rect 8392 5108 8444 5160
rect 6092 4972 6144 5024
rect 9588 4972 9640 5024
rect 16580 4972 16632 5024
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 5858 4870 5910 4922
rect 5922 4870 5974 4922
rect 8766 4870 8818 4922
rect 8830 4870 8882 4922
rect 8894 4870 8946 4922
rect 8958 4870 9010 4922
rect 9022 4870 9074 4922
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 4712 4768 4764 4820
rect 8208 4768 8260 4820
rect 8668 4768 8720 4820
rect 9220 4768 9272 4820
rect 2780 4700 2832 4752
rect 3148 4700 3200 4752
rect 1676 4564 1728 4616
rect 2780 4564 2832 4616
rect 2964 4564 3016 4616
rect 5172 4700 5224 4752
rect 4804 4632 4856 4684
rect 4988 4632 5040 4684
rect 1032 4496 1084 4548
rect 4068 4564 4120 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 4528 4496 4580 4548
rect 8576 4700 8628 4752
rect 6552 4632 6604 4684
rect 8024 4632 8076 4684
rect 8208 4632 8260 4684
rect 9220 4632 9272 4684
rect 9772 4564 9824 4616
rect 2964 4428 3016 4480
rect 3332 4428 3384 4480
rect 6552 4539 6604 4548
rect 6552 4505 6561 4539
rect 6561 4505 6595 4539
rect 6595 4505 6604 4539
rect 6552 4496 6604 4505
rect 4988 4428 5040 4480
rect 5540 4428 5592 4480
rect 6368 4428 6420 4480
rect 6460 4428 6512 4480
rect 8852 4496 8904 4548
rect 7932 4428 7984 4480
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8944 4471 8996 4480
rect 8116 4428 8168 4437
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 4116 4326 4168 4378
rect 4180 4326 4232 4378
rect 4244 4326 4296 4378
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 7216 4326 7268 4378
rect 7280 4326 7332 4378
rect 7344 4326 7396 4378
rect 7408 4326 7460 4378
rect 7472 4326 7524 4378
rect 6736 4224 6788 4276
rect 8116 4224 8168 4276
rect 8944 4224 8996 4276
rect 4436 4156 4488 4208
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3884 4088 3936 4140
rect 4896 4088 4948 4140
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6552 4088 6604 4140
rect 7748 4156 7800 4208
rect 7932 4156 7984 4208
rect 8576 4131 8628 4140
rect 6276 4020 6328 4072
rect 7196 4020 7248 4072
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 8668 4088 8720 4140
rect 7932 4020 7984 4072
rect 8852 4020 8904 4072
rect 9496 4020 9548 4072
rect 5632 3952 5684 4004
rect 9036 3952 9088 4004
rect 10048 3952 10100 4004
rect 3332 3884 3384 3936
rect 3608 3884 3660 3936
rect 4160 3884 4212 3936
rect 6460 3884 6512 3936
rect 6920 3884 6972 3936
rect 16580 3884 16632 3936
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 5858 3782 5910 3834
rect 5922 3782 5974 3834
rect 8766 3782 8818 3834
rect 8830 3782 8882 3834
rect 8894 3782 8946 3834
rect 8958 3782 9010 3834
rect 9022 3782 9074 3834
rect 3056 3680 3108 3732
rect 4252 3680 4304 3732
rect 4436 3680 4488 3732
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 3240 3476 3292 3528
rect 3608 3612 3660 3664
rect 4068 3655 4120 3664
rect 4068 3621 4077 3655
rect 4077 3621 4111 3655
rect 4111 3621 4120 3655
rect 4068 3612 4120 3621
rect 6552 3680 6604 3732
rect 8576 3680 8628 3732
rect 3792 3476 3844 3528
rect 5908 3612 5960 3664
rect 8208 3612 8260 3664
rect 8760 3612 8812 3664
rect 4804 3544 4856 3596
rect 6920 3587 6972 3596
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 8576 3544 8628 3596
rect 9312 3680 9364 3732
rect 5540 3476 5592 3528
rect 6552 3519 6604 3528
rect 5080 3408 5132 3460
rect 5632 3408 5684 3460
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 7840 3476 7892 3528
rect 8484 3476 8536 3528
rect 8208 3408 8260 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 8484 3340 8536 3392
rect 8668 3340 8720 3392
rect 9312 3340 9364 3392
rect 4116 3238 4168 3290
rect 4180 3238 4232 3290
rect 4244 3238 4296 3290
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 7216 3238 7268 3290
rect 7280 3238 7332 3290
rect 7344 3238 7396 3290
rect 7408 3238 7460 3290
rect 7472 3238 7524 3290
rect 3792 3136 3844 3188
rect 5724 3068 5776 3120
rect 5908 3068 5960 3120
rect 7288 3068 7340 3120
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4160 3000 4212 3052
rect 4436 3000 4488 3052
rect 6184 3000 6236 3052
rect 6828 3000 6880 3052
rect 9036 3136 9088 3188
rect 2688 2864 2740 2916
rect 3608 2864 3660 2916
rect 3884 2864 3936 2916
rect 3976 2864 4028 2916
rect 4988 2932 5040 2984
rect 4344 2796 4396 2848
rect 4804 2796 4856 2848
rect 4896 2796 4948 2848
rect 5264 2796 5316 2848
rect 6276 2864 6328 2916
rect 6644 2796 6696 2848
rect 7196 2932 7248 2984
rect 7656 2932 7708 2984
rect 7012 2864 7064 2916
rect 7564 2864 7616 2916
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8944 3068 8996 3120
rect 8852 3000 8904 3052
rect 9036 3000 9088 3052
rect 9220 3000 9272 3052
rect 8668 2932 8720 2984
rect 8116 2796 8168 2848
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 5858 2694 5910 2746
rect 5922 2694 5974 2746
rect 8766 2694 8818 2746
rect 8830 2694 8882 2746
rect 8894 2694 8946 2746
rect 8958 2694 9010 2746
rect 9022 2694 9074 2746
rect 3424 2592 3476 2644
rect 3608 2592 3660 2644
rect 4068 2635 4120 2644
rect 4068 2601 4077 2635
rect 4077 2601 4111 2635
rect 4111 2601 4120 2635
rect 4068 2592 4120 2601
rect 4896 2592 4948 2644
rect 5172 2592 5224 2644
rect 6000 2592 6052 2644
rect 6552 2592 6604 2644
rect 7104 2592 7156 2644
rect 7564 2592 7616 2644
rect 3332 2524 3384 2576
rect 4344 2524 4396 2576
rect 4712 2524 4764 2576
rect 5264 2524 5316 2576
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 6184 2567 6236 2576
rect 6184 2533 6193 2567
rect 6193 2533 6227 2567
rect 6227 2533 6236 2567
rect 6184 2524 6236 2533
rect 6460 2524 6512 2576
rect 2688 2456 2740 2508
rect 3792 2456 3844 2508
rect 4436 2456 4488 2508
rect 3424 2388 3476 2440
rect 2964 2252 3016 2304
rect 3608 2252 3660 2304
rect 4068 2320 4120 2372
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5724 2320 5776 2372
rect 4988 2252 5040 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 5264 2252 5316 2304
rect 5540 2252 5592 2304
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 6092 2252 6144 2304
rect 6736 2320 6788 2372
rect 7656 2320 7708 2372
rect 8024 2456 8076 2508
rect 9220 2592 9272 2644
rect 21364 2592 21416 2644
rect 8300 2431 8352 2440
rect 7012 2252 7064 2304
rect 7748 2252 7800 2304
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8024 2320 8076 2372
rect 9128 2456 9180 2508
rect 8668 2388 8720 2440
rect 9772 2388 9824 2440
rect 8944 2320 8996 2372
rect 16580 2320 16632 2372
rect 9220 2252 9272 2304
rect 16672 2252 16724 2304
rect 4116 2150 4168 2202
rect 4180 2150 4232 2202
rect 4244 2150 4296 2202
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 7216 2150 7268 2202
rect 7280 2150 7332 2202
rect 7344 2150 7396 2202
rect 7408 2150 7460 2202
rect 7472 2150 7524 2202
rect 3148 2048 3200 2100
rect 3792 2091 3844 2100
rect 3792 2057 3801 2091
rect 3801 2057 3835 2091
rect 3835 2057 3844 2091
rect 3792 2048 3844 2057
rect 4620 2048 4672 2100
rect 4712 1980 4764 2032
rect 2688 1912 2740 1964
rect 3608 1955 3660 1964
rect 3608 1921 3617 1955
rect 3617 1921 3651 1955
rect 3651 1921 3660 1955
rect 3608 1912 3660 1921
rect 4068 1955 4120 1964
rect 4068 1921 4077 1955
rect 4077 1921 4111 1955
rect 4111 1921 4120 1955
rect 4068 1912 4120 1921
rect 4528 1912 4580 1964
rect 4252 1844 4304 1896
rect 4804 1844 4856 1896
rect 3700 1776 3752 1828
rect 3976 1776 4028 1828
rect 5356 2048 5408 2100
rect 7104 2048 7156 2100
rect 7840 2091 7892 2100
rect 7840 2057 7849 2091
rect 7849 2057 7883 2091
rect 7883 2057 7892 2091
rect 7840 2048 7892 2057
rect 7932 2048 7984 2100
rect 8208 2048 8260 2100
rect 9036 2048 9088 2100
rect 9404 2091 9456 2100
rect 9404 2057 9413 2091
rect 9413 2057 9447 2091
rect 9447 2057 9456 2091
rect 9404 2048 9456 2057
rect 4988 1980 5040 2032
rect 5448 1980 5500 2032
rect 5540 1980 5592 2032
rect 6736 1980 6788 2032
rect 7564 1980 7616 2032
rect 6920 1912 6972 1964
rect 7656 1955 7708 1964
rect 7656 1921 7665 1955
rect 7665 1921 7699 1955
rect 7699 1921 7708 1955
rect 7656 1912 7708 1921
rect 8024 1912 8076 1964
rect 8484 1955 8536 1964
rect 8484 1921 8493 1955
rect 8493 1921 8527 1955
rect 8527 1921 8536 1955
rect 8484 1912 8536 1921
rect 9312 1980 9364 2032
rect 5080 1844 5132 1896
rect 6736 1844 6788 1896
rect 9496 1776 9548 1828
rect 3608 1708 3660 1760
rect 5264 1708 5316 1760
rect 5666 1606 5718 1658
rect 5730 1606 5782 1658
rect 5794 1606 5846 1658
rect 5858 1606 5910 1658
rect 5922 1606 5974 1658
rect 8766 1606 8818 1658
rect 8830 1606 8882 1658
rect 8894 1606 8946 1658
rect 8958 1606 9010 1658
rect 9022 1606 9074 1658
rect 5172 1504 5224 1556
rect 2872 1436 2924 1488
rect 4068 1436 4120 1488
rect 8116 1504 8168 1556
rect 10968 1436 11020 1488
rect 3516 1300 3568 1352
rect 3608 1343 3660 1352
rect 3608 1309 3617 1343
rect 3617 1309 3651 1343
rect 3651 1309 3660 1343
rect 3884 1343 3936 1352
rect 3608 1300 3660 1309
rect 3884 1309 3893 1343
rect 3893 1309 3927 1343
rect 3927 1309 3936 1343
rect 3884 1300 3936 1309
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 8484 1368 8536 1420
rect 9404 1411 9456 1420
rect 3424 1232 3476 1284
rect 5264 1232 5316 1284
rect 3792 1207 3844 1216
rect 3792 1173 3801 1207
rect 3801 1173 3835 1207
rect 3835 1173 3844 1207
rect 3792 1164 3844 1173
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 8576 1300 8628 1352
rect 9404 1377 9413 1411
rect 9413 1377 9447 1411
rect 9447 1377 9456 1411
rect 9404 1368 9456 1377
rect 7932 1164 7984 1173
rect 8392 1164 8444 1216
rect 8668 1164 8720 1216
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 4116 1062 4168 1114
rect 4180 1062 4232 1114
rect 4244 1062 4296 1114
rect 4308 1062 4360 1114
rect 4372 1062 4424 1114
rect 7216 1062 7268 1114
rect 7280 1062 7332 1114
rect 7344 1062 7396 1114
rect 7408 1062 7460 1114
rect 7472 1062 7524 1114
rect 3792 960 3844 1012
rect 10692 960 10744 1012
rect 7932 892 7984 944
rect 9680 892 9732 944
rect 8576 824 8628 876
rect 16580 824 16632 876
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 22098 12336 22154 12345
rect 22098 12271 22154 12280
rect 952 11234 980 12200
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 768 11206 980 11234
rect 768 7206 796 11206
rect 1320 11150 1348 11562
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 940 11076 992 11082
rect 940 11018 992 11024
rect 846 9616 902 9625
rect 846 9551 902 9560
rect 860 8974 888 9551
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 756 7200 808 7206
rect 756 7142 808 7148
rect 952 5534 980 11018
rect 1412 10690 1440 12200
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11354 1532 11698
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1872 11082 1900 12200
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1768 11008 1820 11014
rect 1766 10976 1768 10985
rect 1820 10976 1822 10985
rect 1766 10911 1822 10920
rect 1858 10840 1914 10849
rect 1676 10804 1728 10810
rect 1858 10775 1860 10784
rect 1676 10746 1728 10752
rect 1912 10775 1914 10784
rect 1860 10746 1912 10752
rect 1228 10662 1440 10690
rect 1584 10736 1636 10742
rect 1688 10713 1716 10746
rect 1584 10678 1636 10684
rect 1674 10704 1730 10713
rect 1124 10600 1176 10606
rect 1124 10542 1176 10548
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 1044 8537 1072 9522
rect 1030 8528 1086 8537
rect 1030 8463 1086 8472
rect 1032 7812 1084 7818
rect 1032 7754 1084 7760
rect 1044 6662 1072 7754
rect 1032 6656 1084 6662
rect 1032 6598 1084 6604
rect 952 5506 1072 5534
rect 1044 4554 1072 5506
rect 1136 5302 1164 10542
rect 1228 5642 1256 10662
rect 1398 10568 1454 10577
rect 1596 10538 1624 10678
rect 1964 10674 1992 11018
rect 1674 10639 1730 10648
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1398 10503 1400 10512
rect 1452 10503 1454 10512
rect 1584 10532 1636 10538
rect 1400 10474 1452 10480
rect 1584 10474 1636 10480
rect 1596 10062 1624 10474
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1308 9920 1360 9926
rect 1308 9862 1360 9868
rect 1320 9654 1348 9862
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1320 8498 1348 9454
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1320 7002 1348 8434
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1320 6458 1348 6938
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6225 1348 6258
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1412 5914 1440 9998
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1490 9480 1546 9489
rect 1490 9415 1546 9424
rect 1504 9178 1532 9415
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1490 8800 1546 8809
rect 1490 8735 1546 8744
rect 1504 7886 1532 8735
rect 1596 7954 1624 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1688 9042 1716 9522
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8090 1716 8978
rect 1780 8514 1808 10202
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9081 1900 9998
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1858 9072 1914 9081
rect 1858 9007 1914 9016
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8634 1900 8910
rect 1964 8673 1992 9318
rect 2056 9178 2084 11086
rect 2148 10810 2176 11086
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 9722 2176 10610
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 9926 2268 10406
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2134 9072 2190 9081
rect 2134 9007 2190 9016
rect 2148 8974 2176 9007
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1950 8664 2006 8673
rect 1860 8628 1912 8634
rect 1950 8599 2006 8608
rect 1860 8570 1912 8576
rect 1780 8486 1900 8514
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1504 5710 1532 7686
rect 1596 7002 1624 7686
rect 1688 7562 1716 8026
rect 1780 7750 1808 8366
rect 1872 8362 1900 8486
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1688 7534 1900 7562
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 5846 1624 6831
rect 1584 5840 1636 5846
rect 1584 5782 1636 5788
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1216 5636 1268 5642
rect 1216 5578 1268 5584
rect 1780 5534 1808 7210
rect 1872 5914 1900 7534
rect 1964 7410 1992 8230
rect 2056 7410 2084 8774
rect 2332 8650 2360 12200
rect 2412 11960 2464 11966
rect 2412 11902 2464 11908
rect 2792 11914 2820 12200
rect 2424 11150 2452 11902
rect 2792 11886 3188 11914
rect 2964 11824 3016 11830
rect 2964 11766 3016 11772
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2976 11354 3004 11766
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10130 2452 10950
rect 2976 10810 3004 11086
rect 3054 10840 3110 10849
rect 2964 10804 3016 10810
rect 3054 10775 3056 10784
rect 2964 10746 3016 10752
rect 3108 10775 3110 10784
rect 3056 10746 3108 10752
rect 3160 10690 3188 11886
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 3068 10662 3188 10690
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2870 10160 2926 10169
rect 2412 10124 2464 10130
rect 2870 10095 2926 10104
rect 2412 10066 2464 10072
rect 2410 10024 2466 10033
rect 2410 9959 2466 9968
rect 2240 8622 2360 8650
rect 2134 7984 2190 7993
rect 2134 7919 2190 7928
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6730 2084 6802
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1872 5817 1900 5850
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1964 5710 1992 6054
rect 2148 5846 2176 7919
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1688 5506 1808 5534
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 2240 5534 2268 8622
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2332 8430 2360 8502
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 7478 2360 8366
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2332 6474 2360 7414
rect 2424 7274 2452 9959
rect 2884 9466 2912 10095
rect 2976 9586 3004 10610
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2884 9438 3004 9466
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2596 8968 2648 8974
rect 2594 8936 2596 8945
rect 2648 8936 2650 8945
rect 2504 8900 2556 8906
rect 2594 8871 2650 8880
rect 2872 8900 2924 8906
rect 2504 8842 2556 8848
rect 2872 8842 2924 8848
rect 2516 8412 2544 8842
rect 2884 8809 2912 8842
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 2884 8566 2912 8735
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2596 8424 2648 8430
rect 2516 8384 2596 8412
rect 2596 8366 2648 8372
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2608 6718 2820 6746
rect 2608 6662 2636 6718
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2332 6446 2452 6474
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5914 2360 6258
rect 2424 6254 2452 6446
rect 2700 6390 2728 6598
rect 2792 6390 2820 6718
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1124 5296 1176 5302
rect 1124 5238 1176 5244
rect 1688 4622 1716 5506
rect 1872 4978 1900 5510
rect 2240 5506 2360 5534
rect 2332 5098 2360 5506
rect 2424 5234 2452 6190
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2976 5828 3004 9438
rect 2792 5800 3004 5828
rect 2686 5672 2742 5681
rect 2686 5607 2742 5616
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 1872 4950 2360 4978
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1032 4548 1084 4554
rect 1032 4490 1084 4496
rect 2332 1986 2360 4950
rect 2516 2417 2544 5238
rect 2608 5137 2636 5510
rect 2594 5128 2650 5137
rect 2594 5063 2650 5072
rect 2594 4720 2650 4729
rect 2594 4655 2650 4664
rect 2608 2496 2636 4655
rect 2700 2922 2728 5607
rect 2792 4758 2820 5800
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2792 3233 2820 4558
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2688 2508 2740 2514
rect 2608 2468 2688 2496
rect 2688 2450 2740 2456
rect 2502 2408 2558 2417
rect 2502 2343 2558 2352
rect 2332 1970 2728 1986
rect 2332 1964 2740 1970
rect 2332 1958 2688 1964
rect 2688 1906 2740 1912
rect 2884 1494 2912 5510
rect 2976 4622 3004 5646
rect 3068 5534 3096 10662
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 8974 3188 10474
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3252 8922 3280 12200
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3436 11150 3464 11630
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 3608 11280 3660 11286
rect 3606 11248 3608 11257
rect 3660 11248 3662 11257
rect 3516 11212 3568 11218
rect 3606 11183 3662 11192
rect 3516 11154 3568 11160
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 9518 3372 10406
rect 3436 10266 3464 10610
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3528 10169 3556 10950
rect 3514 10160 3570 10169
rect 3514 10095 3570 10104
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3252 8894 3372 8922
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7818 3188 8230
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3252 7478 3280 8366
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3160 5846 3188 6326
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3068 5506 3188 5534
rect 3054 5264 3110 5273
rect 3054 5199 3110 5208
rect 3068 5166 3096 5199
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3160 5030 3188 5506
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3054 4584 3110 4593
rect 3054 4519 3110 4528
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 2310 3004 4422
rect 3068 3738 3096 4519
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 3160 2106 3188 4694
rect 3252 3534 3280 7142
rect 3344 5098 3372 8894
rect 3436 8634 3464 9998
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3528 9178 3556 9590
rect 3620 9382 3648 11086
rect 3712 10146 3740 12200
rect 4172 11098 4200 12200
rect 4632 11506 4660 12200
rect 4632 11478 5028 11506
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4632 11150 4660 11290
rect 3896 11070 4200 11098
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4528 11076 4580 11082
rect 3790 10976 3846 10985
rect 3790 10911 3846 10920
rect 3804 10674 3832 10911
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3804 10305 3832 10474
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3712 10118 3832 10146
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3712 9722 3740 9930
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3712 9058 3740 9114
rect 3620 9030 3740 9058
rect 3620 8974 3648 9030
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3514 8664 3570 8673
rect 3424 8628 3476 8634
rect 3514 8599 3516 8608
rect 3424 8570 3476 8576
rect 3568 8599 3570 8608
rect 3516 8570 3568 8576
rect 3436 8412 3464 8570
rect 3608 8424 3660 8430
rect 3436 8384 3608 8412
rect 3436 7886 3464 8384
rect 3608 8366 3660 8372
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 6662 3464 7686
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3436 5914 3464 6151
rect 3620 5930 3648 6734
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3528 5902 3648 5930
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3436 5710 3464 5743
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3528 5642 3556 5902
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3620 5302 3648 5714
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3424 5024 3476 5030
rect 3330 4992 3386 5001
rect 3608 5024 3660 5030
rect 3476 4984 3556 5012
rect 3424 4966 3476 4972
rect 3330 4927 3386 4936
rect 3344 4570 3372 4927
rect 3344 4542 3464 4570
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4146 3372 4422
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3344 3058 3372 3878
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3344 2582 3372 2994
rect 3436 2650 3464 4542
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 2872 1488 2924 1494
rect 2872 1430 2924 1436
rect 3436 1290 3464 2382
rect 3528 1358 3556 4984
rect 3608 4966 3660 4972
rect 3620 3942 3648 4966
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3620 2922 3648 3606
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3606 2816 3662 2825
rect 3606 2751 3662 2760
rect 3620 2650 3648 2751
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3620 1970 3648 2246
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3620 1766 3648 1906
rect 3712 1834 3740 8842
rect 3804 3534 3832 10118
rect 3896 8090 3924 11070
rect 4528 11018 4580 11024
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 9625 4016 10950
rect 4116 10908 4424 10928
rect 4116 10906 4122 10908
rect 4178 10906 4202 10908
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4424 10908
rect 4178 10854 4180 10906
rect 4360 10854 4362 10906
rect 4116 10852 4122 10854
rect 4178 10852 4202 10854
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4424 10854
rect 4116 10832 4424 10852
rect 4116 9820 4424 9840
rect 4116 9818 4122 9820
rect 4178 9818 4202 9820
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4424 9820
rect 4178 9766 4180 9818
rect 4360 9766 4362 9818
rect 4116 9764 4122 9766
rect 4178 9764 4202 9766
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4424 9766
rect 4116 9744 4424 9764
rect 3974 9616 4030 9625
rect 3974 9551 4030 9560
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4448 9042 4476 9522
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3988 8294 4016 8842
rect 4116 8732 4424 8752
rect 4116 8730 4122 8732
rect 4178 8730 4202 8732
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4424 8732
rect 4178 8678 4180 8730
rect 4360 8678 4362 8730
rect 4116 8676 4122 8678
rect 4178 8676 4202 8678
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4424 8678
rect 4116 8656 4424 8676
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 4146 3924 7754
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 6322 4016 7686
rect 4116 7644 4424 7664
rect 4116 7642 4122 7644
rect 4178 7642 4202 7644
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4424 7644
rect 4178 7590 4180 7642
rect 4360 7590 4362 7642
rect 4116 7588 4122 7590
rect 4178 7588 4202 7590
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4424 7590
rect 4116 7568 4424 7588
rect 4540 7274 4568 11018
rect 4896 11008 4948 11014
rect 4816 10968 4896 10996
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 10538 4752 10610
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4116 6556 4424 6576
rect 4116 6554 4122 6556
rect 4178 6554 4202 6556
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4424 6556
rect 4178 6502 4180 6554
rect 4360 6502 4362 6554
rect 4116 6500 4122 6502
rect 4178 6500 4202 6502
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4424 6502
rect 4116 6480 4424 6500
rect 4540 6458 4568 6802
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 4729 4016 6054
rect 4448 5642 4476 6258
rect 4526 6216 4582 6225
rect 4526 6151 4582 6160
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4116 5468 4424 5488
rect 4116 5466 4122 5468
rect 4178 5466 4202 5468
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4424 5468
rect 4178 5414 4180 5466
rect 4360 5414 4362 5466
rect 4116 5412 4122 5414
rect 4178 5412 4202 5414
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4424 5414
rect 4116 5392 4424 5412
rect 4540 4978 4568 6151
rect 4448 4950 4568 4978
rect 3974 4720 4030 4729
rect 3974 4655 4030 4664
rect 4068 4616 4120 4622
rect 4448 4593 4476 4950
rect 4526 4856 4582 4865
rect 4526 4791 4528 4800
rect 4580 4791 4582 4800
rect 4528 4762 4580 4768
rect 4068 4558 4120 4564
rect 4434 4584 4490 4593
rect 4080 4468 4108 4558
rect 4434 4519 4490 4528
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 3988 4440 4108 4468
rect 3988 4264 4016 4440
rect 4116 4380 4424 4400
rect 4116 4378 4122 4380
rect 4178 4378 4202 4380
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4424 4380
rect 4178 4326 4180 4378
rect 4360 4326 4362 4378
rect 4116 4324 4122 4326
rect 4178 4324 4202 4326
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4424 4326
rect 4116 4304 4424 4324
rect 3988 4236 4292 4264
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3790 3360 3846 3369
rect 3790 3295 3846 3304
rect 3804 3194 3832 3295
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3896 3058 3924 3975
rect 4160 3936 4212 3942
rect 4080 3884 4160 3890
rect 4080 3878 4212 3884
rect 4080 3862 4200 3878
rect 4080 3670 4108 3862
rect 4264 3738 4292 4236
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3738 4476 4150
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4116 3292 4424 3312
rect 4116 3290 4122 3292
rect 4178 3290 4202 3292
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4424 3292
rect 4178 3238 4180 3290
rect 4360 3238 4362 3290
rect 4116 3236 4122 3238
rect 4178 3236 4202 3238
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4424 3238
rect 3974 3224 4030 3233
rect 4116 3216 4424 3236
rect 4540 3176 4568 4490
rect 3974 3159 4030 3168
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3988 2922 4016 3159
rect 4448 3148 4568 3176
rect 4066 3088 4122 3097
rect 4448 3058 4476 3148
rect 4632 3074 4660 9862
rect 4724 9178 4752 10066
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4724 8673 4752 8978
rect 4710 8664 4766 8673
rect 4710 8599 4766 8608
rect 4724 8566 4752 8599
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4816 7410 4844 10968
rect 4896 10950 4948 10956
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4908 9489 4936 9590
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4908 8809 4936 8842
rect 4894 8800 4950 8809
rect 4894 8735 4950 8744
rect 5000 8650 5028 11478
rect 4908 8622 5028 8650
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4724 6390 4752 6666
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4816 6118 4844 7210
rect 4804 6112 4856 6118
rect 4710 6080 4766 6089
rect 4804 6054 4856 6060
rect 4710 6015 4766 6024
rect 4724 5001 4752 6015
rect 4802 5944 4858 5953
rect 4802 5879 4858 5888
rect 4710 4992 4766 5001
rect 4710 4927 4766 4936
rect 4816 4842 4844 5879
rect 4908 5030 4936 8622
rect 4988 8424 5040 8430
rect 5092 8412 5120 12200
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5460 11354 5488 11591
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5184 10985 5212 11290
rect 5552 11286 5580 12200
rect 5666 11452 5974 11472
rect 5666 11450 5672 11452
rect 5728 11450 5752 11452
rect 5808 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5974 11452
rect 5728 11398 5730 11450
rect 5910 11398 5912 11450
rect 5666 11396 5672 11398
rect 5728 11396 5752 11398
rect 5808 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5974 11398
rect 5666 11376 5974 11396
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5264 11144 5316 11150
rect 5632 11144 5684 11150
rect 5264 11086 5316 11092
rect 5630 11112 5632 11121
rect 5724 11144 5776 11150
rect 5684 11112 5686 11121
rect 5170 10976 5226 10985
rect 5170 10911 5226 10920
rect 5184 10674 5212 10911
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5276 9466 5304 11086
rect 5724 11086 5776 11092
rect 5630 11047 5686 11056
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10577 5580 10950
rect 5736 10713 5764 11086
rect 5722 10704 5778 10713
rect 5722 10639 5778 10648
rect 5538 10568 5594 10577
rect 5538 10503 5594 10512
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5184 9438 5304 9466
rect 5184 8838 5212 9438
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9178 5304 9318
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5368 9081 5396 10406
rect 5666 10364 5974 10384
rect 5666 10362 5672 10364
rect 5728 10362 5752 10364
rect 5808 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5974 10364
rect 5728 10310 5730 10362
rect 5910 10310 5912 10362
rect 5666 10308 5672 10310
rect 5728 10308 5752 10310
rect 5808 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5974 10310
rect 5666 10288 5974 10308
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9654 5580 9998
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5722 9616 5778 9625
rect 5722 9551 5778 9560
rect 5908 9580 5960 9586
rect 5736 9518 5764 9551
rect 5908 9522 5960 9528
rect 5724 9512 5776 9518
rect 5920 9489 5948 9522
rect 5724 9454 5776 9460
rect 5906 9480 5962 9489
rect 5906 9415 5962 9424
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5354 9072 5410 9081
rect 5354 9007 5410 9016
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5092 8384 5304 8412
rect 4988 8366 5040 8372
rect 5000 7562 5028 8366
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5000 7534 5120 7562
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5000 6254 5028 7346
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5166 5028 6190
rect 5092 5370 5120 7534
rect 5184 5953 5212 8026
rect 5170 5944 5226 5953
rect 5170 5879 5226 5888
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5642 5212 5714
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 4865 5028 4966
rect 4986 4856 5042 4865
rect 4712 4820 4764 4826
rect 4816 4814 4936 4842
rect 4712 4762 4764 4768
rect 4066 3023 4122 3032
rect 4160 3052 4212 3058
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3804 2106 3832 2450
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3700 1828 3752 1834
rect 3700 1770 3752 1776
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3606 1456 3662 1465
rect 3606 1391 3662 1400
rect 3620 1358 3648 1391
rect 3896 1358 3924 2858
rect 4080 2650 4108 3023
rect 4160 2994 4212 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4540 3046 4660 3074
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4172 2553 4200 2994
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2582 4384 2790
rect 4344 2576 4396 2582
rect 4158 2544 4214 2553
rect 4344 2518 4396 2524
rect 4448 2514 4476 2994
rect 4158 2479 4214 2488
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4068 2372 4120 2378
rect 3988 2332 4068 2360
rect 3988 1834 4016 2332
rect 4068 2314 4120 2320
rect 4116 2204 4424 2224
rect 4116 2202 4122 2204
rect 4178 2202 4202 2204
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4424 2204
rect 4178 2150 4180 2202
rect 4360 2150 4362 2202
rect 4116 2148 4122 2150
rect 4178 2148 4202 2150
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4424 2150
rect 4116 2128 4424 2148
rect 4540 1970 4568 3046
rect 4724 2666 4752 4762
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 3602 4844 4626
rect 4908 4570 4936 4814
rect 4986 4791 5042 4800
rect 5000 4690 5028 4791
rect 5092 4729 5120 5306
rect 5184 5166 5212 5578
rect 5276 5386 5304 8384
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 5522 5396 7686
rect 5460 7449 5488 9318
rect 5666 9276 5974 9296
rect 5666 9274 5672 9276
rect 5728 9274 5752 9276
rect 5808 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5974 9276
rect 5728 9222 5730 9274
rect 5910 9222 5912 9274
rect 5666 9220 5672 9222
rect 5728 9220 5752 9222
rect 5808 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5974 9222
rect 5666 9200 5974 9220
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5446 7304 5502 7313
rect 5446 7239 5502 7248
rect 5460 6089 5488 7239
rect 5552 6662 5580 9007
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5920 8634 5948 8842
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5736 8430 5764 8570
rect 5920 8498 5948 8570
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 6012 8378 6040 12200
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6104 10062 6132 11630
rect 6196 11354 6224 11630
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6288 11354 6316 11562
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6274 10976 6330 10985
rect 6274 10911 6330 10920
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6104 9722 6132 9862
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6104 9586 6132 9658
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9081 6132 9318
rect 6090 9072 6146 9081
rect 6090 9007 6146 9016
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6104 8673 6132 8842
rect 6090 8664 6146 8673
rect 6090 8599 6146 8608
rect 6196 8537 6224 10406
rect 6288 10062 6316 10911
rect 6380 10674 6408 11086
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9897 6316 9998
rect 6274 9888 6330 9897
rect 6274 9823 6330 9832
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 8945 6316 9522
rect 6274 8936 6330 8945
rect 6274 8871 6330 8880
rect 6274 8800 6330 8809
rect 6274 8735 6330 8744
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 6012 8350 6132 8378
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5666 8188 5974 8208
rect 5666 8186 5672 8188
rect 5728 8186 5752 8188
rect 5808 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5974 8188
rect 5728 8134 5730 8186
rect 5910 8134 5912 8186
rect 5666 8132 5672 8134
rect 5728 8132 5752 8134
rect 5808 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5974 8134
rect 5666 8112 5974 8132
rect 6012 7954 6040 8230
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7478 5672 7822
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5666 7100 5974 7120
rect 5666 7098 5672 7100
rect 5728 7098 5752 7100
rect 5808 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5974 7100
rect 5728 7046 5730 7098
rect 5910 7046 5912 7098
rect 5666 7044 5672 7046
rect 5728 7044 5752 7046
rect 5808 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5974 7046
rect 5666 7024 5974 7044
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 6474 5672 6598
rect 5552 6446 5672 6474
rect 5446 6080 5502 6089
rect 5446 6015 5502 6024
rect 5552 5778 5580 6446
rect 5736 6225 5764 6870
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6390 5948 6666
rect 6012 6458 6040 7754
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5722 6216 5778 6225
rect 5722 6151 5778 6160
rect 5666 6012 5974 6032
rect 5666 6010 5672 6012
rect 5728 6010 5752 6012
rect 5808 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5974 6012
rect 5728 5958 5730 6010
rect 5910 5958 5912 6010
rect 5666 5956 5672 5958
rect 5728 5956 5752 5958
rect 5808 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5974 5958
rect 5666 5936 5974 5956
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5368 5494 5488 5522
rect 5276 5358 5396 5386
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5172 4752 5224 4758
rect 5078 4720 5134 4729
rect 4988 4684 5040 4690
rect 5172 4694 5224 4700
rect 5078 4655 5134 4664
rect 4988 4626 5040 4632
rect 4908 4542 5120 4570
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4894 3632 4950 3641
rect 4804 3596 4856 3602
rect 4894 3567 4950 3576
rect 4804 3538 4856 3544
rect 4908 2938 4936 3567
rect 5000 2990 5028 4422
rect 5092 3738 5120 4542
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3534 5212 4694
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4816 2910 4936 2938
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4816 2854 4844 2910
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4632 2638 4752 2666
rect 4908 2650 4936 2790
rect 4896 2644 4948 2650
rect 4632 2106 4660 2638
rect 4896 2586 4948 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4802 2544 4858 2553
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 4724 2038 4752 2518
rect 4802 2479 4858 2488
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4528 1964 4580 1970
rect 4528 1906 4580 1912
rect 3976 1828 4028 1834
rect 3976 1770 4028 1776
rect 4080 1494 4108 1906
rect 4816 1902 4844 2479
rect 4896 2440 4948 2446
rect 5092 2428 5120 3402
rect 5184 2650 5212 3470
rect 5276 2854 5304 5170
rect 5368 3641 5396 5358
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5354 3224 5410 3233
rect 5354 3159 5410 3168
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 4948 2400 5120 2428
rect 4896 2382 4948 2388
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5000 2038 5028 2246
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 5092 1902 5120 2400
rect 5276 2310 5304 2518
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4804 1896 4856 1902
rect 4804 1838 4856 1844
rect 5080 1896 5132 1902
rect 5080 1838 5132 1844
rect 4068 1488 4120 1494
rect 4068 1430 4120 1436
rect 4264 1358 4292 1838
rect 5184 1562 5212 2246
rect 5368 2106 5396 3159
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5460 2038 5488 5494
rect 5644 5114 5672 5782
rect 5816 5160 5868 5166
rect 5552 5086 5672 5114
rect 5814 5128 5816 5137
rect 5868 5128 5870 5137
rect 5552 4706 5580 5086
rect 5814 5063 5870 5072
rect 5666 4924 5974 4944
rect 5666 4922 5672 4924
rect 5728 4922 5752 4924
rect 5808 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5974 4924
rect 5728 4870 5730 4922
rect 5910 4870 5912 4922
rect 5666 4868 5672 4870
rect 5728 4868 5752 4870
rect 5808 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5974 4870
rect 5666 4848 5974 4868
rect 5814 4720 5870 4729
rect 5552 4678 5672 4706
rect 5540 4616 5592 4622
rect 5538 4584 5540 4593
rect 5592 4584 5594 4593
rect 5538 4519 5594 4528
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 3534 5580 4422
rect 5644 4010 5672 4678
rect 5814 4655 5870 4664
rect 5828 4049 5856 4655
rect 5906 4584 5962 4593
rect 5906 4519 5962 4528
rect 5814 4040 5870 4049
rect 5632 4004 5684 4010
rect 5814 3975 5870 3984
rect 5632 3946 5684 3952
rect 5920 3924 5948 4519
rect 6012 4146 6040 6258
rect 6104 5114 6132 8350
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6196 6202 6224 7278
rect 6288 6322 6316 8735
rect 6380 6934 6408 10610
rect 6472 7750 6500 12200
rect 8668 11960 8720 11966
rect 8668 11902 8720 11908
rect 20718 11928 20774 11937
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6550 11384 6606 11393
rect 6550 11319 6552 11328
rect 6604 11319 6606 11328
rect 6552 11290 6604 11296
rect 6564 10985 6592 11290
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6550 10976 6606 10985
rect 6550 10911 6606 10920
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 9722 6592 10610
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6550 9480 6606 9489
rect 6550 9415 6606 9424
rect 6564 8022 6592 9415
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8498 6684 8774
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6642 8392 6698 8401
rect 6642 8327 6698 8336
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7002 6592 7686
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6656 6440 6684 8327
rect 6564 6412 6684 6440
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6196 6174 6316 6202
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5234 6224 6054
rect 6288 5710 6316 6174
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5914 6408 6054
rect 6564 5953 6592 6412
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6550 5944 6606 5953
rect 6368 5908 6420 5914
rect 6550 5879 6606 5888
rect 6368 5850 6420 5856
rect 6656 5846 6684 6258
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6104 5086 6224 5114
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5920 3896 6040 3924
rect 5666 3836 5974 3856
rect 5666 3834 5672 3836
rect 5728 3834 5752 3836
rect 5808 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5974 3836
rect 5728 3782 5730 3834
rect 5910 3782 5912 3834
rect 5666 3780 5672 3782
rect 5728 3780 5752 3782
rect 5808 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5974 3782
rect 5666 3760 5974 3780
rect 5908 3664 5960 3670
rect 5814 3632 5870 3641
rect 5908 3606 5960 3612
rect 5814 3567 5870 3576
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5644 3176 5672 3402
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5552 3148 5672 3176
rect 5552 2310 5580 3148
rect 5736 3126 5764 3334
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5828 2961 5856 3567
rect 5920 3126 5948 3606
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5814 2952 5870 2961
rect 5814 2887 5870 2896
rect 5666 2748 5974 2768
rect 5666 2746 5672 2748
rect 5728 2746 5752 2748
rect 5808 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5974 2748
rect 5728 2694 5730 2746
rect 5910 2694 5912 2746
rect 5666 2692 5672 2694
rect 5728 2692 5752 2694
rect 5808 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5974 2694
rect 5666 2672 5974 2692
rect 6012 2650 6040 3896
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5816 2576 5868 2582
rect 5814 2544 5816 2553
rect 5868 2544 5870 2553
rect 5814 2479 5870 2488
rect 5724 2372 5776 2378
rect 5828 2360 5856 2479
rect 5776 2332 5856 2360
rect 5724 2314 5776 2320
rect 6104 2310 6132 4966
rect 6196 3233 6224 5086
rect 6288 4729 6316 5646
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6274 4720 6330 4729
rect 6274 4655 6330 4664
rect 6380 4570 6408 5578
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6288 4542 6408 4570
rect 6472 4570 6500 5510
rect 6564 4690 6592 5714
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6656 4865 6684 5238
rect 6642 4856 6698 4865
rect 6642 4791 6698 4800
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6748 4570 6776 11222
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 11014 6868 11086
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6932 10742 6960 11698
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11354 7420 11562
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7668 11354 7696 11494
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7760 11286 7788 11494
rect 7838 11384 7894 11393
rect 7838 11319 7840 11328
rect 7892 11319 7894 11328
rect 7840 11290 7892 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7564 11144 7616 11150
rect 7010 11112 7066 11121
rect 7564 11086 7616 11092
rect 7010 11047 7066 11056
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6918 9888 6974 9897
rect 6918 9823 6974 9832
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 8566 6868 9454
rect 6932 9160 6960 9823
rect 7024 9364 7052 11047
rect 7216 10908 7524 10928
rect 7216 10906 7222 10908
rect 7278 10906 7302 10908
rect 7358 10906 7382 10908
rect 7438 10906 7462 10908
rect 7518 10906 7524 10908
rect 7278 10854 7280 10906
rect 7460 10854 7462 10906
rect 7216 10852 7222 10854
rect 7278 10852 7302 10854
rect 7358 10852 7382 10854
rect 7438 10852 7462 10854
rect 7518 10852 7524 10854
rect 7216 10832 7524 10852
rect 7194 10704 7250 10713
rect 7194 10639 7250 10648
rect 7208 9908 7236 10639
rect 7470 10296 7526 10305
rect 7470 10231 7526 10240
rect 7484 10130 7512 10231
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7470 10024 7526 10033
rect 7470 9959 7472 9968
rect 7524 9959 7526 9968
rect 7472 9930 7524 9936
rect 7116 9880 7236 9908
rect 7116 9704 7144 9880
rect 7216 9820 7524 9840
rect 7216 9818 7222 9820
rect 7278 9818 7302 9820
rect 7358 9818 7382 9820
rect 7438 9818 7462 9820
rect 7518 9818 7524 9820
rect 7278 9766 7280 9818
rect 7460 9766 7462 9818
rect 7216 9764 7222 9766
rect 7278 9764 7302 9766
rect 7358 9764 7382 9766
rect 7438 9764 7462 9766
rect 7518 9764 7524 9766
rect 7216 9744 7524 9764
rect 7116 9676 7512 9704
rect 7104 9376 7156 9382
rect 7024 9336 7104 9364
rect 7104 9318 7156 9324
rect 6932 9132 7052 9160
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6932 7410 6960 8978
rect 7024 8906 7052 9132
rect 7484 8945 7512 9676
rect 7470 8936 7526 8945
rect 7012 8900 7064 8906
rect 7470 8871 7526 8880
rect 7012 8842 7064 8848
rect 7024 8673 7052 8842
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7886 7052 8230
rect 7116 7886 7144 8774
rect 7216 8732 7524 8752
rect 7216 8730 7222 8732
rect 7278 8730 7302 8732
rect 7358 8730 7382 8732
rect 7438 8730 7462 8732
rect 7518 8730 7524 8732
rect 7278 8678 7280 8730
rect 7460 8678 7462 8730
rect 7216 8676 7222 8678
rect 7278 8676 7302 8678
rect 7358 8676 7382 8678
rect 7438 8676 7462 8678
rect 7518 8676 7524 8678
rect 7216 8656 7524 8676
rect 7576 8634 7604 11086
rect 7852 10538 7880 11290
rect 8022 11248 8078 11257
rect 8022 11183 8078 11192
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7852 10266 7880 10474
rect 7840 10260 7892 10266
rect 7892 10220 7972 10248
rect 7840 10202 7892 10208
rect 7944 10169 7972 10220
rect 7930 10160 7986 10169
rect 7840 10124 7892 10130
rect 7930 10095 7986 10104
rect 7840 10066 7892 10072
rect 7654 9752 7710 9761
rect 7654 9687 7710 9696
rect 7668 9586 7696 9687
rect 7748 9686 7800 9692
rect 7748 9628 7800 9634
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 6860 6880 6866
rect 6932 6848 6960 7346
rect 7116 7002 7144 7822
rect 7216 7644 7524 7664
rect 7216 7642 7222 7644
rect 7278 7642 7302 7644
rect 7358 7642 7382 7644
rect 7438 7642 7462 7644
rect 7518 7642 7524 7644
rect 7278 7590 7280 7642
rect 7460 7590 7462 7642
rect 7216 7588 7222 7590
rect 7278 7588 7302 7590
rect 7358 7588 7382 7590
rect 7438 7588 7462 7590
rect 7518 7588 7524 7590
rect 7216 7568 7524 7588
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6880 6820 6960 6848
rect 6828 6802 6880 6808
rect 6932 5778 6960 6820
rect 7208 6730 7236 7210
rect 7576 6769 7604 8026
rect 7562 6760 7618 6769
rect 7012 6724 7064 6730
rect 7196 6724 7248 6730
rect 7012 6666 7064 6672
rect 7116 6684 7196 6712
rect 7024 5914 7052 6666
rect 7116 6440 7144 6684
rect 7562 6695 7618 6704
rect 7196 6666 7248 6672
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7216 6556 7524 6576
rect 7216 6554 7222 6556
rect 7278 6554 7302 6556
rect 7358 6554 7382 6556
rect 7438 6554 7462 6556
rect 7518 6554 7524 6556
rect 7278 6502 7280 6554
rect 7460 6502 7462 6554
rect 7216 6500 7222 6502
rect 7278 6500 7302 6502
rect 7358 6500 7382 6502
rect 7438 6500 7462 6502
rect 7518 6500 7524 6502
rect 7216 6480 7524 6500
rect 7116 6412 7236 6440
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6472 4554 6592 4570
rect 6472 4548 6604 4554
rect 6472 4542 6552 4548
rect 6288 4078 6316 4542
rect 6552 4490 6604 4496
rect 6735 4542 6776 4570
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6182 3224 6238 3233
rect 6182 3159 6238 3168
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6196 2582 6224 2994
rect 6288 2922 6316 4014
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5552 2038 5580 2246
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5264 1760 5316 1766
rect 5264 1702 5316 1708
rect 5172 1556 5224 1562
rect 5172 1498 5224 1504
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 5276 1290 5304 1702
rect 5666 1660 5974 1680
rect 5666 1658 5672 1660
rect 5728 1658 5752 1660
rect 5808 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5974 1660
rect 5728 1606 5730 1658
rect 5910 1606 5912 1658
rect 5666 1604 5672 1606
rect 5728 1604 5752 1606
rect 5808 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5974 1606
rect 5666 1584 5974 1604
rect 6288 1465 6316 2751
rect 6380 2446 6408 4422
rect 6472 4026 6500 4422
rect 6564 4146 6592 4490
rect 6735 4468 6763 4542
rect 6656 4440 6763 4468
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6472 3998 6592 4026
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 2582 6500 3878
rect 6564 3738 6592 3998
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 2650 6592 3470
rect 6656 2961 6684 4440
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6642 2952 6698 2961
rect 6642 2887 6698 2896
rect 6748 2904 6776 4218
rect 6840 3058 6868 5510
rect 7116 5352 7144 6054
rect 7208 5710 7236 6412
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7216 5468 7524 5488
rect 7216 5466 7222 5468
rect 7278 5466 7302 5468
rect 7358 5466 7382 5468
rect 7438 5466 7462 5468
rect 7518 5466 7524 5468
rect 7278 5414 7280 5466
rect 7460 5414 7462 5466
rect 7216 5412 7222 5414
rect 7278 5412 7302 5414
rect 7358 5412 7382 5414
rect 7438 5412 7462 5414
rect 7518 5412 7524 5414
rect 7216 5392 7524 5412
rect 6932 5324 7144 5352
rect 6932 4049 6960 5324
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7010 4584 7066 4593
rect 7010 4519 7066 4528
rect 6918 4040 6974 4049
rect 6918 3975 6974 3984
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3602 6960 3878
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 7024 2922 7052 4519
rect 7012 2916 7064 2922
rect 6748 2876 6960 2904
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6826 2816 6882 2825
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6656 1884 6684 2790
rect 6826 2751 6882 2760
rect 6840 2446 6868 2751
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 2038 6776 2314
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6932 1970 6960 2876
rect 7012 2858 7064 2864
rect 7116 2650 7144 5170
rect 7216 4380 7524 4400
rect 7216 4378 7222 4380
rect 7278 4378 7302 4380
rect 7358 4378 7382 4380
rect 7438 4378 7462 4380
rect 7518 4378 7524 4380
rect 7278 4326 7280 4378
rect 7460 4326 7462 4378
rect 7216 4324 7222 4326
rect 7278 4324 7302 4326
rect 7358 4324 7382 4326
rect 7438 4324 7462 4326
rect 7518 4324 7524 4326
rect 7216 4304 7524 4324
rect 7194 4176 7250 4185
rect 7194 4111 7250 4120
rect 7208 4078 7236 4111
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7216 3292 7524 3312
rect 7216 3290 7222 3292
rect 7278 3290 7302 3292
rect 7358 3290 7382 3292
rect 7438 3290 7462 3292
rect 7518 3290 7524 3292
rect 7278 3238 7280 3290
rect 7460 3238 7462 3290
rect 7216 3236 7222 3238
rect 7278 3236 7302 3238
rect 7358 3236 7382 3238
rect 7438 3236 7462 3238
rect 7518 3236 7524 3238
rect 7216 3216 7524 3236
rect 7576 3176 7604 6598
rect 7668 4457 7696 9318
rect 7760 6458 7788 9628
rect 7852 9042 7880 10066
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8090 7880 8774
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7944 7834 7972 9998
rect 8036 8566 8064 11183
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10742 8156 11086
rect 8116 10736 8168 10742
rect 8114 10704 8116 10713
rect 8168 10704 8170 10713
rect 8114 10639 8170 10648
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 9568 8156 10474
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10266 8248 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 8220 9722 8248 9959
rect 8312 9722 8340 11766
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8404 11354 8432 11698
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8128 9540 8340 9568
rect 8206 9480 8262 9489
rect 8206 9415 8262 9424
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 7852 7806 7972 7834
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7852 6338 7880 7806
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7760 6310 7880 6338
rect 7760 5409 7788 6310
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7654 4448 7710 4457
rect 7654 4383 7710 4392
rect 7760 4298 7788 5238
rect 7392 3148 7604 3176
rect 7668 4270 7788 4298
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7196 2984 7248 2990
rect 7300 2961 7328 3062
rect 7196 2926 7248 2932
rect 7286 2952 7342 2961
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7010 2408 7066 2417
rect 7208 2394 7236 2926
rect 7286 2887 7342 2896
rect 7300 2446 7328 2887
rect 7010 2343 7066 2352
rect 7116 2366 7236 2394
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7392 2394 7420 3148
rect 7668 2990 7696 4270
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2650 7604 2858
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7760 2446 7788 4150
rect 7852 3777 7880 6190
rect 7944 4570 7972 7686
rect 8128 7206 8156 7958
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8036 6866 8064 7142
rect 8024 6860 8076 6866
rect 8076 6820 8156 6848
rect 8024 6802 8076 6808
rect 8022 6760 8078 6769
rect 8022 6695 8078 6704
rect 8036 4690 8064 6695
rect 8128 6497 8156 6820
rect 8114 6488 8170 6497
rect 8114 6423 8170 6432
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8128 5370 8156 6326
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8220 4826 8248 9415
rect 8312 7993 8340 9540
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 7041 8340 7278
rect 8298 7032 8354 7041
rect 8298 6967 8354 6976
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8312 5642 8340 6870
rect 8404 6730 8432 11086
rect 8496 9926 8524 11222
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9382 8524 9862
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8496 8090 8524 8910
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8496 6866 8524 7822
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6225 8524 6598
rect 8588 6390 8616 11290
rect 8680 10810 8708 11902
rect 20718 11863 20774 11872
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 8766 11452 9074 11472
rect 8766 11450 8772 11452
rect 8828 11450 8852 11452
rect 8908 11450 8932 11452
rect 8988 11450 9012 11452
rect 9068 11450 9074 11452
rect 8828 11398 8830 11450
rect 9010 11398 9012 11450
rect 8766 11396 8772 11398
rect 8828 11396 8852 11398
rect 8908 11396 8932 11398
rect 8988 11396 9012 11398
rect 9068 11396 9074 11398
rect 8766 11376 9074 11396
rect 9140 11206 9352 11234
rect 9140 11150 9168 11206
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8680 8838 8708 10542
rect 8766 10364 9074 10384
rect 8766 10362 8772 10364
rect 8828 10362 8852 10364
rect 8908 10362 8932 10364
rect 8988 10362 9012 10364
rect 9068 10362 9074 10364
rect 8828 10310 8830 10362
rect 9010 10310 9012 10362
rect 8766 10308 8772 10310
rect 8828 10308 8852 10310
rect 8908 10308 8932 10310
rect 8988 10308 9012 10310
rect 9068 10308 9074 10310
rect 8766 10288 9074 10308
rect 8942 10160 8998 10169
rect 8942 10095 8998 10104
rect 8956 10062 8984 10095
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8766 9276 9074 9296
rect 8766 9274 8772 9276
rect 8828 9274 8852 9276
rect 8908 9274 8932 9276
rect 8988 9274 9012 9276
rect 9068 9274 9074 9276
rect 8828 9222 8830 9274
rect 9010 9222 9012 9274
rect 8766 9220 8772 9222
rect 8828 9220 8852 9222
rect 8908 9220 8932 9222
rect 8988 9220 9012 9222
rect 9068 9220 9074 9222
rect 8766 9200 9074 9220
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8482 6216 8538 6225
rect 8482 6151 8538 6160
rect 8680 5914 8708 8366
rect 8766 8188 9074 8208
rect 8766 8186 8772 8188
rect 8828 8186 8852 8188
rect 8908 8186 8932 8188
rect 8988 8186 9012 8188
rect 9068 8186 9074 8188
rect 8828 8134 8830 8186
rect 9010 8134 9012 8186
rect 8766 8132 8772 8134
rect 8828 8132 8852 8134
rect 8908 8132 8932 8134
rect 8988 8132 9012 8134
rect 9068 8132 9074 8134
rect 8766 8112 9074 8132
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 7313 9076 7346
rect 9034 7304 9090 7313
rect 9034 7239 9090 7248
rect 8766 7100 9074 7120
rect 8766 7098 8772 7100
rect 8828 7098 8852 7100
rect 8908 7098 8932 7100
rect 8988 7098 9012 7100
rect 9068 7098 9074 7100
rect 8828 7046 8830 7098
rect 9010 7046 9012 7098
rect 8766 7044 8772 7046
rect 8828 7044 8852 7046
rect 8908 7044 8932 7046
rect 8988 7044 9012 7046
rect 9068 7044 9074 7046
rect 8766 7024 9074 7044
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6186 8892 6598
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8766 6012 9074 6032
rect 8766 6010 8772 6012
rect 8828 6010 8852 6012
rect 8908 6010 8932 6012
rect 8988 6010 9012 6012
rect 9068 6010 9074 6012
rect 8828 5958 8830 6010
rect 9010 5958 9012 6010
rect 8766 5956 8772 5958
rect 8828 5956 8852 5958
rect 8908 5956 8932 5958
rect 8988 5956 9012 5958
rect 9068 5956 9074 5958
rect 8766 5936 9074 5956
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7944 4542 8064 4570
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4214 7972 4422
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7838 3768 7894 3777
rect 7838 3703 7894 3712
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7748 2440 7800 2446
rect 7392 2366 7604 2394
rect 7748 2382 7800 2388
rect 7024 2310 7052 2343
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7116 2106 7144 2366
rect 7216 2204 7524 2224
rect 7216 2202 7222 2204
rect 7278 2202 7302 2204
rect 7358 2202 7382 2204
rect 7438 2202 7462 2204
rect 7518 2202 7524 2204
rect 7278 2150 7280 2202
rect 7460 2150 7462 2202
rect 7216 2148 7222 2150
rect 7278 2148 7302 2150
rect 7358 2148 7382 2150
rect 7438 2148 7462 2150
rect 7518 2148 7524 2150
rect 7216 2128 7524 2148
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7576 2038 7604 2366
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7668 1970 7696 2314
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 2145 7788 2246
rect 7746 2136 7802 2145
rect 7852 2106 7880 3470
rect 7944 2106 7972 4014
rect 8036 3380 8064 4542
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4282 8156 4422
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8114 4176 8170 4185
rect 8114 4111 8170 4120
rect 8128 3505 8156 4111
rect 8220 3670 8248 4626
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8036 3352 8156 3380
rect 8022 3088 8078 3097
rect 8022 3023 8024 3032
rect 8076 3023 8078 3032
rect 8024 2994 8076 3000
rect 8128 2938 8156 3352
rect 8036 2910 8156 2938
rect 8220 2938 8248 3402
rect 8220 2910 8340 2938
rect 8036 2514 8064 2910
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8036 2281 8064 2314
rect 8022 2272 8078 2281
rect 8022 2207 8078 2216
rect 7746 2071 7802 2080
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8036 1970 8064 2207
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 6736 1896 6788 1902
rect 6656 1856 6736 1884
rect 6736 1838 6788 1844
rect 8128 1562 8156 2790
rect 8312 2666 8340 2910
rect 8220 2638 8340 2666
rect 8220 2106 8248 2638
rect 8300 2440 8352 2446
rect 8298 2408 8300 2417
rect 8352 2408 8354 2417
rect 8298 2343 8354 2352
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 6274 1456 6330 1465
rect 6274 1391 6330 1400
rect 8404 1442 8432 5102
rect 8496 3534 8524 5170
rect 8588 4758 8616 5850
rect 8666 5808 8722 5817
rect 8666 5743 8722 5752
rect 8680 4826 8708 5743
rect 8766 4924 9074 4944
rect 8766 4922 8772 4924
rect 8828 4922 8852 4924
rect 8908 4922 8932 4924
rect 8988 4922 9012 4924
rect 9068 4922 9074 4924
rect 8828 4870 8830 4922
rect 9010 4870 9012 4922
rect 8766 4868 8772 4870
rect 8828 4868 8852 4870
rect 8908 4868 8932 4870
rect 8988 4868 9012 4870
rect 9068 4868 9074 4870
rect 8766 4848 9074 4868
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8588 3738 8616 4082
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 1970 8524 3334
rect 8588 2417 8616 3538
rect 8680 3398 8708 4082
rect 8864 4078 8892 4490
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4282 8984 4422
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9140 4185 9168 10950
rect 9232 8498 9260 11018
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9232 7342 9260 8026
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6866 9260 7278
rect 9324 7274 9352 11206
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9416 9625 9444 10542
rect 9402 9616 9458 9625
rect 9508 9586 9536 11154
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 10713 9628 11086
rect 9586 10704 9642 10713
rect 9586 10639 9642 10648
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9402 9551 9458 9560
rect 9496 9580 9548 9586
rect 9416 9466 9444 9551
rect 9496 9522 9548 9528
rect 9416 9438 9536 9466
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 9178 9444 9318
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 7970 9536 9438
rect 9600 8090 9628 10474
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8265 9720 8842
rect 9784 8673 9812 11494
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9678 8256 9734 8265
rect 9678 8191 9734 8200
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9508 7942 9720 7970
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 4826 9260 6598
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 9034 4040 9090 4049
rect 9034 3975 9036 3984
rect 9088 3975 9090 3984
rect 9036 3946 9088 3952
rect 8766 3836 9074 3856
rect 8766 3834 8772 3836
rect 8828 3834 8852 3836
rect 8908 3834 8932 3836
rect 8988 3834 9012 3836
rect 9068 3834 9074 3836
rect 8828 3782 8830 3834
rect 9010 3782 9012 3834
rect 8766 3780 8772 3782
rect 8828 3780 8852 3782
rect 8908 3780 8932 3782
rect 8988 3780 9012 3782
rect 9068 3780 9074 3782
rect 8766 3760 9074 3780
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8850 3632 8906 3641
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8666 3088 8722 3097
rect 8666 3023 8722 3032
rect 8680 2990 8708 3023
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8772 2836 8800 3606
rect 8850 3567 8906 3576
rect 8864 3058 8892 3567
rect 9034 3496 9090 3505
rect 9034 3431 9090 3440
rect 9048 3194 9076 3431
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8956 2961 8984 3062
rect 9232 3058 9260 4626
rect 9324 3738 9352 6054
rect 9416 5710 9444 7686
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9508 5409 9536 7754
rect 9692 6746 9720 7942
rect 9876 7857 9904 11562
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9968 7041 9996 8570
rect 9954 7032 10010 7041
rect 9954 6967 10010 6976
rect 9600 6718 9720 6746
rect 9600 5930 9628 6718
rect 9600 5902 9812 5930
rect 9678 5808 9734 5817
rect 9678 5743 9734 5752
rect 9494 5400 9550 5409
rect 9494 5335 9550 5344
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9402 3360 9458 3369
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8942 2952 8998 2961
rect 8942 2887 8998 2896
rect 8680 2808 8800 2836
rect 9048 2836 9076 2994
rect 9218 2952 9274 2961
rect 9218 2887 9274 2896
rect 9048 2808 9168 2836
rect 8680 2632 8708 2808
rect 8766 2748 9074 2768
rect 8766 2746 8772 2748
rect 8828 2746 8852 2748
rect 8908 2746 8932 2748
rect 8988 2746 9012 2748
rect 9068 2746 9074 2748
rect 8828 2694 8830 2746
rect 9010 2694 9012 2746
rect 8766 2692 8772 2694
rect 8828 2692 8852 2694
rect 8908 2692 8932 2694
rect 8988 2692 9012 2694
rect 9068 2692 9074 2694
rect 8766 2672 9074 2692
rect 9140 2632 9168 2808
rect 9232 2650 9260 2887
rect 8680 2604 8800 2632
rect 8666 2544 8722 2553
rect 8666 2479 8722 2488
rect 8772 2496 8800 2604
rect 9048 2604 9168 2632
rect 9220 2644 9272 2650
rect 8680 2446 8708 2479
rect 8772 2468 8892 2496
rect 8668 2440 8720 2446
rect 8574 2408 8630 2417
rect 8668 2382 8720 2388
rect 8574 2343 8630 2352
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8864 1748 8892 2468
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8956 2281 8984 2314
rect 8942 2272 8998 2281
rect 8942 2207 8998 2216
rect 9048 2106 9076 2604
rect 9220 2586 9272 2592
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9140 2417 9168 2450
rect 9126 2408 9182 2417
rect 9126 2343 9182 2352
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 8680 1720 8892 1748
rect 8404 1426 8524 1442
rect 8404 1420 8536 1426
rect 8404 1414 8484 1420
rect 3424 1284 3476 1290
rect 3424 1226 3476 1232
rect 5264 1284 5316 1290
rect 5264 1226 5316 1232
rect 8404 1222 8432 1414
rect 8484 1362 8536 1368
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 3804 1018 3832 1158
rect 4116 1116 4424 1136
rect 4116 1114 4122 1116
rect 4178 1114 4202 1116
rect 4258 1114 4282 1116
rect 4338 1114 4362 1116
rect 4418 1114 4424 1116
rect 4178 1062 4180 1114
rect 4360 1062 4362 1114
rect 4116 1060 4122 1062
rect 4178 1060 4202 1062
rect 4258 1060 4282 1062
rect 4338 1060 4362 1062
rect 4418 1060 4424 1062
rect 4116 1040 4424 1060
rect 7216 1116 7524 1136
rect 7216 1114 7222 1116
rect 7278 1114 7302 1116
rect 7358 1114 7382 1116
rect 7438 1114 7462 1116
rect 7518 1114 7524 1116
rect 7278 1062 7280 1114
rect 7460 1062 7462 1114
rect 7216 1060 7222 1062
rect 7278 1060 7302 1062
rect 7358 1060 7382 1062
rect 7438 1060 7462 1062
rect 7518 1060 7524 1062
rect 7216 1040 7524 1060
rect 3792 1012 3844 1018
rect 3792 954 3844 960
rect 7944 950 7972 1158
rect 7932 944 7984 950
rect 7932 886 7984 892
rect 8588 882 8616 1294
rect 8680 1222 8708 1720
rect 8766 1660 9074 1680
rect 8766 1658 8772 1660
rect 8828 1658 8852 1660
rect 8908 1658 8932 1660
rect 8988 1658 9012 1660
rect 9068 1658 9074 1660
rect 8828 1606 8830 1658
rect 9010 1606 9012 1658
rect 8766 1604 8772 1606
rect 8828 1604 8852 1606
rect 8908 1604 8932 1606
rect 8988 1604 9012 1606
rect 9068 1604 9074 1606
rect 8766 1584 9074 1604
rect 9232 1222 9260 2246
rect 9324 2038 9352 3334
rect 9402 3295 9458 3304
rect 9416 2106 9444 3295
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9312 2032 9364 2038
rect 9312 1974 9364 1980
rect 9508 1834 9536 4014
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9232 921 9260 1158
rect 9218 912 9274 921
rect 8576 876 8628 882
rect 9218 847 9274 856
rect 8576 818 8628 824
rect 9416 513 9444 1362
rect 9600 1329 9628 4966
rect 9586 1320 9642 1329
rect 9586 1255 9642 1264
rect 9692 950 9720 5743
rect 9784 4622 9812 5902
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9876 2553 9904 5510
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9862 2544 9918 2553
rect 9862 2479 9918 2488
rect 9772 2440 9824 2446
rect 9968 2417 9996 5306
rect 10060 4010 10088 9823
rect 10428 6633 10456 11698
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16592 10334 16620 11047
rect 15200 10328 15252 10334
rect 15200 10270 15252 10276
rect 16580 10328 16632 10334
rect 16684 10305 16712 11630
rect 16580 10270 16632 10276
rect 16670 10296 16726 10305
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 10692 7676 10744 7682
rect 10692 7618 10744 7624
rect 10414 6624 10470 6633
rect 10414 6559 10470 6568
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9772 2382 9824 2388
rect 9954 2408 10010 2417
rect 9784 2145 9812 2382
rect 9954 2343 10010 2352
rect 9770 2136 9826 2145
rect 9770 2071 9826 2080
rect 10704 1018 10732 7618
rect 11060 7608 11112 7614
rect 11060 7550 11112 7556
rect 11072 5216 11100 7550
rect 13832 7546 13860 9007
rect 15212 7682 15240 10270
rect 16670 10231 16726 10240
rect 20732 8378 20760 11863
rect 22112 9722 22140 12271
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 20640 8350 20760 8378
rect 20640 7682 20668 8350
rect 15200 7676 15252 7682
rect 15200 7618 15252 7624
rect 20628 7676 20680 7682
rect 20628 7618 20680 7624
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 10980 5188 11100 5216
rect 10980 1494 11008 5188
rect 16580 5024 16632 5030
rect 16684 5001 16712 6054
rect 16580 4966 16632 4972
rect 16670 4992 16726 5001
rect 16592 4185 16620 4966
rect 16670 4927 16726 4936
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3777 16620 3878
rect 16578 3768 16634 3777
rect 16578 3703 16634 3712
rect 21376 2650 21404 9658
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 16670 2544 16726 2553
rect 16670 2479 16726 2488
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16592 2145 16620 2314
rect 16684 2310 16712 2479
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 16578 1728 16634 1737
rect 16578 1663 16634 1672
rect 10968 1488 11020 1494
rect 10968 1430 11020 1436
rect 10692 1012 10744 1018
rect 10692 954 10744 960
rect 9680 944 9732 950
rect 9680 886 9732 892
rect 16592 882 16620 1663
rect 16580 876 16632 882
rect 16580 818 16632 824
rect 9402 504 9458 513
rect 9402 439 9458 448
<< via2 >>
rect 22098 12280 22154 12336
rect 846 9560 902 9616
rect 1766 10956 1768 10976
rect 1768 10956 1820 10976
rect 1820 10956 1822 10976
rect 1766 10920 1822 10956
rect 1858 10804 1914 10840
rect 1858 10784 1860 10804
rect 1860 10784 1912 10804
rect 1912 10784 1914 10804
rect 1030 8472 1086 8528
rect 1398 10532 1454 10568
rect 1674 10648 1730 10704
rect 1398 10512 1400 10532
rect 1400 10512 1452 10532
rect 1452 10512 1454 10532
rect 1306 6160 1362 6216
rect 1490 9424 1546 9480
rect 1490 8744 1546 8800
rect 1858 9016 1914 9072
rect 2134 9016 2190 9072
rect 1950 8608 2006 8664
rect 1582 6840 1638 6896
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 3054 10804 3110 10840
rect 3054 10784 3056 10804
rect 3056 10784 3108 10804
rect 3108 10784 3110 10804
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2870 10104 2926 10160
rect 2410 9968 2466 10024
rect 2134 7928 2190 7984
rect 1858 5752 1914 5808
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2594 8916 2596 8936
rect 2596 8916 2648 8936
rect 2648 8916 2650 8936
rect 2594 8880 2650 8916
rect 2870 8744 2926 8800
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2686 5616 2742 5672
rect 2594 5072 2650 5128
rect 2594 4664 2650 4720
rect 2778 3168 2834 3224
rect 2502 2352 2558 2408
rect 3606 11228 3608 11248
rect 3608 11228 3660 11248
rect 3660 11228 3662 11248
rect 3606 11192 3662 11228
rect 3514 10104 3570 10160
rect 3054 5208 3110 5264
rect 3054 4528 3110 4584
rect 3790 10920 3846 10976
rect 3790 10240 3846 10296
rect 3514 8628 3570 8664
rect 3514 8608 3516 8628
rect 3516 8608 3568 8628
rect 3568 8608 3570 8628
rect 3422 6160 3478 6216
rect 3422 5752 3478 5808
rect 3330 4936 3386 4992
rect 3606 2760 3662 2816
rect 4122 10906 4178 10908
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4122 10854 4168 10906
rect 4168 10854 4178 10906
rect 4202 10854 4232 10906
rect 4232 10854 4244 10906
rect 4244 10854 4258 10906
rect 4282 10854 4296 10906
rect 4296 10854 4308 10906
rect 4308 10854 4338 10906
rect 4362 10854 4372 10906
rect 4372 10854 4418 10906
rect 4122 10852 4178 10854
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 4122 9818 4178 9820
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4122 9766 4168 9818
rect 4168 9766 4178 9818
rect 4202 9766 4232 9818
rect 4232 9766 4244 9818
rect 4244 9766 4258 9818
rect 4282 9766 4296 9818
rect 4296 9766 4308 9818
rect 4308 9766 4338 9818
rect 4362 9766 4372 9818
rect 4372 9766 4418 9818
rect 4122 9764 4178 9766
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 3974 9560 4030 9616
rect 4122 8730 4178 8732
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4122 8678 4168 8730
rect 4168 8678 4178 8730
rect 4202 8678 4232 8730
rect 4232 8678 4244 8730
rect 4244 8678 4258 8730
rect 4282 8678 4296 8730
rect 4296 8678 4308 8730
rect 4308 8678 4338 8730
rect 4362 8678 4372 8730
rect 4372 8678 4418 8730
rect 4122 8676 4178 8678
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4122 7642 4178 7644
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4122 7590 4168 7642
rect 4168 7590 4178 7642
rect 4202 7590 4232 7642
rect 4232 7590 4244 7642
rect 4244 7590 4258 7642
rect 4282 7590 4296 7642
rect 4296 7590 4308 7642
rect 4308 7590 4338 7642
rect 4362 7590 4372 7642
rect 4372 7590 4418 7642
rect 4122 7588 4178 7590
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 4122 6554 4178 6556
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4122 6502 4168 6554
rect 4168 6502 4178 6554
rect 4202 6502 4232 6554
rect 4232 6502 4244 6554
rect 4244 6502 4258 6554
rect 4282 6502 4296 6554
rect 4296 6502 4308 6554
rect 4308 6502 4338 6554
rect 4362 6502 4372 6554
rect 4372 6502 4418 6554
rect 4122 6500 4178 6502
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4526 6160 4582 6216
rect 4122 5466 4178 5468
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4122 5414 4168 5466
rect 4168 5414 4178 5466
rect 4202 5414 4232 5466
rect 4232 5414 4244 5466
rect 4244 5414 4258 5466
rect 4282 5414 4296 5466
rect 4296 5414 4308 5466
rect 4308 5414 4338 5466
rect 4362 5414 4372 5466
rect 4372 5414 4418 5466
rect 4122 5412 4178 5414
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 3974 4664 4030 4720
rect 4526 4820 4582 4856
rect 4526 4800 4528 4820
rect 4528 4800 4580 4820
rect 4580 4800 4582 4820
rect 4434 4528 4490 4584
rect 4122 4378 4178 4380
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4122 4326 4168 4378
rect 4168 4326 4178 4378
rect 4202 4326 4232 4378
rect 4232 4326 4244 4378
rect 4244 4326 4258 4378
rect 4282 4326 4296 4378
rect 4296 4326 4308 4378
rect 4308 4326 4338 4378
rect 4362 4326 4372 4378
rect 4372 4326 4418 4378
rect 4122 4324 4178 4326
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 3882 3984 3938 4040
rect 3790 3304 3846 3360
rect 4122 3290 4178 3292
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4122 3238 4168 3290
rect 4168 3238 4178 3290
rect 4202 3238 4232 3290
rect 4232 3238 4244 3290
rect 4244 3238 4258 3290
rect 4282 3238 4296 3290
rect 4296 3238 4308 3290
rect 4308 3238 4338 3290
rect 4362 3238 4372 3290
rect 4372 3238 4418 3290
rect 4122 3236 4178 3238
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 3974 3168 4030 3224
rect 4066 3032 4122 3088
rect 4710 8608 4766 8664
rect 4894 9424 4950 9480
rect 4894 8744 4950 8800
rect 4710 6024 4766 6080
rect 4802 5888 4858 5944
rect 4710 4936 4766 4992
rect 5446 11600 5502 11656
rect 5672 11450 5728 11452
rect 5752 11450 5808 11452
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5672 11398 5718 11450
rect 5718 11398 5728 11450
rect 5752 11398 5782 11450
rect 5782 11398 5794 11450
rect 5794 11398 5808 11450
rect 5832 11398 5846 11450
rect 5846 11398 5858 11450
rect 5858 11398 5888 11450
rect 5912 11398 5922 11450
rect 5922 11398 5968 11450
rect 5672 11396 5728 11398
rect 5752 11396 5808 11398
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5630 11092 5632 11112
rect 5632 11092 5684 11112
rect 5684 11092 5686 11112
rect 5170 10920 5226 10976
rect 5630 11056 5686 11092
rect 5722 10648 5778 10704
rect 5538 10512 5594 10568
rect 5672 10362 5728 10364
rect 5752 10362 5808 10364
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5672 10310 5718 10362
rect 5718 10310 5728 10362
rect 5752 10310 5782 10362
rect 5782 10310 5794 10362
rect 5794 10310 5808 10362
rect 5832 10310 5846 10362
rect 5846 10310 5858 10362
rect 5858 10310 5888 10362
rect 5912 10310 5922 10362
rect 5922 10310 5968 10362
rect 5672 10308 5728 10310
rect 5752 10308 5808 10310
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5722 9560 5778 9616
rect 5906 9424 5962 9480
rect 5354 9016 5410 9072
rect 5170 5888 5226 5944
rect 3606 1400 3662 1456
rect 4158 2488 4214 2544
rect 4122 2202 4178 2204
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4122 2150 4168 2202
rect 4168 2150 4178 2202
rect 4202 2150 4232 2202
rect 4232 2150 4244 2202
rect 4244 2150 4258 2202
rect 4282 2150 4296 2202
rect 4296 2150 4308 2202
rect 4308 2150 4338 2202
rect 4362 2150 4372 2202
rect 4372 2150 4418 2202
rect 4122 2148 4178 2150
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 4986 4800 5042 4856
rect 5672 9274 5728 9276
rect 5752 9274 5808 9276
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5672 9222 5718 9274
rect 5718 9222 5728 9274
rect 5752 9222 5782 9274
rect 5782 9222 5794 9274
rect 5794 9222 5808 9274
rect 5832 9222 5846 9274
rect 5846 9222 5858 9274
rect 5858 9222 5888 9274
rect 5912 9222 5922 9274
rect 5922 9222 5968 9274
rect 5672 9220 5728 9222
rect 5752 9220 5808 9222
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5538 9016 5594 9072
rect 5446 7384 5502 7440
rect 5446 7248 5502 7304
rect 6274 10920 6330 10976
rect 6090 9016 6146 9072
rect 6090 8608 6146 8664
rect 6274 9832 6330 9888
rect 6274 8880 6330 8936
rect 6274 8744 6330 8800
rect 6182 8472 6238 8528
rect 5672 8186 5728 8188
rect 5752 8186 5808 8188
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5672 8134 5718 8186
rect 5718 8134 5728 8186
rect 5752 8134 5782 8186
rect 5782 8134 5794 8186
rect 5794 8134 5808 8186
rect 5832 8134 5846 8186
rect 5846 8134 5858 8186
rect 5858 8134 5888 8186
rect 5912 8134 5922 8186
rect 5922 8134 5968 8186
rect 5672 8132 5728 8134
rect 5752 8132 5808 8134
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5672 7098 5728 7100
rect 5752 7098 5808 7100
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5672 7046 5718 7098
rect 5718 7046 5728 7098
rect 5752 7046 5782 7098
rect 5782 7046 5794 7098
rect 5794 7046 5808 7098
rect 5832 7046 5846 7098
rect 5846 7046 5858 7098
rect 5858 7046 5888 7098
rect 5912 7046 5922 7098
rect 5922 7046 5968 7098
rect 5672 7044 5728 7046
rect 5752 7044 5808 7046
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5446 6024 5502 6080
rect 5722 6160 5778 6216
rect 5672 6010 5728 6012
rect 5752 6010 5808 6012
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5672 5958 5718 6010
rect 5718 5958 5728 6010
rect 5752 5958 5782 6010
rect 5782 5958 5794 6010
rect 5794 5958 5808 6010
rect 5832 5958 5846 6010
rect 5846 5958 5858 6010
rect 5858 5958 5888 6010
rect 5912 5958 5922 6010
rect 5922 5958 5968 6010
rect 5672 5956 5728 5958
rect 5752 5956 5808 5958
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5078 4664 5134 4720
rect 4894 3576 4950 3632
rect 4802 2488 4858 2544
rect 5354 3576 5410 3632
rect 5354 3168 5410 3224
rect 5814 5108 5816 5128
rect 5816 5108 5868 5128
rect 5868 5108 5870 5128
rect 5814 5072 5870 5108
rect 5672 4922 5728 4924
rect 5752 4922 5808 4924
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5672 4870 5718 4922
rect 5718 4870 5728 4922
rect 5752 4870 5782 4922
rect 5782 4870 5794 4922
rect 5794 4870 5808 4922
rect 5832 4870 5846 4922
rect 5846 4870 5858 4922
rect 5858 4870 5888 4922
rect 5912 4870 5922 4922
rect 5922 4870 5968 4922
rect 5672 4868 5728 4870
rect 5752 4868 5808 4870
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5538 4564 5540 4584
rect 5540 4564 5592 4584
rect 5592 4564 5594 4584
rect 5538 4528 5594 4564
rect 5814 4664 5870 4720
rect 5906 4528 5962 4584
rect 5814 3984 5870 4040
rect 6550 11348 6606 11384
rect 6550 11328 6552 11348
rect 6552 11328 6604 11348
rect 6604 11328 6606 11348
rect 6550 10920 6606 10976
rect 6550 9424 6606 9480
rect 6642 8336 6698 8392
rect 6550 5888 6606 5944
rect 5672 3834 5728 3836
rect 5752 3834 5808 3836
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5672 3782 5718 3834
rect 5718 3782 5728 3834
rect 5752 3782 5782 3834
rect 5782 3782 5794 3834
rect 5794 3782 5808 3834
rect 5832 3782 5846 3834
rect 5846 3782 5858 3834
rect 5858 3782 5888 3834
rect 5912 3782 5922 3834
rect 5922 3782 5968 3834
rect 5672 3780 5728 3782
rect 5752 3780 5808 3782
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5814 3576 5870 3632
rect 5814 2896 5870 2952
rect 5672 2746 5728 2748
rect 5752 2746 5808 2748
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5672 2694 5718 2746
rect 5718 2694 5728 2746
rect 5752 2694 5782 2746
rect 5782 2694 5794 2746
rect 5794 2694 5808 2746
rect 5832 2694 5846 2746
rect 5846 2694 5858 2746
rect 5858 2694 5888 2746
rect 5912 2694 5922 2746
rect 5922 2694 5968 2746
rect 5672 2692 5728 2694
rect 5752 2692 5808 2694
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 5814 2524 5816 2544
rect 5816 2524 5868 2544
rect 5868 2524 5870 2544
rect 5814 2488 5870 2524
rect 6274 4664 6330 4720
rect 6642 4800 6698 4856
rect 7838 11348 7894 11384
rect 7838 11328 7840 11348
rect 7840 11328 7892 11348
rect 7892 11328 7894 11348
rect 7010 11056 7066 11112
rect 6918 9832 6974 9888
rect 7222 10906 7278 10908
rect 7302 10906 7358 10908
rect 7382 10906 7438 10908
rect 7462 10906 7518 10908
rect 7222 10854 7268 10906
rect 7268 10854 7278 10906
rect 7302 10854 7332 10906
rect 7332 10854 7344 10906
rect 7344 10854 7358 10906
rect 7382 10854 7396 10906
rect 7396 10854 7408 10906
rect 7408 10854 7438 10906
rect 7462 10854 7472 10906
rect 7472 10854 7518 10906
rect 7222 10852 7278 10854
rect 7302 10852 7358 10854
rect 7382 10852 7438 10854
rect 7462 10852 7518 10854
rect 7194 10648 7250 10704
rect 7470 10240 7526 10296
rect 7470 9988 7526 10024
rect 7470 9968 7472 9988
rect 7472 9968 7524 9988
rect 7524 9968 7526 9988
rect 7222 9818 7278 9820
rect 7302 9818 7358 9820
rect 7382 9818 7438 9820
rect 7462 9818 7518 9820
rect 7222 9766 7268 9818
rect 7268 9766 7278 9818
rect 7302 9766 7332 9818
rect 7332 9766 7344 9818
rect 7344 9766 7358 9818
rect 7382 9766 7396 9818
rect 7396 9766 7408 9818
rect 7408 9766 7438 9818
rect 7462 9766 7472 9818
rect 7472 9766 7518 9818
rect 7222 9764 7278 9766
rect 7302 9764 7358 9766
rect 7382 9764 7438 9766
rect 7462 9764 7518 9766
rect 7470 8880 7526 8936
rect 7010 8608 7066 8664
rect 7222 8730 7278 8732
rect 7302 8730 7358 8732
rect 7382 8730 7438 8732
rect 7462 8730 7518 8732
rect 7222 8678 7268 8730
rect 7268 8678 7278 8730
rect 7302 8678 7332 8730
rect 7332 8678 7344 8730
rect 7344 8678 7358 8730
rect 7382 8678 7396 8730
rect 7396 8678 7408 8730
rect 7408 8678 7438 8730
rect 7462 8678 7472 8730
rect 7472 8678 7518 8730
rect 7222 8676 7278 8678
rect 7302 8676 7358 8678
rect 7382 8676 7438 8678
rect 7462 8676 7518 8678
rect 8022 11192 8078 11248
rect 7930 10104 7986 10160
rect 7654 9696 7710 9752
rect 7222 7642 7278 7644
rect 7302 7642 7358 7644
rect 7382 7642 7438 7644
rect 7462 7642 7518 7644
rect 7222 7590 7268 7642
rect 7268 7590 7278 7642
rect 7302 7590 7332 7642
rect 7332 7590 7344 7642
rect 7344 7590 7358 7642
rect 7382 7590 7396 7642
rect 7396 7590 7408 7642
rect 7408 7590 7438 7642
rect 7462 7590 7472 7642
rect 7472 7590 7518 7642
rect 7222 7588 7278 7590
rect 7302 7588 7358 7590
rect 7382 7588 7438 7590
rect 7462 7588 7518 7590
rect 7562 6704 7618 6760
rect 7222 6554 7278 6556
rect 7302 6554 7358 6556
rect 7382 6554 7438 6556
rect 7462 6554 7518 6556
rect 7222 6502 7268 6554
rect 7268 6502 7278 6554
rect 7302 6502 7332 6554
rect 7332 6502 7344 6554
rect 7344 6502 7358 6554
rect 7382 6502 7396 6554
rect 7396 6502 7408 6554
rect 7408 6502 7438 6554
rect 7462 6502 7472 6554
rect 7472 6502 7518 6554
rect 7222 6500 7278 6502
rect 7302 6500 7358 6502
rect 7382 6500 7438 6502
rect 7462 6500 7518 6502
rect 6182 3168 6238 3224
rect 6274 2760 6330 2816
rect 5672 1658 5728 1660
rect 5752 1658 5808 1660
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5672 1606 5718 1658
rect 5718 1606 5728 1658
rect 5752 1606 5782 1658
rect 5782 1606 5794 1658
rect 5794 1606 5808 1658
rect 5832 1606 5846 1658
rect 5846 1606 5858 1658
rect 5858 1606 5888 1658
rect 5912 1606 5922 1658
rect 5922 1606 5968 1658
rect 5672 1604 5728 1606
rect 5752 1604 5808 1606
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 6642 2896 6698 2952
rect 7222 5466 7278 5468
rect 7302 5466 7358 5468
rect 7382 5466 7438 5468
rect 7462 5466 7518 5468
rect 7222 5414 7268 5466
rect 7268 5414 7278 5466
rect 7302 5414 7332 5466
rect 7332 5414 7344 5466
rect 7344 5414 7358 5466
rect 7382 5414 7396 5466
rect 7396 5414 7408 5466
rect 7408 5414 7438 5466
rect 7462 5414 7472 5466
rect 7472 5414 7518 5466
rect 7222 5412 7278 5414
rect 7302 5412 7358 5414
rect 7382 5412 7438 5414
rect 7462 5412 7518 5414
rect 7010 4528 7066 4584
rect 6918 3984 6974 4040
rect 6826 2760 6882 2816
rect 7222 4378 7278 4380
rect 7302 4378 7358 4380
rect 7382 4378 7438 4380
rect 7462 4378 7518 4380
rect 7222 4326 7268 4378
rect 7268 4326 7278 4378
rect 7302 4326 7332 4378
rect 7332 4326 7344 4378
rect 7344 4326 7358 4378
rect 7382 4326 7396 4378
rect 7396 4326 7408 4378
rect 7408 4326 7438 4378
rect 7462 4326 7472 4378
rect 7472 4326 7518 4378
rect 7222 4324 7278 4326
rect 7302 4324 7358 4326
rect 7382 4324 7438 4326
rect 7462 4324 7518 4326
rect 7194 4120 7250 4176
rect 7222 3290 7278 3292
rect 7302 3290 7358 3292
rect 7382 3290 7438 3292
rect 7462 3290 7518 3292
rect 7222 3238 7268 3290
rect 7268 3238 7278 3290
rect 7302 3238 7332 3290
rect 7332 3238 7344 3290
rect 7344 3238 7358 3290
rect 7382 3238 7396 3290
rect 7396 3238 7408 3290
rect 7408 3238 7438 3290
rect 7462 3238 7472 3290
rect 7472 3238 7518 3290
rect 7222 3236 7278 3238
rect 7302 3236 7358 3238
rect 7382 3236 7438 3238
rect 7462 3236 7518 3238
rect 8114 10684 8116 10704
rect 8116 10684 8168 10704
rect 8168 10684 8170 10704
rect 8114 10648 8170 10684
rect 8206 9968 8262 10024
rect 8206 9424 8262 9480
rect 7746 5344 7802 5400
rect 7654 4392 7710 4448
rect 7010 2352 7066 2408
rect 7286 2896 7342 2952
rect 8022 6704 8078 6760
rect 8114 6432 8170 6488
rect 8298 7928 8354 7984
rect 8298 6976 8354 7032
rect 20718 11872 20774 11928
rect 8772 11450 8828 11452
rect 8852 11450 8908 11452
rect 8932 11450 8988 11452
rect 9012 11450 9068 11452
rect 8772 11398 8818 11450
rect 8818 11398 8828 11450
rect 8852 11398 8882 11450
rect 8882 11398 8894 11450
rect 8894 11398 8908 11450
rect 8932 11398 8946 11450
rect 8946 11398 8958 11450
rect 8958 11398 8988 11450
rect 9012 11398 9022 11450
rect 9022 11398 9068 11450
rect 8772 11396 8828 11398
rect 8852 11396 8908 11398
rect 8932 11396 8988 11398
rect 9012 11396 9068 11398
rect 8772 10362 8828 10364
rect 8852 10362 8908 10364
rect 8932 10362 8988 10364
rect 9012 10362 9068 10364
rect 8772 10310 8818 10362
rect 8818 10310 8828 10362
rect 8852 10310 8882 10362
rect 8882 10310 8894 10362
rect 8894 10310 8908 10362
rect 8932 10310 8946 10362
rect 8946 10310 8958 10362
rect 8958 10310 8988 10362
rect 9012 10310 9022 10362
rect 9022 10310 9068 10362
rect 8772 10308 8828 10310
rect 8852 10308 8908 10310
rect 8932 10308 8988 10310
rect 9012 10308 9068 10310
rect 8942 10104 8998 10160
rect 8772 9274 8828 9276
rect 8852 9274 8908 9276
rect 8932 9274 8988 9276
rect 9012 9274 9068 9276
rect 8772 9222 8818 9274
rect 8818 9222 8828 9274
rect 8852 9222 8882 9274
rect 8882 9222 8894 9274
rect 8894 9222 8908 9274
rect 8932 9222 8946 9274
rect 8946 9222 8958 9274
rect 8958 9222 8988 9274
rect 9012 9222 9022 9274
rect 9022 9222 9068 9274
rect 8772 9220 8828 9222
rect 8852 9220 8908 9222
rect 8932 9220 8988 9222
rect 9012 9220 9068 9222
rect 8482 6160 8538 6216
rect 8772 8186 8828 8188
rect 8852 8186 8908 8188
rect 8932 8186 8988 8188
rect 9012 8186 9068 8188
rect 8772 8134 8818 8186
rect 8818 8134 8828 8186
rect 8852 8134 8882 8186
rect 8882 8134 8894 8186
rect 8894 8134 8908 8186
rect 8932 8134 8946 8186
rect 8946 8134 8958 8186
rect 8958 8134 8988 8186
rect 9012 8134 9022 8186
rect 9022 8134 9068 8186
rect 8772 8132 8828 8134
rect 8852 8132 8908 8134
rect 8932 8132 8988 8134
rect 9012 8132 9068 8134
rect 9034 7248 9090 7304
rect 8772 7098 8828 7100
rect 8852 7098 8908 7100
rect 8932 7098 8988 7100
rect 9012 7098 9068 7100
rect 8772 7046 8818 7098
rect 8818 7046 8828 7098
rect 8852 7046 8882 7098
rect 8882 7046 8894 7098
rect 8894 7046 8908 7098
rect 8932 7046 8946 7098
rect 8946 7046 8958 7098
rect 8958 7046 8988 7098
rect 9012 7046 9022 7098
rect 9022 7046 9068 7098
rect 8772 7044 8828 7046
rect 8852 7044 8908 7046
rect 8932 7044 8988 7046
rect 9012 7044 9068 7046
rect 8772 6010 8828 6012
rect 8852 6010 8908 6012
rect 8932 6010 8988 6012
rect 9012 6010 9068 6012
rect 8772 5958 8818 6010
rect 8818 5958 8828 6010
rect 8852 5958 8882 6010
rect 8882 5958 8894 6010
rect 8894 5958 8908 6010
rect 8932 5958 8946 6010
rect 8946 5958 8958 6010
rect 8958 5958 8988 6010
rect 9012 5958 9022 6010
rect 9022 5958 9068 6010
rect 8772 5956 8828 5958
rect 8852 5956 8908 5958
rect 8932 5956 8988 5958
rect 9012 5956 9068 5958
rect 7838 3712 7894 3768
rect 7222 2202 7278 2204
rect 7302 2202 7358 2204
rect 7382 2202 7438 2204
rect 7462 2202 7518 2204
rect 7222 2150 7268 2202
rect 7268 2150 7278 2202
rect 7302 2150 7332 2202
rect 7332 2150 7344 2202
rect 7344 2150 7358 2202
rect 7382 2150 7396 2202
rect 7396 2150 7408 2202
rect 7408 2150 7438 2202
rect 7462 2150 7472 2202
rect 7472 2150 7518 2202
rect 7222 2148 7278 2150
rect 7302 2148 7358 2150
rect 7382 2148 7438 2150
rect 7462 2148 7518 2150
rect 7746 2080 7802 2136
rect 8114 4120 8170 4176
rect 8114 3440 8170 3496
rect 8022 3052 8078 3088
rect 8022 3032 8024 3052
rect 8024 3032 8076 3052
rect 8076 3032 8078 3052
rect 8022 2216 8078 2272
rect 8298 2388 8300 2408
rect 8300 2388 8352 2408
rect 8352 2388 8354 2408
rect 8298 2352 8354 2388
rect 6274 1400 6330 1456
rect 8666 5752 8722 5808
rect 8772 4922 8828 4924
rect 8852 4922 8908 4924
rect 8932 4922 8988 4924
rect 9012 4922 9068 4924
rect 8772 4870 8818 4922
rect 8818 4870 8828 4922
rect 8852 4870 8882 4922
rect 8882 4870 8894 4922
rect 8894 4870 8908 4922
rect 8932 4870 8946 4922
rect 8946 4870 8958 4922
rect 8958 4870 8988 4922
rect 9012 4870 9022 4922
rect 9022 4870 9068 4922
rect 8772 4868 8828 4870
rect 8852 4868 8908 4870
rect 8932 4868 8988 4870
rect 9012 4868 9068 4870
rect 9402 9560 9458 9616
rect 9586 10648 9642 10704
rect 9770 8608 9826 8664
rect 9678 8200 9734 8256
rect 9126 4120 9182 4176
rect 9034 4004 9090 4040
rect 9034 3984 9036 4004
rect 9036 3984 9088 4004
rect 9088 3984 9090 4004
rect 8772 3834 8828 3836
rect 8852 3834 8908 3836
rect 8932 3834 8988 3836
rect 9012 3834 9068 3836
rect 8772 3782 8818 3834
rect 8818 3782 8828 3834
rect 8852 3782 8882 3834
rect 8882 3782 8894 3834
rect 8894 3782 8908 3834
rect 8932 3782 8946 3834
rect 8946 3782 8958 3834
rect 8958 3782 8988 3834
rect 9012 3782 9022 3834
rect 9022 3782 9068 3834
rect 8772 3780 8828 3782
rect 8852 3780 8908 3782
rect 8932 3780 8988 3782
rect 9012 3780 9068 3782
rect 8666 3032 8722 3088
rect 8850 3576 8906 3632
rect 9034 3440 9090 3496
rect 10046 9832 10102 9888
rect 9862 7792 9918 7848
rect 9954 6976 10010 7032
rect 9678 5752 9734 5808
rect 9494 5344 9550 5400
rect 8942 2896 8998 2952
rect 9218 2896 9274 2952
rect 8772 2746 8828 2748
rect 8852 2746 8908 2748
rect 8932 2746 8988 2748
rect 9012 2746 9068 2748
rect 8772 2694 8818 2746
rect 8818 2694 8828 2746
rect 8852 2694 8882 2746
rect 8882 2694 8894 2746
rect 8894 2694 8908 2746
rect 8932 2694 8946 2746
rect 8946 2694 8958 2746
rect 8958 2694 8988 2746
rect 9012 2694 9022 2746
rect 9022 2694 9068 2746
rect 8772 2692 8828 2694
rect 8852 2692 8908 2694
rect 8932 2692 8988 2694
rect 9012 2692 9068 2694
rect 8666 2488 8722 2544
rect 8574 2352 8630 2408
rect 8942 2216 8998 2272
rect 9126 2352 9182 2408
rect 4122 1114 4178 1116
rect 4202 1114 4258 1116
rect 4282 1114 4338 1116
rect 4362 1114 4418 1116
rect 4122 1062 4168 1114
rect 4168 1062 4178 1114
rect 4202 1062 4232 1114
rect 4232 1062 4244 1114
rect 4244 1062 4258 1114
rect 4282 1062 4296 1114
rect 4296 1062 4308 1114
rect 4308 1062 4338 1114
rect 4362 1062 4372 1114
rect 4372 1062 4418 1114
rect 4122 1060 4178 1062
rect 4202 1060 4258 1062
rect 4282 1060 4338 1062
rect 4362 1060 4418 1062
rect 7222 1114 7278 1116
rect 7302 1114 7358 1116
rect 7382 1114 7438 1116
rect 7462 1114 7518 1116
rect 7222 1062 7268 1114
rect 7268 1062 7278 1114
rect 7302 1062 7332 1114
rect 7332 1062 7344 1114
rect 7344 1062 7358 1114
rect 7382 1062 7396 1114
rect 7396 1062 7408 1114
rect 7408 1062 7438 1114
rect 7462 1062 7472 1114
rect 7472 1062 7518 1114
rect 7222 1060 7278 1062
rect 7302 1060 7358 1062
rect 7382 1060 7438 1062
rect 7462 1060 7518 1062
rect 8772 1658 8828 1660
rect 8852 1658 8908 1660
rect 8932 1658 8988 1660
rect 9012 1658 9068 1660
rect 8772 1606 8818 1658
rect 8818 1606 8828 1658
rect 8852 1606 8882 1658
rect 8882 1606 8894 1658
rect 8894 1606 8908 1658
rect 8932 1606 8946 1658
rect 8946 1606 8958 1658
rect 8958 1606 8988 1658
rect 9012 1606 9022 1658
rect 9022 1606 9068 1658
rect 8772 1604 8828 1606
rect 8852 1604 8908 1606
rect 8932 1604 8988 1606
rect 9012 1604 9068 1606
rect 9402 3304 9458 3360
rect 9218 856 9274 912
rect 9586 1264 9642 1320
rect 9862 2488 9918 2544
rect 16578 11056 16634 11112
rect 13818 9016 13874 9072
rect 10414 6568 10470 6624
rect 9954 2352 10010 2408
rect 9770 2080 9826 2136
rect 16670 10240 16726 10296
rect 16670 4936 16726 4992
rect 16578 4120 16634 4176
rect 16578 3712 16634 3768
rect 16670 2488 16726 2544
rect 16578 2080 16634 2136
rect 16578 1672 16634 1728
rect 9402 448 9458 504
<< metal3 >>
rect 14000 12336 34000 12368
rect 14000 12280 22098 12336
rect 22154 12280 34000 12336
rect 14000 12248 34000 12280
rect 14000 11928 34000 11960
rect 14000 11872 20718 11928
rect 20774 11872 34000 11928
rect 14000 11840 34000 11872
rect 5441 11658 5507 11661
rect 5441 11656 12450 11658
rect 5441 11600 5446 11656
rect 5502 11600 12450 11656
rect 5441 11598 12450 11600
rect 5441 11595 5507 11598
rect 12390 11522 12450 11598
rect 14000 11522 34000 11552
rect 12390 11462 34000 11522
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 5660 11456 5980 11457
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 11391 5980 11392
rect 8760 11456 9080 11457
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 14000 11432 34000 11462
rect 8760 11391 9080 11392
rect 6545 11386 6611 11389
rect 7833 11386 7899 11389
rect 6545 11384 7899 11386
rect 6545 11328 6550 11384
rect 6606 11328 7838 11384
rect 7894 11328 7899 11384
rect 6545 11326 7899 11328
rect 6545 11323 6611 11326
rect 7833 11323 7899 11326
rect 3601 11250 3667 11253
rect 8017 11250 8083 11253
rect 3601 11248 8083 11250
rect 3601 11192 3606 11248
rect 3662 11192 8022 11248
rect 8078 11192 8083 11248
rect 3601 11190 8083 11192
rect 3601 11187 3667 11190
rect 8017 11187 8083 11190
rect 5625 11114 5691 11117
rect 7005 11114 7071 11117
rect 5625 11112 7071 11114
rect 5625 11056 5630 11112
rect 5686 11056 7010 11112
rect 7066 11056 7071 11112
rect 5625 11054 7071 11056
rect 5625 11051 5691 11054
rect 7005 11051 7071 11054
rect 14000 11112 34000 11144
rect 14000 11056 16578 11112
rect 16634 11056 34000 11112
rect 14000 11024 34000 11056
rect 1761 10978 1827 10981
rect 3785 10978 3851 10981
rect 1761 10976 3851 10978
rect 1761 10920 1766 10976
rect 1822 10920 3790 10976
rect 3846 10920 3851 10976
rect 1761 10918 3851 10920
rect 1761 10915 1827 10918
rect 3785 10915 3851 10918
rect 5165 10978 5231 10981
rect 6269 10978 6335 10981
rect 6545 10978 6611 10981
rect 5165 10976 6611 10978
rect 5165 10920 5170 10976
rect 5226 10920 6274 10976
rect 6330 10920 6550 10976
rect 6606 10920 6611 10976
rect 5165 10918 6611 10920
rect 5165 10915 5231 10918
rect 6269 10915 6335 10918
rect 6545 10915 6611 10918
rect 4110 10912 4430 10913
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10847 4430 10848
rect 7210 10912 7530 10913
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 10847 7530 10848
rect 1853 10842 1919 10845
rect 3049 10842 3115 10845
rect 1853 10840 3115 10842
rect 1853 10784 1858 10840
rect 1914 10784 3054 10840
rect 3110 10784 3115 10840
rect 1853 10782 3115 10784
rect 1853 10779 1919 10782
rect 3049 10779 3115 10782
rect 1669 10706 1735 10709
rect 5717 10706 5783 10709
rect 1669 10704 5783 10706
rect 1669 10648 1674 10704
rect 1730 10648 5722 10704
rect 5778 10648 5783 10704
rect 1669 10646 5783 10648
rect 1669 10643 1735 10646
rect 5717 10643 5783 10646
rect 7189 10706 7255 10709
rect 8109 10706 8175 10709
rect 7189 10704 8175 10706
rect 7189 10648 7194 10704
rect 7250 10648 8114 10704
rect 8170 10648 8175 10704
rect 7189 10646 8175 10648
rect 7189 10643 7255 10646
rect 8109 10643 8175 10646
rect 9581 10706 9647 10709
rect 14000 10706 34000 10736
rect 9581 10704 34000 10706
rect 9581 10648 9586 10704
rect 9642 10648 34000 10704
rect 9581 10646 34000 10648
rect 9581 10643 9647 10646
rect 14000 10616 34000 10646
rect 1393 10570 1459 10573
rect 5533 10570 5599 10573
rect 1393 10568 5599 10570
rect 1393 10512 1398 10568
rect 1454 10512 5538 10568
rect 5594 10512 5599 10568
rect 1393 10510 5599 10512
rect 1393 10507 1459 10510
rect 5533 10507 5599 10510
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 5660 10368 5980 10369
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 10303 5980 10304
rect 8760 10368 9080 10369
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 10303 9080 10304
rect 3785 10298 3851 10301
rect 3190 10296 3851 10298
rect 3190 10240 3790 10296
rect 3846 10240 3851 10296
rect 3190 10238 3851 10240
rect 2865 10162 2931 10165
rect 3190 10162 3250 10238
rect 3785 10235 3851 10238
rect 7465 10298 7531 10301
rect 7465 10296 7850 10298
rect 7465 10240 7470 10296
rect 7526 10240 7850 10296
rect 7465 10238 7850 10240
rect 7465 10235 7531 10238
rect 2865 10160 3250 10162
rect 2865 10104 2870 10160
rect 2926 10104 3250 10160
rect 2865 10102 3250 10104
rect 3509 10162 3575 10165
rect 3509 10160 7666 10162
rect 3509 10104 3514 10160
rect 3570 10104 7666 10160
rect 3509 10102 7666 10104
rect 2865 10099 2931 10102
rect 3509 10099 3575 10102
rect 2405 10026 2471 10029
rect 7465 10026 7531 10029
rect 2405 10024 7531 10026
rect 2405 9968 2410 10024
rect 2466 9968 7470 10024
rect 7526 9968 7531 10024
rect 2405 9966 7531 9968
rect 2405 9963 2471 9966
rect 7465 9963 7531 9966
rect 6269 9890 6335 9893
rect 6913 9890 6979 9893
rect 6269 9888 6979 9890
rect 6269 9832 6274 9888
rect 6330 9832 6918 9888
rect 6974 9832 6979 9888
rect 6269 9830 6979 9832
rect 6269 9827 6335 9830
rect 6913 9827 6979 9830
rect 4110 9824 4430 9825
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 9759 4430 9760
rect 7210 9824 7530 9825
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 7210 9759 7530 9760
rect 7606 9757 7666 10102
rect 7790 10026 7850 10238
rect 14000 10296 34000 10328
rect 14000 10240 16670 10296
rect 16726 10240 34000 10296
rect 14000 10208 34000 10240
rect 7925 10162 7991 10165
rect 8937 10162 9003 10165
rect 7925 10160 9003 10162
rect 7925 10104 7930 10160
rect 7986 10104 8942 10160
rect 8998 10104 9003 10160
rect 7925 10102 9003 10104
rect 7925 10099 7991 10102
rect 8937 10099 9003 10102
rect 8201 10026 8267 10029
rect 7790 10024 8267 10026
rect 7790 9968 8206 10024
rect 8262 9968 8267 10024
rect 7790 9966 8267 9968
rect 8201 9963 8267 9966
rect 10041 9890 10107 9893
rect 14000 9890 34000 9920
rect 10041 9888 34000 9890
rect 10041 9832 10046 9888
rect 10102 9832 34000 9888
rect 10041 9830 34000 9832
rect 10041 9827 10107 9830
rect 14000 9800 34000 9830
rect 7606 9752 7715 9757
rect 7606 9696 7654 9752
rect 7710 9696 7715 9752
rect 7606 9694 7715 9696
rect 7649 9691 7715 9694
rect 841 9618 907 9621
rect 3969 9618 4035 9621
rect 841 9616 4035 9618
rect 841 9560 846 9616
rect 902 9560 3974 9616
rect 4030 9560 4035 9616
rect 841 9558 4035 9560
rect 841 9555 907 9558
rect 3969 9555 4035 9558
rect 5717 9618 5783 9621
rect 9397 9618 9463 9621
rect 5717 9616 9463 9618
rect 5717 9560 5722 9616
rect 5778 9560 9402 9616
rect 9458 9560 9463 9616
rect 5717 9558 9463 9560
rect 5717 9555 5783 9558
rect 9397 9555 9463 9558
rect 1485 9482 1551 9485
rect 4889 9482 4955 9485
rect 1485 9480 4955 9482
rect 1485 9424 1490 9480
rect 1546 9424 4894 9480
rect 4950 9424 4955 9480
rect 1485 9422 4955 9424
rect 1485 9419 1551 9422
rect 4889 9419 4955 9422
rect 5901 9482 5967 9485
rect 6545 9482 6611 9485
rect 5901 9480 6611 9482
rect 5901 9424 5906 9480
rect 5962 9424 6550 9480
rect 6606 9424 6611 9480
rect 5901 9422 6611 9424
rect 5901 9419 5967 9422
rect 6545 9419 6611 9422
rect 8201 9482 8267 9485
rect 14000 9482 34000 9512
rect 8201 9480 34000 9482
rect 8201 9424 8206 9480
rect 8262 9424 34000 9480
rect 8201 9422 34000 9424
rect 8201 9419 8267 9422
rect 14000 9392 34000 9422
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 5660 9280 5980 9281
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 9215 5980 9216
rect 8760 9280 9080 9281
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 9215 9080 9216
rect 1853 9074 1919 9077
rect 2129 9074 2195 9077
rect 5349 9074 5415 9077
rect 1853 9072 1962 9074
rect 1853 9016 1858 9072
rect 1914 9016 1962 9072
rect 1853 9011 1962 9016
rect 2129 9072 5415 9074
rect 2129 9016 2134 9072
rect 2190 9016 5354 9072
rect 5410 9016 5415 9072
rect 2129 9014 5415 9016
rect 2129 9011 2195 9014
rect 5349 9011 5415 9014
rect 5533 9074 5599 9077
rect 6085 9074 6151 9077
rect 5533 9072 6151 9074
rect 5533 9016 5538 9072
rect 5594 9016 6090 9072
rect 6146 9016 6151 9072
rect 5533 9014 6151 9016
rect 5533 9011 5599 9014
rect 6085 9011 6151 9014
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 1485 8802 1551 8805
rect 1902 8802 1962 9011
rect 14000 8984 34000 9014
rect 2589 8938 2655 8941
rect 6269 8938 6335 8941
rect 2589 8936 6335 8938
rect 2589 8880 2594 8936
rect 2650 8880 6274 8936
rect 6330 8880 6335 8936
rect 2589 8878 6335 8880
rect 2589 8875 2655 8878
rect 6269 8875 6335 8878
rect 7465 8938 7531 8941
rect 7465 8936 7666 8938
rect 7465 8880 7470 8936
rect 7526 8880 7666 8936
rect 7465 8878 7666 8880
rect 7465 8875 7531 8878
rect 2865 8802 2931 8805
rect 1485 8800 2931 8802
rect 1485 8744 1490 8800
rect 1546 8744 2870 8800
rect 2926 8744 2931 8800
rect 1485 8742 2931 8744
rect 1485 8739 1551 8742
rect 2865 8739 2931 8742
rect 4889 8802 4955 8805
rect 6269 8802 6335 8805
rect 4889 8800 6335 8802
rect 4889 8744 4894 8800
rect 4950 8744 6274 8800
rect 6330 8744 6335 8800
rect 4889 8742 6335 8744
rect 4889 8739 4955 8742
rect 6269 8739 6335 8742
rect 4110 8736 4430 8737
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 8671 4430 8672
rect 7210 8736 7530 8737
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 8671 7530 8672
rect 1945 8666 2011 8669
rect 3509 8666 3575 8669
rect 1945 8664 3575 8666
rect 1945 8608 1950 8664
rect 2006 8608 3514 8664
rect 3570 8608 3575 8664
rect 1945 8606 3575 8608
rect 1945 8603 2011 8606
rect 3509 8603 3575 8606
rect 4705 8666 4771 8669
rect 6085 8666 6151 8669
rect 7005 8666 7071 8669
rect 4705 8664 7071 8666
rect 4705 8608 4710 8664
rect 4766 8608 6090 8664
rect 6146 8608 7010 8664
rect 7066 8608 7071 8664
rect 4705 8606 7071 8608
rect 4705 8603 4771 8606
rect 6085 8603 6151 8606
rect 7005 8603 7071 8606
rect 1025 8530 1091 8533
rect 6177 8530 6243 8533
rect 1025 8528 6243 8530
rect 1025 8472 1030 8528
rect 1086 8472 6182 8528
rect 6238 8472 6243 8528
rect 1025 8470 6243 8472
rect 1025 8467 1091 8470
rect 6177 8467 6243 8470
rect 6637 8394 6703 8397
rect 7606 8394 7666 8878
rect 9765 8666 9831 8669
rect 14000 8666 34000 8696
rect 9765 8664 34000 8666
rect 9765 8608 9770 8664
rect 9826 8608 34000 8664
rect 9765 8606 34000 8608
rect 9765 8603 9831 8606
rect 14000 8576 34000 8606
rect 6637 8392 7666 8394
rect 6637 8336 6642 8392
rect 6698 8336 7666 8392
rect 6637 8334 7666 8336
rect 6637 8331 6703 8334
rect 9673 8258 9739 8261
rect 14000 8258 34000 8288
rect 9673 8256 34000 8258
rect 9673 8200 9678 8256
rect 9734 8200 34000 8256
rect 9673 8198 34000 8200
rect 9673 8195 9739 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 5660 8192 5980 8193
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 8127 5980 8128
rect 8760 8192 9080 8193
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 14000 8168 34000 8198
rect 8760 8127 9080 8128
rect 2129 7986 2195 7989
rect 8293 7986 8359 7989
rect 2129 7984 8359 7986
rect 2129 7928 2134 7984
rect 2190 7928 8298 7984
rect 8354 7928 8359 7984
rect 2129 7926 8359 7928
rect 2129 7923 2195 7926
rect 8293 7923 8359 7926
rect 9857 7850 9923 7853
rect 14000 7850 34000 7880
rect 9857 7848 34000 7850
rect 9857 7792 9862 7848
rect 9918 7792 34000 7848
rect 9857 7790 34000 7792
rect 9857 7787 9923 7790
rect 14000 7760 34000 7790
rect 4110 7648 4430 7649
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7583 4430 7584
rect 7210 7648 7530 7649
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 7583 7530 7584
rect 5441 7442 5507 7445
rect 14000 7442 34000 7472
rect 5441 7440 34000 7442
rect 5441 7384 5446 7440
rect 5502 7384 34000 7440
rect 5441 7382 34000 7384
rect 5441 7379 5507 7382
rect 14000 7352 34000 7382
rect 5441 7306 5507 7309
rect 9029 7306 9095 7309
rect 5441 7304 9095 7306
rect 5441 7248 5446 7304
rect 5502 7248 9034 7304
rect 9090 7248 9095 7304
rect 5441 7246 9095 7248
rect 5441 7243 5507 7246
rect 9029 7243 9095 7246
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 5660 7104 5980 7105
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 7039 5980 7040
rect 8760 7104 9080 7105
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 7039 9080 7040
rect 8293 7034 8359 7037
rect 6134 7032 8359 7034
rect 6134 6976 8298 7032
rect 8354 6976 8359 7032
rect 6134 6974 8359 6976
rect 1577 6898 1643 6901
rect 6134 6898 6194 6974
rect 8293 6971 8359 6974
rect 9949 7034 10015 7037
rect 14000 7034 34000 7064
rect 9949 7032 34000 7034
rect 9949 6976 9954 7032
rect 10010 6976 34000 7032
rect 9949 6974 34000 6976
rect 9949 6971 10015 6974
rect 14000 6944 34000 6974
rect 1577 6896 6194 6898
rect 1577 6840 1582 6896
rect 1638 6840 6194 6896
rect 1577 6838 6194 6840
rect 1577 6835 1643 6838
rect 7557 6762 7623 6765
rect 8017 6762 8083 6765
rect 7557 6760 8083 6762
rect 7557 6704 7562 6760
rect 7618 6704 8022 6760
rect 8078 6704 8083 6760
rect 7557 6702 8083 6704
rect 7557 6699 7623 6702
rect 8017 6699 8083 6702
rect 10409 6626 10475 6629
rect 14000 6626 34000 6656
rect 10409 6624 34000 6626
rect 10409 6568 10414 6624
rect 10470 6568 34000 6624
rect 10409 6566 34000 6568
rect 10409 6563 10475 6566
rect 4110 6560 4430 6561
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 6495 4430 6496
rect 7210 6560 7530 6561
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 14000 6536 34000 6566
rect 7210 6495 7530 6496
rect 8109 6490 8175 6493
rect 8109 6488 8218 6490
rect 8109 6432 8114 6488
rect 8170 6432 8218 6488
rect 8109 6427 8218 6432
rect 1301 6218 1367 6221
rect 3417 6218 3483 6221
rect 1301 6216 3483 6218
rect 1301 6160 1306 6216
rect 1362 6160 3422 6216
rect 3478 6160 3483 6216
rect 1301 6158 3483 6160
rect 1301 6155 1367 6158
rect 3417 6155 3483 6158
rect 4521 6218 4587 6221
rect 5717 6218 5783 6221
rect 4521 6216 5783 6218
rect 4521 6160 4526 6216
rect 4582 6160 5722 6216
rect 5778 6160 5783 6216
rect 4521 6158 5783 6160
rect 4521 6155 4587 6158
rect 5717 6155 5783 6158
rect 4705 6082 4771 6085
rect 5441 6082 5507 6085
rect 4705 6080 5507 6082
rect 4705 6024 4710 6080
rect 4766 6024 5446 6080
rect 5502 6024 5507 6080
rect 4705 6022 5507 6024
rect 4705 6019 4771 6022
rect 5441 6019 5507 6022
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 5660 6016 5980 6017
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5951 5980 5952
rect 4797 5946 4863 5949
rect 5165 5946 5231 5949
rect 4797 5944 5231 5946
rect 4797 5888 4802 5944
rect 4858 5888 5170 5944
rect 5226 5888 5231 5944
rect 4797 5886 5231 5888
rect 4797 5883 4863 5886
rect 5165 5883 5231 5886
rect 6545 5944 6611 5949
rect 6545 5888 6550 5944
rect 6606 5888 6611 5944
rect 6545 5883 6611 5888
rect 1853 5810 1919 5813
rect 3417 5810 3483 5813
rect 6548 5810 6608 5883
rect 1853 5808 3483 5810
rect 1853 5752 1858 5808
rect 1914 5752 3422 5808
rect 3478 5752 3483 5808
rect 1853 5750 3483 5752
rect 1853 5747 1919 5750
rect 3417 5747 3483 5750
rect 5490 5750 6608 5810
rect 8158 5810 8218 6427
rect 8477 6218 8543 6221
rect 14000 6218 34000 6248
rect 8477 6216 34000 6218
rect 8477 6160 8482 6216
rect 8538 6160 34000 6216
rect 8477 6158 34000 6160
rect 8477 6155 8543 6158
rect 14000 6128 34000 6158
rect 8760 6016 9080 6017
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 5951 9080 5952
rect 8661 5810 8727 5813
rect 8158 5808 8727 5810
rect 8158 5752 8666 5808
rect 8722 5752 8727 5808
rect 8158 5750 8727 5752
rect 2681 5674 2747 5677
rect 5490 5674 5550 5750
rect 8661 5747 8727 5750
rect 9673 5810 9739 5813
rect 14000 5810 34000 5840
rect 9673 5808 34000 5810
rect 9673 5752 9678 5808
rect 9734 5752 34000 5808
rect 9673 5750 34000 5752
rect 9673 5747 9739 5750
rect 14000 5720 34000 5750
rect 2681 5672 5550 5674
rect 2681 5616 2686 5672
rect 2742 5616 5550 5672
rect 2681 5614 5550 5616
rect 2681 5611 2747 5614
rect 4110 5472 4430 5473
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 5407 4430 5408
rect 7210 5472 7530 5473
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 5407 7530 5408
rect 7741 5402 7807 5405
rect 7606 5400 7807 5402
rect 7606 5344 7746 5400
rect 7802 5344 7807 5400
rect 7606 5342 7807 5344
rect 3049 5266 3115 5269
rect 7606 5266 7666 5342
rect 7741 5339 7807 5342
rect 9489 5402 9555 5405
rect 14000 5402 34000 5432
rect 9489 5400 34000 5402
rect 9489 5344 9494 5400
rect 9550 5344 34000 5400
rect 9489 5342 34000 5344
rect 9489 5339 9555 5342
rect 14000 5312 34000 5342
rect 3049 5264 7666 5266
rect 3049 5208 3054 5264
rect 3110 5208 7666 5264
rect 3049 5206 7666 5208
rect 3049 5203 3115 5206
rect 2589 5130 2655 5133
rect 5809 5130 5875 5133
rect 2589 5128 5875 5130
rect 2589 5072 2594 5128
rect 2650 5072 5814 5128
rect 5870 5072 5875 5128
rect 2589 5070 5875 5072
rect 2589 5067 2655 5070
rect 5809 5067 5875 5070
rect 3325 4994 3391 4997
rect 4705 4994 4771 4997
rect 3325 4992 4771 4994
rect 3325 4936 3330 4992
rect 3386 4936 4710 4992
rect 4766 4936 4771 4992
rect 3325 4934 4771 4936
rect 3325 4931 3391 4934
rect 4705 4931 4771 4934
rect 14000 4992 34000 5024
rect 14000 4936 16670 4992
rect 16726 4936 34000 4992
rect 5660 4928 5980 4929
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4863 5980 4864
rect 8760 4928 9080 4929
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 14000 4904 34000 4936
rect 8760 4863 9080 4864
rect 4521 4858 4587 4861
rect 4981 4858 5047 4861
rect 4521 4856 5047 4858
rect 4521 4800 4526 4856
rect 4582 4800 4986 4856
rect 5042 4800 5047 4856
rect 4521 4798 5047 4800
rect 4521 4795 4587 4798
rect 4981 4795 5047 4798
rect 6637 4856 6703 4861
rect 6637 4800 6642 4856
rect 6698 4800 6703 4856
rect 6637 4795 6703 4800
rect 2589 4722 2655 4725
rect 3969 4722 4035 4725
rect 2589 4720 4035 4722
rect 2589 4664 2594 4720
rect 2650 4664 3974 4720
rect 4030 4664 4035 4720
rect 2589 4662 4035 4664
rect 2589 4659 2655 4662
rect 3969 4659 4035 4662
rect 5073 4722 5139 4725
rect 5809 4722 5875 4725
rect 6269 4722 6335 4725
rect 5073 4720 5458 4722
rect 5073 4664 5078 4720
rect 5134 4664 5458 4720
rect 5073 4662 5458 4664
rect 5073 4659 5139 4662
rect 3049 4586 3115 4589
rect 4429 4586 4495 4589
rect 3049 4584 4495 4586
rect 3049 4528 3054 4584
rect 3110 4528 4434 4584
rect 4490 4528 4495 4584
rect 3049 4526 4495 4528
rect 5398 4586 5458 4662
rect 5809 4720 6335 4722
rect 5809 4664 5814 4720
rect 5870 4664 6274 4720
rect 6330 4664 6335 4720
rect 5809 4662 6335 4664
rect 5809 4659 5875 4662
rect 6269 4659 6335 4662
rect 5533 4586 5599 4589
rect 5398 4584 5599 4586
rect 5398 4528 5538 4584
rect 5594 4528 5599 4584
rect 5398 4526 5599 4528
rect 3049 4523 3115 4526
rect 4429 4523 4495 4526
rect 5533 4523 5599 4526
rect 5901 4586 5967 4589
rect 6640 4586 6700 4795
rect 5901 4584 6700 4586
rect 5901 4528 5906 4584
rect 5962 4528 6700 4584
rect 5901 4526 6700 4528
rect 7005 4586 7071 4589
rect 14000 4586 34000 4616
rect 7005 4584 34000 4586
rect 7005 4528 7010 4584
rect 7066 4528 34000 4584
rect 7005 4526 34000 4528
rect 5901 4523 5967 4526
rect 7005 4523 7071 4526
rect 14000 4496 34000 4526
rect 7649 4448 7715 4453
rect 7649 4392 7654 4448
rect 7710 4392 7715 4448
rect 7649 4387 7715 4392
rect 4110 4384 4430 4385
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4319 4430 4320
rect 7210 4384 7530 4385
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 4319 7530 4320
rect 7189 4178 7255 4181
rect 3926 4176 7255 4178
rect 3926 4120 7194 4176
rect 7250 4120 7255 4176
rect 3926 4118 7255 4120
rect 7652 4178 7712 4387
rect 8109 4178 8175 4181
rect 9121 4178 9187 4181
rect 7652 4176 8175 4178
rect 7652 4120 8114 4176
rect 8170 4120 8175 4176
rect 7652 4118 8175 4120
rect 3926 4045 3986 4118
rect 7189 4115 7255 4118
rect 8109 4115 8175 4118
rect 8894 4176 9187 4178
rect 8894 4120 9126 4176
rect 9182 4120 9187 4176
rect 8894 4118 9187 4120
rect 3877 4040 3986 4045
rect 5809 4042 5875 4045
rect 3877 3984 3882 4040
rect 3938 3984 3986 4040
rect 3877 3982 3986 3984
rect 4708 4040 5875 4042
rect 4708 3984 5814 4040
rect 5870 3984 5875 4040
rect 4708 3982 5875 3984
rect 3877 3979 3943 3982
rect 3785 3362 3851 3365
rect 2484 3360 3851 3362
rect 2484 3304 3790 3360
rect 3846 3304 3851 3360
rect 2484 3302 3851 3304
rect 3785 3299 3851 3302
rect 4110 3296 4430 3297
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3231 4430 3232
rect 2773 3226 2839 3229
rect 3969 3226 4035 3229
rect 2773 3224 4035 3226
rect 2773 3168 2778 3224
rect 2834 3168 3974 3224
rect 4030 3168 4035 3224
rect 2773 3166 4035 3168
rect 2773 3163 2839 3166
rect 3969 3163 4035 3166
rect 4061 3090 4127 3093
rect 4708 3090 4768 3982
rect 5809 3979 5875 3982
rect 6913 4040 6979 4045
rect 8894 4042 8954 4118
rect 9121 4115 9187 4118
rect 14000 4176 34000 4208
rect 14000 4120 16578 4176
rect 16634 4120 34000 4176
rect 14000 4088 34000 4120
rect 6913 3984 6918 4040
rect 6974 3984 6979 4040
rect 6913 3979 6979 3984
rect 7054 3982 8954 4042
rect 9029 4042 9095 4045
rect 9029 4040 9276 4042
rect 9029 3984 9034 4040
rect 9090 3984 9276 4040
rect 9029 3982 9276 3984
rect 5660 3840 5980 3841
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 3775 5980 3776
rect 4889 3634 4955 3637
rect 5349 3634 5415 3637
rect 4889 3632 5415 3634
rect 4889 3576 4894 3632
rect 4950 3576 5354 3632
rect 5410 3576 5415 3632
rect 4889 3574 5415 3576
rect 4889 3571 4955 3574
rect 5349 3571 5415 3574
rect 5809 3634 5875 3637
rect 6916 3634 6976 3979
rect 5809 3632 6976 3634
rect 5809 3576 5814 3632
rect 5870 3576 6976 3632
rect 5809 3574 6976 3576
rect 5809 3571 5875 3574
rect 5349 3226 5415 3229
rect 6177 3226 6243 3229
rect 5349 3224 6243 3226
rect 5349 3168 5354 3224
rect 5410 3168 6182 3224
rect 6238 3168 6243 3224
rect 5349 3166 6243 3168
rect 5349 3163 5415 3166
rect 6177 3163 6243 3166
rect 7054 3090 7114 3982
rect 9029 3979 9095 3982
rect 8760 3840 9080 3841
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 3775 9080 3776
rect 7833 3770 7899 3773
rect 7833 3768 8586 3770
rect 7833 3712 7838 3768
rect 7894 3712 8586 3768
rect 7833 3710 8586 3712
rect 7833 3707 7899 3710
rect 8109 3498 8175 3501
rect 8526 3498 8586 3710
rect 8845 3634 8911 3637
rect 9216 3634 9276 3982
rect 14000 3768 34000 3800
rect 14000 3712 16578 3768
rect 16634 3712 34000 3768
rect 14000 3680 34000 3712
rect 8845 3632 9276 3634
rect 8845 3576 8850 3632
rect 8906 3576 9276 3632
rect 8845 3574 9276 3576
rect 8845 3571 8911 3574
rect 9029 3498 9095 3501
rect 8109 3496 8218 3498
rect 8109 3440 8114 3496
rect 8170 3440 8218 3496
rect 8109 3435 8218 3440
rect 8526 3496 9095 3498
rect 8526 3440 9034 3496
rect 9090 3440 9095 3496
rect 8526 3438 9095 3440
rect 9029 3435 9095 3438
rect 7210 3296 7530 3297
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 3231 7530 3232
rect 4061 3088 4768 3090
rect 4061 3032 4066 3088
rect 4122 3032 4768 3088
rect 4061 3030 4768 3032
rect 6272 3030 7114 3090
rect 8017 3090 8083 3093
rect 8158 3090 8218 3435
rect 9397 3362 9463 3365
rect 14000 3362 34000 3392
rect 9397 3360 34000 3362
rect 9397 3304 9402 3360
rect 9458 3304 34000 3360
rect 9397 3302 34000 3304
rect 9397 3299 9463 3302
rect 14000 3272 34000 3302
rect 8661 3090 8727 3093
rect 8017 3088 8218 3090
rect 8017 3032 8022 3088
rect 8078 3032 8218 3088
rect 8017 3030 8218 3032
rect 8342 3088 8727 3090
rect 8342 3032 8666 3088
rect 8722 3032 8727 3088
rect 8342 3030 8727 3032
rect 4061 3027 4127 3030
rect 5809 2954 5875 2957
rect 3742 2952 5875 2954
rect 3742 2896 5814 2952
rect 5870 2896 5875 2952
rect 3742 2894 5875 2896
rect 3601 2818 3667 2821
rect 3742 2818 3802 2894
rect 5809 2891 5875 2894
rect 6272 2821 6332 3030
rect 8017 3027 8083 3030
rect 6637 2952 6703 2957
rect 6637 2896 6642 2952
rect 6698 2896 6703 2952
rect 6637 2891 6703 2896
rect 7281 2954 7347 2957
rect 8342 2954 8402 3030
rect 8661 3027 8727 3030
rect 8937 2954 9003 2957
rect 7281 2952 8402 2954
rect 7281 2896 7286 2952
rect 7342 2896 8402 2952
rect 7281 2894 8402 2896
rect 8480 2952 9003 2954
rect 8480 2896 8942 2952
rect 8998 2896 9003 2952
rect 8480 2894 9003 2896
rect 7281 2891 7347 2894
rect 3601 2816 3802 2818
rect 3601 2760 3606 2816
rect 3662 2760 3802 2816
rect 3601 2758 3802 2760
rect 6269 2816 6335 2821
rect 6269 2760 6274 2816
rect 6330 2760 6335 2816
rect 3601 2755 3667 2758
rect 6269 2755 6335 2760
rect 5660 2752 5980 2753
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 2687 5980 2688
rect 4153 2546 4219 2549
rect 4797 2546 4863 2549
rect 4153 2544 4863 2546
rect 4153 2488 4158 2544
rect 4214 2488 4802 2544
rect 4858 2488 4863 2544
rect 4153 2486 4863 2488
rect 4153 2483 4219 2486
rect 4797 2483 4863 2486
rect 5809 2546 5875 2549
rect 6640 2546 6700 2891
rect 6821 2818 6887 2821
rect 8480 2818 8540 2894
rect 8937 2891 9003 2894
rect 9213 2954 9279 2957
rect 14000 2954 34000 2984
rect 9213 2952 34000 2954
rect 9213 2896 9218 2952
rect 9274 2896 34000 2952
rect 9213 2894 34000 2896
rect 9213 2891 9279 2894
rect 14000 2864 34000 2894
rect 6821 2816 8540 2818
rect 6821 2760 6826 2816
rect 6882 2760 8540 2816
rect 6821 2758 8540 2760
rect 6821 2755 6887 2758
rect 8760 2752 9080 2753
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 2687 9080 2688
rect 5809 2544 6700 2546
rect 5809 2488 5814 2544
rect 5870 2488 6700 2544
rect 5809 2486 6700 2488
rect 8661 2546 8727 2549
rect 9857 2546 9923 2549
rect 8661 2544 9923 2546
rect 8661 2488 8666 2544
rect 8722 2488 9862 2544
rect 9918 2488 9923 2544
rect 8661 2486 9923 2488
rect 5809 2483 5875 2486
rect 8661 2483 8727 2486
rect 9857 2483 9923 2486
rect 14000 2544 34000 2576
rect 14000 2488 16670 2544
rect 16726 2488 34000 2544
rect 14000 2456 34000 2488
rect 2497 2410 2563 2413
rect 7005 2410 7071 2413
rect 2497 2408 7071 2410
rect 2497 2352 2502 2408
rect 2558 2352 7010 2408
rect 7066 2352 7071 2408
rect 2497 2350 7071 2352
rect 2497 2347 2563 2350
rect 7005 2347 7071 2350
rect 8293 2410 8359 2413
rect 8569 2410 8635 2413
rect 8293 2408 8635 2410
rect 8293 2352 8298 2408
rect 8354 2352 8574 2408
rect 8630 2352 8635 2408
rect 8293 2350 8635 2352
rect 8293 2347 8359 2350
rect 8569 2347 8635 2350
rect 9121 2410 9187 2413
rect 9949 2410 10015 2413
rect 9121 2408 10015 2410
rect 9121 2352 9126 2408
rect 9182 2352 9954 2408
rect 10010 2352 10015 2408
rect 9121 2350 10015 2352
rect 9121 2347 9187 2350
rect 9949 2347 10015 2350
rect 8017 2274 8083 2277
rect 8937 2274 9003 2277
rect 8017 2272 9003 2274
rect 8017 2216 8022 2272
rect 8078 2216 8942 2272
rect 8998 2216 9003 2272
rect 8017 2214 9003 2216
rect 8017 2211 8083 2214
rect 8937 2211 9003 2214
rect 4110 2208 4430 2209
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 2143 4430 2144
rect 7210 2208 7530 2209
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 2143 7530 2144
rect 7741 2138 7807 2141
rect 9765 2138 9831 2141
rect 7741 2136 9831 2138
rect 7741 2080 7746 2136
rect 7802 2080 9770 2136
rect 9826 2080 9831 2136
rect 7741 2078 9831 2080
rect 7741 2075 7807 2078
rect 9765 2075 9831 2078
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 16578 1728
rect 16634 1672 34000 1728
rect 5660 1664 5980 1665
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1599 5980 1600
rect 8760 1664 9080 1665
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 14000 1640 34000 1672
rect 8760 1599 9080 1600
rect 3601 1458 3667 1461
rect 6269 1458 6335 1461
rect 3601 1456 6335 1458
rect 3601 1400 3606 1456
rect 3662 1400 6274 1456
rect 6330 1400 6335 1456
rect 3601 1398 6335 1400
rect 3601 1395 3667 1398
rect 6269 1395 6335 1398
rect 9581 1322 9647 1325
rect 14000 1322 34000 1352
rect 9581 1320 34000 1322
rect 9581 1264 9586 1320
rect 9642 1264 34000 1320
rect 9581 1262 34000 1264
rect 9581 1259 9647 1262
rect 14000 1232 34000 1262
rect 4110 1120 4430 1121
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 4110 1055 4430 1056
rect 7210 1120 7530 1121
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 7210 1055 7530 1056
rect 9213 914 9279 917
rect 14000 914 34000 944
rect 9213 912 34000 914
rect 9213 856 9218 912
rect 9274 856 34000 912
rect 9213 854 34000 856
rect 9213 851 9279 854
rect 14000 824 34000 854
rect 9397 506 9463 509
rect 14000 506 34000 536
rect 9397 504 34000 506
rect 9397 448 9402 504
rect 9458 448 34000 504
rect 9397 446 34000 448
rect 9397 443 9463 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 5668 11452 5732 11456
rect 5668 11396 5672 11452
rect 5672 11396 5728 11452
rect 5728 11396 5732 11452
rect 5668 11392 5732 11396
rect 5748 11452 5812 11456
rect 5748 11396 5752 11452
rect 5752 11396 5808 11452
rect 5808 11396 5812 11452
rect 5748 11392 5812 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 8768 11452 8832 11456
rect 8768 11396 8772 11452
rect 8772 11396 8828 11452
rect 8828 11396 8832 11452
rect 8768 11392 8832 11396
rect 8848 11452 8912 11456
rect 8848 11396 8852 11452
rect 8852 11396 8908 11452
rect 8908 11396 8912 11452
rect 8848 11392 8912 11396
rect 8928 11452 8992 11456
rect 8928 11396 8932 11452
rect 8932 11396 8988 11452
rect 8988 11396 8992 11452
rect 8928 11392 8992 11396
rect 9008 11452 9072 11456
rect 9008 11396 9012 11452
rect 9012 11396 9068 11452
rect 9068 11396 9072 11452
rect 9008 11392 9072 11396
rect 4118 10908 4182 10912
rect 4118 10852 4122 10908
rect 4122 10852 4178 10908
rect 4178 10852 4182 10908
rect 4118 10848 4182 10852
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 7218 10908 7282 10912
rect 7218 10852 7222 10908
rect 7222 10852 7278 10908
rect 7278 10852 7282 10908
rect 7218 10848 7282 10852
rect 7298 10908 7362 10912
rect 7298 10852 7302 10908
rect 7302 10852 7358 10908
rect 7358 10852 7362 10908
rect 7298 10848 7362 10852
rect 7378 10908 7442 10912
rect 7378 10852 7382 10908
rect 7382 10852 7438 10908
rect 7438 10852 7442 10908
rect 7378 10848 7442 10852
rect 7458 10908 7522 10912
rect 7458 10852 7462 10908
rect 7462 10852 7518 10908
rect 7518 10852 7522 10908
rect 7458 10848 7522 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 5668 10364 5732 10368
rect 5668 10308 5672 10364
rect 5672 10308 5728 10364
rect 5728 10308 5732 10364
rect 5668 10304 5732 10308
rect 5748 10364 5812 10368
rect 5748 10308 5752 10364
rect 5752 10308 5808 10364
rect 5808 10308 5812 10364
rect 5748 10304 5812 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 8768 10364 8832 10368
rect 8768 10308 8772 10364
rect 8772 10308 8828 10364
rect 8828 10308 8832 10364
rect 8768 10304 8832 10308
rect 8848 10364 8912 10368
rect 8848 10308 8852 10364
rect 8852 10308 8908 10364
rect 8908 10308 8912 10364
rect 8848 10304 8912 10308
rect 8928 10364 8992 10368
rect 8928 10308 8932 10364
rect 8932 10308 8988 10364
rect 8988 10308 8992 10364
rect 8928 10304 8992 10308
rect 9008 10364 9072 10368
rect 9008 10308 9012 10364
rect 9012 10308 9068 10364
rect 9068 10308 9072 10364
rect 9008 10304 9072 10308
rect 4118 9820 4182 9824
rect 4118 9764 4122 9820
rect 4122 9764 4178 9820
rect 4178 9764 4182 9820
rect 4118 9760 4182 9764
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 7218 9820 7282 9824
rect 7218 9764 7222 9820
rect 7222 9764 7278 9820
rect 7278 9764 7282 9820
rect 7218 9760 7282 9764
rect 7298 9820 7362 9824
rect 7298 9764 7302 9820
rect 7302 9764 7358 9820
rect 7358 9764 7362 9820
rect 7298 9760 7362 9764
rect 7378 9820 7442 9824
rect 7378 9764 7382 9820
rect 7382 9764 7438 9820
rect 7438 9764 7442 9820
rect 7378 9760 7442 9764
rect 7458 9820 7522 9824
rect 7458 9764 7462 9820
rect 7462 9764 7518 9820
rect 7518 9764 7522 9820
rect 7458 9760 7522 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 5668 9276 5732 9280
rect 5668 9220 5672 9276
rect 5672 9220 5728 9276
rect 5728 9220 5732 9276
rect 5668 9216 5732 9220
rect 5748 9276 5812 9280
rect 5748 9220 5752 9276
rect 5752 9220 5808 9276
rect 5808 9220 5812 9276
rect 5748 9216 5812 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 8768 9276 8832 9280
rect 8768 9220 8772 9276
rect 8772 9220 8828 9276
rect 8828 9220 8832 9276
rect 8768 9216 8832 9220
rect 8848 9276 8912 9280
rect 8848 9220 8852 9276
rect 8852 9220 8908 9276
rect 8908 9220 8912 9276
rect 8848 9216 8912 9220
rect 8928 9276 8992 9280
rect 8928 9220 8932 9276
rect 8932 9220 8988 9276
rect 8988 9220 8992 9276
rect 8928 9216 8992 9220
rect 9008 9276 9072 9280
rect 9008 9220 9012 9276
rect 9012 9220 9068 9276
rect 9068 9220 9072 9276
rect 9008 9216 9072 9220
rect 4118 8732 4182 8736
rect 4118 8676 4122 8732
rect 4122 8676 4178 8732
rect 4178 8676 4182 8732
rect 4118 8672 4182 8676
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 7218 8732 7282 8736
rect 7218 8676 7222 8732
rect 7222 8676 7278 8732
rect 7278 8676 7282 8732
rect 7218 8672 7282 8676
rect 7298 8732 7362 8736
rect 7298 8676 7302 8732
rect 7302 8676 7358 8732
rect 7358 8676 7362 8732
rect 7298 8672 7362 8676
rect 7378 8732 7442 8736
rect 7378 8676 7382 8732
rect 7382 8676 7438 8732
rect 7438 8676 7442 8732
rect 7378 8672 7442 8676
rect 7458 8732 7522 8736
rect 7458 8676 7462 8732
rect 7462 8676 7518 8732
rect 7518 8676 7522 8732
rect 7458 8672 7522 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 5668 8188 5732 8192
rect 5668 8132 5672 8188
rect 5672 8132 5728 8188
rect 5728 8132 5732 8188
rect 5668 8128 5732 8132
rect 5748 8188 5812 8192
rect 5748 8132 5752 8188
rect 5752 8132 5808 8188
rect 5808 8132 5812 8188
rect 5748 8128 5812 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 8768 8188 8832 8192
rect 8768 8132 8772 8188
rect 8772 8132 8828 8188
rect 8828 8132 8832 8188
rect 8768 8128 8832 8132
rect 8848 8188 8912 8192
rect 8848 8132 8852 8188
rect 8852 8132 8908 8188
rect 8908 8132 8912 8188
rect 8848 8128 8912 8132
rect 8928 8188 8992 8192
rect 8928 8132 8932 8188
rect 8932 8132 8988 8188
rect 8988 8132 8992 8188
rect 8928 8128 8992 8132
rect 9008 8188 9072 8192
rect 9008 8132 9012 8188
rect 9012 8132 9068 8188
rect 9068 8132 9072 8188
rect 9008 8128 9072 8132
rect 4118 7644 4182 7648
rect 4118 7588 4122 7644
rect 4122 7588 4178 7644
rect 4178 7588 4182 7644
rect 4118 7584 4182 7588
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 7218 7644 7282 7648
rect 7218 7588 7222 7644
rect 7222 7588 7278 7644
rect 7278 7588 7282 7644
rect 7218 7584 7282 7588
rect 7298 7644 7362 7648
rect 7298 7588 7302 7644
rect 7302 7588 7358 7644
rect 7358 7588 7362 7644
rect 7298 7584 7362 7588
rect 7378 7644 7442 7648
rect 7378 7588 7382 7644
rect 7382 7588 7438 7644
rect 7438 7588 7442 7644
rect 7378 7584 7442 7588
rect 7458 7644 7522 7648
rect 7458 7588 7462 7644
rect 7462 7588 7518 7644
rect 7518 7588 7522 7644
rect 7458 7584 7522 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 5668 7100 5732 7104
rect 5668 7044 5672 7100
rect 5672 7044 5728 7100
rect 5728 7044 5732 7100
rect 5668 7040 5732 7044
rect 5748 7100 5812 7104
rect 5748 7044 5752 7100
rect 5752 7044 5808 7100
rect 5808 7044 5812 7100
rect 5748 7040 5812 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 8768 7100 8832 7104
rect 8768 7044 8772 7100
rect 8772 7044 8828 7100
rect 8828 7044 8832 7100
rect 8768 7040 8832 7044
rect 8848 7100 8912 7104
rect 8848 7044 8852 7100
rect 8852 7044 8908 7100
rect 8908 7044 8912 7100
rect 8848 7040 8912 7044
rect 8928 7100 8992 7104
rect 8928 7044 8932 7100
rect 8932 7044 8988 7100
rect 8988 7044 8992 7100
rect 8928 7040 8992 7044
rect 9008 7100 9072 7104
rect 9008 7044 9012 7100
rect 9012 7044 9068 7100
rect 9068 7044 9072 7100
rect 9008 7040 9072 7044
rect 4118 6556 4182 6560
rect 4118 6500 4122 6556
rect 4122 6500 4178 6556
rect 4178 6500 4182 6556
rect 4118 6496 4182 6500
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 7218 6556 7282 6560
rect 7218 6500 7222 6556
rect 7222 6500 7278 6556
rect 7278 6500 7282 6556
rect 7218 6496 7282 6500
rect 7298 6556 7362 6560
rect 7298 6500 7302 6556
rect 7302 6500 7358 6556
rect 7358 6500 7362 6556
rect 7298 6496 7362 6500
rect 7378 6556 7442 6560
rect 7378 6500 7382 6556
rect 7382 6500 7438 6556
rect 7438 6500 7442 6556
rect 7378 6496 7442 6500
rect 7458 6556 7522 6560
rect 7458 6500 7462 6556
rect 7462 6500 7518 6556
rect 7518 6500 7522 6556
rect 7458 6496 7522 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 5668 6012 5732 6016
rect 5668 5956 5672 6012
rect 5672 5956 5728 6012
rect 5728 5956 5732 6012
rect 5668 5952 5732 5956
rect 5748 6012 5812 6016
rect 5748 5956 5752 6012
rect 5752 5956 5808 6012
rect 5808 5956 5812 6012
rect 5748 5952 5812 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 8768 6012 8832 6016
rect 8768 5956 8772 6012
rect 8772 5956 8828 6012
rect 8828 5956 8832 6012
rect 8768 5952 8832 5956
rect 8848 6012 8912 6016
rect 8848 5956 8852 6012
rect 8852 5956 8908 6012
rect 8908 5956 8912 6012
rect 8848 5952 8912 5956
rect 8928 6012 8992 6016
rect 8928 5956 8932 6012
rect 8932 5956 8988 6012
rect 8988 5956 8992 6012
rect 8928 5952 8992 5956
rect 9008 6012 9072 6016
rect 9008 5956 9012 6012
rect 9012 5956 9068 6012
rect 9068 5956 9072 6012
rect 9008 5952 9072 5956
rect 4118 5468 4182 5472
rect 4118 5412 4122 5468
rect 4122 5412 4178 5468
rect 4178 5412 4182 5468
rect 4118 5408 4182 5412
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 7218 5468 7282 5472
rect 7218 5412 7222 5468
rect 7222 5412 7278 5468
rect 7278 5412 7282 5468
rect 7218 5408 7282 5412
rect 7298 5468 7362 5472
rect 7298 5412 7302 5468
rect 7302 5412 7358 5468
rect 7358 5412 7362 5468
rect 7298 5408 7362 5412
rect 7378 5468 7442 5472
rect 7378 5412 7382 5468
rect 7382 5412 7438 5468
rect 7438 5412 7442 5468
rect 7378 5408 7442 5412
rect 7458 5468 7522 5472
rect 7458 5412 7462 5468
rect 7462 5412 7518 5468
rect 7518 5412 7522 5468
rect 7458 5408 7522 5412
rect 5668 4924 5732 4928
rect 5668 4868 5672 4924
rect 5672 4868 5728 4924
rect 5728 4868 5732 4924
rect 5668 4864 5732 4868
rect 5748 4924 5812 4928
rect 5748 4868 5752 4924
rect 5752 4868 5808 4924
rect 5808 4868 5812 4924
rect 5748 4864 5812 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 8768 4924 8832 4928
rect 8768 4868 8772 4924
rect 8772 4868 8828 4924
rect 8828 4868 8832 4924
rect 8768 4864 8832 4868
rect 8848 4924 8912 4928
rect 8848 4868 8852 4924
rect 8852 4868 8908 4924
rect 8908 4868 8912 4924
rect 8848 4864 8912 4868
rect 8928 4924 8992 4928
rect 8928 4868 8932 4924
rect 8932 4868 8988 4924
rect 8988 4868 8992 4924
rect 8928 4864 8992 4868
rect 9008 4924 9072 4928
rect 9008 4868 9012 4924
rect 9012 4868 9068 4924
rect 9068 4868 9072 4924
rect 9008 4864 9072 4868
rect 4118 4380 4182 4384
rect 4118 4324 4122 4380
rect 4122 4324 4178 4380
rect 4178 4324 4182 4380
rect 4118 4320 4182 4324
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 7218 4380 7282 4384
rect 7218 4324 7222 4380
rect 7222 4324 7278 4380
rect 7278 4324 7282 4380
rect 7218 4320 7282 4324
rect 7298 4380 7362 4384
rect 7298 4324 7302 4380
rect 7302 4324 7358 4380
rect 7358 4324 7362 4380
rect 7298 4320 7362 4324
rect 7378 4380 7442 4384
rect 7378 4324 7382 4380
rect 7382 4324 7438 4380
rect 7438 4324 7442 4380
rect 7378 4320 7442 4324
rect 7458 4380 7522 4384
rect 7458 4324 7462 4380
rect 7462 4324 7518 4380
rect 7518 4324 7522 4380
rect 7458 4320 7522 4324
rect 4118 3292 4182 3296
rect 4118 3236 4122 3292
rect 4122 3236 4178 3292
rect 4178 3236 4182 3292
rect 4118 3232 4182 3236
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 5668 3836 5732 3840
rect 5668 3780 5672 3836
rect 5672 3780 5728 3836
rect 5728 3780 5732 3836
rect 5668 3776 5732 3780
rect 5748 3836 5812 3840
rect 5748 3780 5752 3836
rect 5752 3780 5808 3836
rect 5808 3780 5812 3836
rect 5748 3776 5812 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 8768 3836 8832 3840
rect 8768 3780 8772 3836
rect 8772 3780 8828 3836
rect 8828 3780 8832 3836
rect 8768 3776 8832 3780
rect 8848 3836 8912 3840
rect 8848 3780 8852 3836
rect 8852 3780 8908 3836
rect 8908 3780 8912 3836
rect 8848 3776 8912 3780
rect 8928 3836 8992 3840
rect 8928 3780 8932 3836
rect 8932 3780 8988 3836
rect 8988 3780 8992 3836
rect 8928 3776 8992 3780
rect 9008 3836 9072 3840
rect 9008 3780 9012 3836
rect 9012 3780 9068 3836
rect 9068 3780 9072 3836
rect 9008 3776 9072 3780
rect 7218 3292 7282 3296
rect 7218 3236 7222 3292
rect 7222 3236 7278 3292
rect 7278 3236 7282 3292
rect 7218 3232 7282 3236
rect 7298 3292 7362 3296
rect 7298 3236 7302 3292
rect 7302 3236 7358 3292
rect 7358 3236 7362 3292
rect 7298 3232 7362 3236
rect 7378 3292 7442 3296
rect 7378 3236 7382 3292
rect 7382 3236 7438 3292
rect 7438 3236 7442 3292
rect 7378 3232 7442 3236
rect 7458 3292 7522 3296
rect 7458 3236 7462 3292
rect 7462 3236 7518 3292
rect 7518 3236 7522 3292
rect 7458 3232 7522 3236
rect 5668 2748 5732 2752
rect 5668 2692 5672 2748
rect 5672 2692 5728 2748
rect 5728 2692 5732 2748
rect 5668 2688 5732 2692
rect 5748 2748 5812 2752
rect 5748 2692 5752 2748
rect 5752 2692 5808 2748
rect 5808 2692 5812 2748
rect 5748 2688 5812 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 8768 2748 8832 2752
rect 8768 2692 8772 2748
rect 8772 2692 8828 2748
rect 8828 2692 8832 2748
rect 8768 2688 8832 2692
rect 8848 2748 8912 2752
rect 8848 2692 8852 2748
rect 8852 2692 8908 2748
rect 8908 2692 8912 2748
rect 8848 2688 8912 2692
rect 8928 2748 8992 2752
rect 8928 2692 8932 2748
rect 8932 2692 8988 2748
rect 8988 2692 8992 2748
rect 8928 2688 8992 2692
rect 9008 2748 9072 2752
rect 9008 2692 9012 2748
rect 9012 2692 9068 2748
rect 9068 2692 9072 2748
rect 9008 2688 9072 2692
rect 4118 2204 4182 2208
rect 4118 2148 4122 2204
rect 4122 2148 4178 2204
rect 4178 2148 4182 2204
rect 4118 2144 4182 2148
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 7218 2204 7282 2208
rect 7218 2148 7222 2204
rect 7222 2148 7278 2204
rect 7278 2148 7282 2204
rect 7218 2144 7282 2148
rect 7298 2204 7362 2208
rect 7298 2148 7302 2204
rect 7302 2148 7358 2204
rect 7358 2148 7362 2204
rect 7298 2144 7362 2148
rect 7378 2204 7442 2208
rect 7378 2148 7382 2204
rect 7382 2148 7438 2204
rect 7438 2148 7442 2204
rect 7378 2144 7442 2148
rect 7458 2204 7522 2208
rect 7458 2148 7462 2204
rect 7462 2148 7518 2204
rect 7518 2148 7522 2204
rect 7458 2144 7522 2148
rect 5668 1660 5732 1664
rect 5668 1604 5672 1660
rect 5672 1604 5728 1660
rect 5728 1604 5732 1660
rect 5668 1600 5732 1604
rect 5748 1660 5812 1664
rect 5748 1604 5752 1660
rect 5752 1604 5808 1660
rect 5808 1604 5812 1660
rect 5748 1600 5812 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 8768 1660 8832 1664
rect 8768 1604 8772 1660
rect 8772 1604 8828 1660
rect 8828 1604 8832 1660
rect 8768 1600 8832 1604
rect 8848 1660 8912 1664
rect 8848 1604 8852 1660
rect 8852 1604 8908 1660
rect 8908 1604 8912 1660
rect 8848 1600 8912 1604
rect 8928 1660 8992 1664
rect 8928 1604 8932 1660
rect 8932 1604 8988 1660
rect 8988 1604 8992 1660
rect 8928 1600 8992 1604
rect 9008 1660 9072 1664
rect 9008 1604 9012 1660
rect 9012 1604 9068 1660
rect 9068 1604 9072 1660
rect 9008 1600 9072 1604
rect 4118 1116 4182 1120
rect 4118 1060 4122 1116
rect 4122 1060 4178 1116
rect 4178 1060 4182 1116
rect 4118 1056 4182 1060
rect 4198 1116 4262 1120
rect 4198 1060 4202 1116
rect 4202 1060 4258 1116
rect 4258 1060 4262 1116
rect 4198 1056 4262 1060
rect 4278 1116 4342 1120
rect 4278 1060 4282 1116
rect 4282 1060 4338 1116
rect 4338 1060 4342 1116
rect 4278 1056 4342 1060
rect 4358 1116 4422 1120
rect 4358 1060 4362 1116
rect 4362 1060 4418 1116
rect 4418 1060 4422 1116
rect 4358 1056 4422 1060
rect 7218 1116 7282 1120
rect 7218 1060 7222 1116
rect 7222 1060 7278 1116
rect 7278 1060 7282 1116
rect 7218 1056 7282 1060
rect 7298 1116 7362 1120
rect 7298 1060 7302 1116
rect 7302 1060 7358 1116
rect 7358 1060 7362 1116
rect 7298 1056 7362 1060
rect 7378 1116 7442 1120
rect 7378 1060 7382 1116
rect 7382 1060 7438 1116
rect 7438 1060 7442 1116
rect 7378 1056 7442 1060
rect 7458 1116 7522 1120
rect 7458 1060 7462 1116
rect 7462 1060 7518 1116
rect 7518 1060 7522 1116
rect 7458 1056 7522 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 4110 10912 4430 11472
rect 5660 11456 5980 11472
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 9908 4430 10848
rect 4110 9824 4152 9908
rect 4388 9824 4430 9908
rect 4110 9760 4118 9824
rect 4422 9760 4430 9824
rect 4110 9672 4152 9760
rect 4388 9672 4430 9760
rect 4110 8736 4430 9672
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 7648 4430 8672
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 6560 4430 7584
rect 4110 6496 4118 6560
rect 4182 6528 4198 6560
rect 4262 6528 4278 6560
rect 4342 6528 4358 6560
rect 4422 6496 4430 6560
rect 4110 6292 4152 6496
rect 4388 6292 4430 6496
rect 4110 5472 4430 6292
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 4384 4430 5408
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 3296 4430 4320
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3148 4430 3232
rect 4110 2912 4152 3148
rect 4388 2912 4430 3148
rect 4110 2208 4430 2912
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 1120 4430 2144
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 5110 10956 5430 11424
rect 5110 10720 5152 10956
rect 5388 10720 5430 10956
rect 5110 7576 5430 10720
rect 5110 7340 5152 7576
rect 5388 7340 5430 7576
rect 5110 4196 5430 7340
rect 5110 3960 5152 4196
rect 5388 3960 5430 4196
rect 5110 1088 5430 3960
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 10368 5980 11392
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 9280 5980 10304
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 8218 5980 9216
rect 5660 8192 5702 8218
rect 5938 8192 5980 8218
rect 5660 8128 5668 8192
rect 5972 8128 5980 8192
rect 5660 7982 5702 8128
rect 5938 7982 5980 8128
rect 5660 7104 5980 7982
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 6016 5980 7040
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 4928 5980 5952
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4838 5980 4864
rect 5660 4602 5702 4838
rect 5938 4602 5980 4838
rect 5660 3840 5980 4602
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 2752 5980 3776
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 1664 5980 2688
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1458 5980 1600
rect 5660 1222 5702 1458
rect 5938 1222 5980 1458
rect 4110 1040 4430 1056
rect 5660 1040 5980 1222
rect 6660 9266 6980 11424
rect 6660 9030 6702 9266
rect 6938 9030 6980 9266
rect 6660 5886 6980 9030
rect 6660 5650 6702 5886
rect 6938 5650 6980 5886
rect 6660 2506 6980 5650
rect 6660 2270 6702 2506
rect 6938 2270 6980 2506
rect 6660 1088 6980 2270
rect 7210 10912 7530 11472
rect 8760 11456 9080 11472
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 9908 7530 10848
rect 7210 9824 7252 9908
rect 7488 9824 7530 9908
rect 7210 9760 7218 9824
rect 7522 9760 7530 9824
rect 7210 9672 7252 9760
rect 7488 9672 7530 9760
rect 7210 8736 7530 9672
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 7648 7530 8672
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 6560 7530 7584
rect 7210 6496 7218 6560
rect 7282 6528 7298 6560
rect 7362 6528 7378 6560
rect 7442 6528 7458 6560
rect 7522 6496 7530 6560
rect 7210 6292 7252 6496
rect 7488 6292 7530 6496
rect 7210 5472 7530 6292
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 4384 7530 5408
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 3296 7530 4320
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 3148 7530 3232
rect 7210 2912 7252 3148
rect 7488 2912 7530 3148
rect 7210 2208 7530 2912
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 1120 7530 2144
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 8210 10956 8530 11424
rect 8210 10720 8252 10956
rect 8488 10720 8530 10956
rect 8210 7576 8530 10720
rect 8210 7340 8252 7576
rect 8488 7340 8530 7576
rect 8210 4196 8530 7340
rect 8210 3960 8252 4196
rect 8488 3960 8530 4196
rect 8210 1088 8530 3960
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 10368 9080 11392
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 9280 9080 10304
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 8218 9080 9216
rect 8760 8192 8802 8218
rect 9038 8192 9080 8218
rect 8760 8128 8768 8192
rect 9072 8128 9080 8192
rect 8760 7982 8802 8128
rect 9038 7982 9080 8128
rect 8760 7104 9080 7982
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 6016 9080 7040
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 4928 9080 5952
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 8760 4838 9080 4864
rect 8760 4602 8802 4838
rect 9038 4602 9080 4838
rect 8760 3840 9080 4602
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 2752 9080 3776
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 1664 9080 2688
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 8760 1458 9080 1600
rect 8760 1222 8802 1458
rect 9038 1222 9080 1458
rect 7210 1040 7530 1056
rect 8760 1040 9080 1222
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 4152 9824 4388 9908
rect 4152 9760 4182 9824
rect 4182 9760 4198 9824
rect 4198 9760 4262 9824
rect 4262 9760 4278 9824
rect 4278 9760 4342 9824
rect 4342 9760 4358 9824
rect 4358 9760 4388 9824
rect 4152 9672 4388 9760
rect 4152 6496 4182 6528
rect 4182 6496 4198 6528
rect 4198 6496 4262 6528
rect 4262 6496 4278 6528
rect 4278 6496 4342 6528
rect 4342 6496 4358 6528
rect 4358 6496 4388 6528
rect 4152 6292 4388 6496
rect 4152 2912 4388 3148
rect 5152 10720 5388 10956
rect 5152 7340 5388 7576
rect 5152 3960 5388 4196
rect 5702 8192 5938 8218
rect 5702 8128 5732 8192
rect 5732 8128 5748 8192
rect 5748 8128 5812 8192
rect 5812 8128 5828 8192
rect 5828 8128 5892 8192
rect 5892 8128 5908 8192
rect 5908 8128 5938 8192
rect 5702 7982 5938 8128
rect 5702 4602 5938 4838
rect 5702 1222 5938 1458
rect 6702 9030 6938 9266
rect 6702 5650 6938 5886
rect 6702 2270 6938 2506
rect 7252 9824 7488 9908
rect 7252 9760 7282 9824
rect 7282 9760 7298 9824
rect 7298 9760 7362 9824
rect 7362 9760 7378 9824
rect 7378 9760 7442 9824
rect 7442 9760 7458 9824
rect 7458 9760 7488 9824
rect 7252 9672 7488 9760
rect 7252 6496 7282 6528
rect 7282 6496 7298 6528
rect 7298 6496 7362 6528
rect 7362 6496 7378 6528
rect 7378 6496 7442 6528
rect 7442 6496 7458 6528
rect 7458 6496 7488 6528
rect 7252 6292 7488 6496
rect 7252 2912 7488 3148
rect 8252 10720 8488 10956
rect 8252 7340 8488 7576
rect 8252 3960 8488 4196
rect 8802 8192 9038 8218
rect 8802 8128 8832 8192
rect 8832 8128 8848 8192
rect 8848 8128 8912 8192
rect 8912 8128 8928 8192
rect 8928 8128 8992 8192
rect 8992 8128 9008 8192
rect 9008 8128 9038 8192
rect 8802 7982 9038 8128
rect 8802 4602 9038 4838
rect 8802 1222 9038 1458
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 5152 10956
rect 5388 10720 8252 10956
rect 8488 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 4152 9908
rect 4388 9672 7252 9908
rect 7488 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 6702 9266
rect 6938 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 5702 8218
rect 5938 7982 8802 8218
rect 9038 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 5152 7576
rect 5388 7340 8252 7576
rect 8488 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 4152 6528
rect 4388 6292 7252 6528
rect 7488 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 6702 5886
rect 6938 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 5702 4838
rect 5938 4602 8802 4838
rect 9038 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 5152 4196
rect 5388 3960 8252 4196
rect 8488 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 4152 3148
rect 4388 2912 7252 3148
rect 7488 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 6702 2506
rect 6938 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 5702 1458
rect 5938 1222 8802 1458
rect 9038 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__clkbuf_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635271187
transform -1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635271187
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635271187
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635271187
transform -1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635271187
transform -1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635271187
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use gpio_logic_high  gpio_logic_high
timestamp 1636130125
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 4600 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1635271187
transform -1 0 4048 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1635271187
transform -1 0 4232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1635271187
transform -1 0 4416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1635271187
transform -1 0 4600 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635271187
transform -1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635271187
transform 1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1635271187
transform -1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1635271187
transform -1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1635271187
transform -1 0 4784 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1635271187
transform -1 0 5336 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1635271187
transform -1 0 5152 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1635271187
transform -1 0 4968 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1635271187
transform -1 0 4784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1635271187
transform -1 0 5520 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5520 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52
timestamp 1635271187
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4784 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635271187
transform -1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635271187
transform -1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1635271187
transform -1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635271187
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635271187
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1635271187
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635271187
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1635271187
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1635271187
transform -1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1635271187
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635271187
transform -1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635271187
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4232 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1635271187
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635271187
transform -1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635271187
transform -1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1635271187
transform -1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1635271187
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1635271187
transform -1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1635271187
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1635271187
transform -1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1635271187
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1635271187
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _208_
timestamp 1635271187
transform 1 0 3588 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1635271187
transform -1 0 6900 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64
timestamp 1635271187
transform 1 0 6808 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_65
timestamp 1635271187
transform 1 0 6900 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1635271187
transform -1 0 8188 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1635271187
transform -1 0 8004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp 1635271187
transform 1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1635271187
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1635271187
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1635271187
transform 1 0 8280 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1635271187
transform -1 0 7912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635271187
transform -1 0 8188 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635271187
transform -1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1635271187
transform 1 0 7084 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _131_
timestamp 1635271187
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1635271187
transform -1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1635271187
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1635271187
transform 1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_63
timestamp 1635271187
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7544 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1635271187
transform 1 0 8280 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1635271187
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1635271187
transform 1 0 6532 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1635271187
transform -1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1635271187
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1635271187
transform -1 0 6716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1635271187
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1635271187
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635271187
transform -1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1635271187
transform 1 0 8832 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1635271187
transform 1 0 8556 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_89
timestamp 1635271187
transform 1 0 9108 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1635271187
transform 1 0 8556 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1635271187
transform 1 0 9476 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1635271187
transform 1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1635271187
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1635271187
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1635271187
transform -1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1635271187
transform 1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1635271187
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1635271187
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1635271187
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635271187
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1635271187
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635271187
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1635271187
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635271187
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1635271187
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635271187
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1635271187
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__5_A
timestamp 1635271187
transform 1 0 1932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1635271187
transform -1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1635271187
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _124_
timestamp 1635271187
transform -1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1635271187
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _107_
timestamp 1635271187
transform -1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 1635271187
transform -1 0 3496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1635271187
transform 1 0 2392 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1635271187
transform -1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1635271187
transform 1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1635271187
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _118_
timestamp 1635271187
transform -1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635271187
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1635271187
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1635271187
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 1635271187
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635271187
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1635271187
transform 1 0 1196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1635271187
transform -1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1635271187
transform 1 0 3680 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1635271187
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1635271187
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1635271187
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1635271187
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1635271187
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1635271187
transform 1 0 5796 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1635271187
transform 1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1635271187
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1635271187
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _145_
timestamp 1635271187
transform -1 0 4140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1635271187
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1635271187
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1635271187
transform -1 0 6072 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1
timestamp 1635271187
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1635271187
transform -1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1635271187
transform 1 0 4968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1635271187
transform 1 0 3588 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1635271187
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1635271187
transform 1 0 6256 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1635271187
transform -1 0 8648 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1635271187
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1635271187
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1635271187
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1635271187
transform -1 0 8648 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1635271187
transform 1 0 6256 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1635271187
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp 1635271187
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1635271187
transform 1 0 6808 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1635271187
transform -1 0 6716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1635271187
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1635271187
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1635271187
transform 1 0 8280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1635271187
transform 1 0 6440 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1635271187
transform 1 0 5980 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1635271187
transform -1 0 9476 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635271187
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1635271187
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635271187
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1635271187
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1635271187
transform -1 0 9476 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1635271187
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635271187
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1635271187
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1635271187
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635271187
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1635271187
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1635271187
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635271187
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1635271187
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _202_
timestamp 1635271187
transform 1 0 2576 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635271187
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1635271187
transform 1 0 1196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1635271187
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1635271187
transform -1 0 3496 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _106__1
timestamp 1635271187
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635271187
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__1_A
timestamp 1635271187
transform -1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1635271187
transform -1 0 2300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1635271187
transform 1 0 2300 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp 1635271187
transform 1 0 1288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635271187
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1635271187
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635271187
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635271187
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1635271187
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__2_A
timestamp 1635271187
transform -1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1635271187
transform -1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1635271187
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1635271187
transform -1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1635271187
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1635271187
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__3
timestamp 1635271187
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1635271187
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1635271187
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _106__2
timestamp 1635271187
transform -1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp 1635271187
transform -1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1635271187
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1635271187
transform -1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1635271187
transform -1 0 3496 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1635271187
transform 1 0 2760 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1635271187
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1635271187
transform -1 0 6072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1635271187
transform -1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1635271187
transform 1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1635271187
transform 1 0 5152 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1635271187
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1635271187
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1635271187
transform 1 0 4140 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1635271187
transform -1 0 5704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1635271187
transform -1 0 6072 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1635271187
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1635271187
transform 1 0 5336 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _151_
timestamp 1635271187
transform -1 0 4140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1635271187
transform 1 0 4876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1635271187
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1635271187
transform -1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8004 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1635271187
transform 1 0 8004 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1635271187
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1635271187
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1635271187
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1635271187
transform 1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1635271187
transform -1 0 9568 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1635271187
transform -1 0 7176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1635271187
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635271187
transform 1 0 5980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7176 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1635271187
transform 1 0 6164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1635271187
transform -1 0 9568 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  _106__4
timestamp 1635271187
transform -1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1635271187
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1635271187
transform 1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1635271187
transform -1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635271187
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1635271187
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1635271187
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1635271187
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635271187
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1635271187
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1635271187
transform 1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1635271187
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635271187
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635271187
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1635271187
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635271187
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1635271187
transform -1 0 3496 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _189_
timestamp 1635271187
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635271187
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__3_A
timestamp 1635271187
transform -1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1635271187
transform -1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1635271187
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1635271187
transform -1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1635271187
transform -1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1635271187
transform -1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1635271187
transform 1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1635271187
transform -1 0 3404 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635271187
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1635271187
transform 1 0 1196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635271187
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1635271187
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1635271187
transform -1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1635271187
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1635271187
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1635271187
transform -1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1635271187
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1635271187
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1635271187
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1635271187
transform 1 0 3680 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1635271187
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1635271187
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1635271187
transform 1 0 3496 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1635271187
transform 1 0 4232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1635271187
transform -1 0 6072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1635271187
transform 1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1635271187
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1635271187
transform 1 0 3404 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1635271187
transform -1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1635271187
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1635271187
transform 1 0 4416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1635271187
transform -1 0 4416 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1635271187
transform 1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1635271187
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1635271187
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1635271187
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1635271187
transform -1 0 7912 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1635271187
transform -1 0 8464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1635271187
transform 1 0 6164 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1635271187
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1635271187
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1635271187
transform -1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1635271187
transform -1 0 8648 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1635271187
transform -1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1635271187
transform -1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1635271187
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1635271187
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp 1635271187
transform 1 0 7176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1635271187
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1635271187
transform 1 0 8740 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1635271187
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__4_A
timestamp 1635271187
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1635271187
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635271187
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _192_
timestamp 1635271187
transform -1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1635271187
transform -1 0 9476 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1635271187
transform 1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1635271187
transform 1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1635271187
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635271187
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635271187
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1635271187
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1635271187
transform -1 0 9568 0 1 10880
box -38 -48 222 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 5660 1040 5980 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 8760 1040 9080 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 6660 1088 6980 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 4110 1040 4430 11472 6 vssd
port 44 nsew ground input
rlabel metal4 s 7210 1040 7530 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 5110 1088 5430 11424 6 vssd1
port 45 nsew ground input
rlabel metal4 s 8210 1088 8530 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
