VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io_alt
  CLASS BLOCK ;
  FOREIGN chip_io_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN mprj_gpio_analog[5]
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_gpio_analog[5]
  PIN mprj_gpio_noesd[5]
    PORT
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
    END
  END mprj_gpio_noesd[5]
  PIN mprj_io_analog_en[12]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in_3v3[12]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
    END
  END mprj_io_in_3v3[12]
  PIN mprj_gpio_analog[6]
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_gpio_analog[6]
  PIN mprj_gpio_noesd[6]
    PORT
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
    END
  END mprj_gpio_noesd[6]
  PIN mprj_io_analog_en[13]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in_3v3[13]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
    END
  END mprj_io_in_3v3[13]
  PIN mprj_io_one[12]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3876.615 3379.435 3876.895 ;
    END
  END mprj_io_one[12]
  PIN mprj_io_one[13]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4322.615 3379.435 4322.895 ;
    END
  END mprj_io_one[13]
  PIN mprj_clamp_high[0]
    ANTENNADIFFAREA 2045.300781 ;
    PORT
      LAYER met2 ;
        RECT 1979.815 5013.660 1982.020 5015.865 ;
    END
  END mprj_clamp_high[0]
  PIN mprj_clamp_low[0]
    ANTENNADIFFAREA 3339.692627 ;
    PORT
      LAYER met2 ;
        RECT 1924.495 4990.055 1925.005 4990.565 ;
    END
  END mprj_clamp_low[0]
  PIN mprj_io_analog_sel[10]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in_3v3[10]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
    END
  END mprj_io_in_3v3[10]
  PIN mprj_gpio_analog[4]
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_gpio_analog[4]
  PIN mprj_gpio_noesd[4]
    PORT
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
    END
  END mprj_gpio_noesd[4]
  PIN mprj_io_analog_en[11]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in_3v3[11]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
    END
  END mprj_io_in_3v3[11]
  PIN mprj_gpio_analog[0]
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_gpio_analog[0]
  PIN mprj_gpio_noesd[0]
    PORT
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
    END
  END mprj_gpio_noesd[0]
  PIN mprj_io_analog_en[7]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in_3v3[7]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
    END
  END mprj_io_in_3v3[7]
  PIN mprj_gpio_analog[1]
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_gpio_analog[1]
  PIN mprj_gpio_noesd[1]
    PORT
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
    END
  END mprj_gpio_noesd[1]
  PIN mprj_io_analog_en[8]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in_3v3[8]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
    END
  END mprj_io_in_3v3[8]
  PIN mprj_gpio_analog[2]
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_gpio_analog[2]
  PIN mprj_gpio_noesd[2]
    PORT
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
    END
  END mprj_gpio_noesd[2]
  PIN mprj_io_analog_en[9]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_in_3v3[9]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
    END
  END mprj_io_in_3v3[9]
  PIN mprj_gpio_analog[3]
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_gpio_analog[3]
  PIN mprj_gpio_noesd[3]
    PORT
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
    END
  END mprj_gpio_noesd[3]
  PIN mprj_io_one[7]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2749.615 3379.435 2749.895 ;
    END
  END mprj_io_one[7]
  PIN mprj_io_one[8]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2975.615 3379.435 2975.895 ;
    END
  END mprj_io_one[8]
  PIN mprj_io_one[9]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3200.615 3379.435 3200.895 ;
    END
  END mprj_io_one[9]
  PIN mprj_io_one[10]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3426.615 3379.435 3426.895 ;
    END
  END mprj_io_one[10]
  PIN mprj_io_one[11]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3651.615 3379.435 3651.895 ;
    END
  END mprj_io_one[11]
  PIN mprj_io_analog_en[10]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_clamp_high[1]
    ANTENNADIFFAREA 2045.300781 ;
    PORT
      LAYER met2 ;
        RECT 1470.815 5013.660 1473.020 5015.865 ;
    END
  END mprj_clamp_high[1]
  PIN mprj_clamp_low[1]
    ANTENNADIFFAREA 3339.692627 ;
    PORT
      LAYER met2 ;
        RECT 1415.495 4990.055 1416.005 4990.565 ;
    END
  END mprj_clamp_low[1]
  PIN mprj_clamp_high[2]
    ANTENNADIFFAREA 2045.300781 ;
    PORT
      LAYER met2 ;
        RECT 1207.815 5013.660 1210.020 5015.865 ;
    END
  END mprj_clamp_high[2]
  PIN mprj_clamp_low[2]
    ANTENNADIFFAREA 3339.692627 ;
    PORT
      LAYER met2 ;
        RECT 1152.495 4990.055 1153.005 4990.565 ;
    END
  END mprj_clamp_low[2]
  PIN mprj_io_slow_sel[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in_3v3[14]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
    END
  END mprj_io_in_3v3[14]
  PIN mprj_gpio_analog[7]
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_gpio_analog[7]
  PIN mprj_gpio_noesd[7]
    PORT
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
    END
  END mprj_gpio_noesd[7]
  PIN mprj_io_ib_mode_sel[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_analog_en[14]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_one[14]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
    END
  END mprj_io_one[14]
  PIN mprj_io_vtrip_sel[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in_3v3[15]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
    END
  END mprj_io_in_3v3[15]
  PIN mprj_gpio_analog[9]
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_gpio_analog[9]
  PIN mprj_gpio_noesd[9]
    PORT
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
    END
  END mprj_gpio_noesd[9]
  PIN mprj_io_analog_en[16]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in_3v3[16]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
    END
  END mprj_io_in_3v3[16]
  PIN mprj_gpio_analog[10]
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_gpio_analog[10]
  PIN mprj_gpio_noesd[10]
    PORT
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
    END
  END mprj_gpio_noesd[10]
  PIN mprj_io_analog_en[17]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in_3v3[17]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
    END
  END mprj_io_in_3v3[17]
  PIN mprj_gpio_analog[8]
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_gpio_analog[8]
  PIN mprj_gpio_noesd[8]
    PORT
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
    END
  END mprj_gpio_noesd[8]
  PIN mprj_io_analog_en[15]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_one[15]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
    END
  END mprj_io_one[15]
  PIN mprj_io_one[16]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
    END
  END mprj_io_one[16]
  PIN mprj_io_one[17]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
    END
  END mprj_io_one[17]
  PIN mprj_gpio_analog[12]
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_gpio_analog[12]
  PIN mprj_gpio_noesd[12]
    PORT
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
    END
  END mprj_gpio_noesd[12]
  PIN mprj_io_analog_en[19]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in_3v3[19]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
    END
  END mprj_io_in_3v3[19]
  PIN mprj_gpio_analog[13]
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_gpio_analog[13]
  PIN mprj_gpio_noesd[13]
    PORT
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
    END
  END mprj_gpio_noesd[13]
  PIN mprj_io_analog_en[20]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in_3v3[20]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
    END
  END mprj_io_in_3v3[20]
  PIN mprj_gpio_analog[11]
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_gpio_analog[11]
  PIN mprj_gpio_noesd[11]
    PORT
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
    END
  END mprj_gpio_noesd[11]
  PIN mprj_io_analog_en[18]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in_3v3[18]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
    END
  END mprj_io_in_3v3[18]
  PIN mprj_io_one[18]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
    END
  END mprj_io_one[18]
  PIN mprj_io_one[19]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
    END
  END mprj_io_one[19]
  PIN mprj_io_one[20]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
    END
  END mprj_io_one[20]
  PIN mprj_gpio_analog[17]
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_gpio_analog[17]
  PIN mprj_gpio_analog[14]
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_gpio_analog[14]
  PIN mprj_gpio_noesd[14]
    PORT
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
    END
  END mprj_gpio_noesd[14]
  PIN mprj_io_analog_en[21]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in_3v3[21]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
    END
  END mprj_io_in_3v3[21]
  PIN mprj_gpio_analog[15]
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_gpio_analog[15]
  PIN mprj_gpio_noesd[15]
    PORT
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
    END
  END mprj_gpio_noesd[15]
  PIN mprj_io_analog_en[22]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in_3v3[22]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
    END
  END mprj_io_in_3v3[22]
  PIN mprj_gpio_analog[16]
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_gpio_analog[16]
  PIN mprj_gpio_noesd[16]
    PORT
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
    END
  END mprj_gpio_noesd[16]
  PIN mprj_io_analog_en[23]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in_3v3[23]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
    END
  END mprj_io_in_3v3[23]
  PIN mprj_io_slow_sel[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_in[24]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_one[21]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
    END
  END mprj_io_one[21]
  PIN mprj_io_one[22]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
    END
  END mprj_io_one[22]
  PIN mprj_io_one[23]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
    END
  END mprj_io_one[23]
  PIN mprj_io_one[24]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
    END
  END mprj_io_one[24]
  PIN mprj_io_ib_mode_sel[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in_3v3[25]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
    END
  END mprj_io_in_3v3[25]
  PIN mprj_io_analog_en[26]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[26]
  PIN resetb_core_h
    ANTENNADIFFAREA 3.024000 ;
    PORT
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
    END
  END resetb_core_h
  PIN mprj_io_analog_en[24]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_in_3v3[26]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
    END
  END mprj_io_in_3v3[26]
  PIN mprj_io_vtrip_sel[24]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN clock_core
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN mprj_io_in_3v3[24]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
    END
  END mprj_io_in_3v3[24]
  PIN mprj_io_analog_en[25]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[76]
  PIN por
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN mprj_io_dm[77]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_gpio_noesd[17]
    PORT
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
    END
  END mprj_gpio_noesd[17]
  PIN mprj_io_holdover[25]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_one[25]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
    END
  END mprj_io_one[25]
  PIN mprj_io_one[26]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 208.565 977.105 210.965 977.385 ;
    END
  END mprj_io_one[26]
  PIN flash_csb_core
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_csb_oeb_core
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 1551.295 195.525 1551.395 195.625 ;
    END
  END flash_csb_oeb_core
  PIN porb_h
    ANTENNAGATEAREA 281.500000 ;
    PORT
      LAYER met2 ;
        RECT 1541.275 208.730 1541.555 211.130 ;
    END
  END porb_h
  PIN mprj_io_analog_en[4]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in_3v3[4]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
    END
  END mprj_io_in_3v3[4]
  PIN mprj_io_analog_en[5]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in_3v3[5]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
    END
  END mprj_io_in_3v3[5]
  PIN mprj_io_analog_en[6]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in_3v3[6]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
    END
  END mprj_io_in_3v3[6]
  PIN mprj_io_one[4]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1412.615 3379.435 1412.895 ;
    END
  END mprj_io_one[4]
  PIN mprj_io_one[5]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1637.615 3379.435 1637.895 ;
    END
  END mprj_io_one[5]
  PIN mprj_io_one[6]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1863.615 3379.435 1863.895 ;
    END
  END mprj_io_one[6]
  PIN flash_io0_oeb_core
    ANTENNAGATEAREA 1.750000 ;
    PORT
      LAYER met2 ;
        RECT 2098.475 208.565 2098.755 210.965 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1_di_core
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER met2 ;
        RECT 2335.215 208.565 2335.495 210.965 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    ANTENNAGATEAREA 1.750000 ;
    PORT
      LAYER met2 ;
        RECT 2372.475 208.565 2372.755 210.965 ;
    END
  END flash_io1_oeb_core
  PIN gpio_in_core
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN flash_clk_oeb_core
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 1825.295 195.525 1825.395 195.625 ;
    END
  END flash_clk_oeb_core
  PIN flash_clk_core
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_io0_di_core
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER met2 ;
        RECT 2061.215 208.565 2061.495 210.965 ;
    END
  END flash_io0_ieb_core
  PIN mprj_io_analog_sel[0]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in_3v3[0]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
    END
  END mprj_io_in_3v3[0]
  PIN mprj_io_dm[9]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN gpio_inenb_core
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_out_core
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN mprj_io_analog_en[1]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_in_3v3[3]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
    END
  END mprj_io_in_3v3[3]
  PIN mprj_io_dm[11]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_vtrip_sel[1]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_one[0]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 510.615 3379.435 510.895 ;
    END
  END mprj_io_one[0]
  PIN mprj_io_one[1]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 736.615 3379.435 736.895 ;
    END
  END mprj_io_one[1]
  PIN mprj_io_one[2]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 961.615 3379.435 961.895 ;
    END
  END mprj_io_one[2]
  PIN mprj_io_one[3]
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1187.615 3379.435 1187.895 ;
    END
  END mprj_io_one[3]
  PIN gpio_outenb_core
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 2647.295 195.525 2647.395 195.625 ;
    END
  END gpio_outenb_core
  PIN mprj_io_analog_en[0]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_in[1]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in_3v3[1]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
    END
  END mprj_io_in_3v3[1]
  PIN mprj_io_analog_en[2]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    ANTENNAGATEAREA 1.529000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in_3v3[2]
    ANTENNADIFFAREA 6.850000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
    END
  END mprj_io_in_3v3[2]
  PIN mprj_io_analog_en[3]
    ANTENNAGATEAREA 0.640000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    ANTENNAGATEAREA 0.500000 ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN gpio_mode1_core
    ANTENNAGATEAREA 1.000000 ;
    PORT
      LAYER met2 ;
        RECT 2624.855 208.730 2625.135 211.130 ;
    END
  END gpio_mode1_core
  PIN vdda
    ANTENNADIFFAREA 4850.636719 ;
    PORT
      LAYER met4 ;
        RECT 192.160 185.065 194.155 187.060 ;
    END
  END vdda
  PIN vdda1
    ANTENNADIFFAREA 11026.780273 ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2299.000 3406.385 2299.960 ;
    END
  END vdda1
  PIN vssa1
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 14070.980469 ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2299.000 3444.735 2374.000 ;
    END
  END vssa1
  PIN vdda2
    ANTENNADIFFAREA 6809.279785 ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2278.995 ;
    END
  END vdda2
  PIN vssa2
    ANTENNAGATEAREA 9.750000 ;
    ANTENNADIFFAREA 7340.723145 ;
    PORT
      LAYER met4 ;
        RECT 143.265 2204.000 143.595 2279.000 ;
    END
  END vssa2
  PIN vccd
    ANTENNAGATEAREA 3801.599854 ;
    ANTENNADIFFAREA 4661.507324 ;
    PORT
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2279.000 ;
    END
  END vccd
  PIN vddio
    ANTENNAGATEAREA 296.339996 ;
    ANTENNADIFFAREA 19164.962891 ;
    PORT
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2279.000 ;
    END
  END vddio
  PIN vssa
    ANTENNAGATEAREA 4.500000 ;
    ANTENNADIFFAREA 7164.618164 ;
    PORT
      LAYER met4 ;
        RECT 176.665 143.595 176.965 143.895 ;
    END
  END vssa
  PIN vssd
    ANTENNAGATEAREA 910.000000 ;
    ANTENNADIFFAREA 9171.701172 ;
    PORT
      LAYER met4 ;
        RECT 663.000 153.765 664.270 158.415 ;
    END
  END vssd
  PIN vssio
    ANTENNAGATEAREA 110.879997 ;
    ANTENNADIFFAREA 36807.734375 ;
    PORT
      LAYER met4 ;
        RECT 0.000 2278.225 24.215 2280.470 ;
    END
  END vssio
  PIN clock
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 936.855 95.440 938.470 97.055 ;
    END
  END clock
  PIN flash_clk
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 1753.855 95.440 1755.470 97.055 ;
    END
  END flash_clk
  PIN flash_csb
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 1479.855 95.440 1481.470 97.055 ;
    END
  END flash_csb
  PIN flash_io0
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 2027.855 95.440 2029.470 97.055 ;
    END
  END flash_io0
  PIN flash_io1
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 2301.855 95.440 2303.470 97.055 ;
    END
  END flash_io1
  PIN gpio
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 2575.855 95.440 2577.470 97.055 ;
    END
  END gpio
  PIN vccd_pad
    ANTENNAGATEAREA 3801.599854 ;
    ANTENNADIFFAREA 4661.507324 ;
    PORT
      LAYER met5 ;
        RECT 99.105 405.265 100.705 406.865 ;
    END
  END vccd_pad
  PIN vdda_pad
    ANTENNADIFFAREA 4850.636719 ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.875 ;
    END
  END vdda_pad
  PIN vddio_pad
    ANTENNAGATEAREA 296.339996 ;
    ANTENNADIFFAREA 19164.962891 ;
    PORT
      LAYER met5 ;
        RECT 95.890 619.465 97.505 621.080 ;
    END
  END vddio_pad
  PIN vddio_pad2
    ANTENNAGATEAREA 296.339996 ;
    ANTENNADIFFAREA 19164.962891 ;
    PORT
      LAYER met5 ;
        RECT 95.890 4417.465 97.505 4419.080 ;
    END
  END vddio_pad2
  PIN vssa_pad
    ANTENNAGATEAREA 4.500000 ;
    ANTENNADIFFAREA 7164.618164 ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.875 ;
    END
  END vssa_pad
  PIN vssd_pad
    ANTENNAGATEAREA 910.000000 ;
    ANTENNADIFFAREA 9171.701172 ;
    PORT
      LAYER met5 ;
        RECT 1271.600 98.770 1273.200 100.370 ;
    END
  END vssd_pad
  PIN vssio_pad
    ANTENNAGATEAREA 110.879997 ;
    ANTENNADIFFAREA 36807.734375 ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.875 ;
    END
  END vssio_pad
  PIN vssio_pad2
    ANTENNAGATEAREA 110.879997 ;
    ANTENNADIFFAREA 36807.734375 ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.940 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 568.735 3492.615 570.200 ;
    END
  END mprj_io[0]
  PIN mprj_io[10]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 3484.735 3492.615 3486.200 ;
    END
  END mprj_io[10]
  PIN mprj_io[11]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 3709.735 3492.615 3711.200 ;
    END
  END mprj_io[11]
  PIN mprj_io[12]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 3934.735 3492.615 3936.200 ;
    END
  END mprj_io[12]
  PIN mprj_io[13]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 4380.735 3492.615 4382.200 ;
    END
  END mprj_io[13]
  PIN mprj_io[1]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 794.735 3492.615 796.200 ;
    END
  END mprj_io[1]
  PIN mprj_io[2]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 1019.735 3492.615 1021.200 ;
    END
  END mprj_io[2]
  PIN mprj_io[3]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 1245.735 3492.615 1247.200 ;
    END
  END mprj_io[3]
  PIN mprj_io[4]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 1470.735 3492.615 1472.200 ;
    END
  END mprj_io[4]
  PIN mprj_io[5]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 1695.735 3492.615 1697.200 ;
    END
  END mprj_io[5]
  PIN mprj_io[6]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 1921.735 3492.615 1923.200 ;
    END
  END mprj_io[6]
  PIN mprj_io[7]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 2807.735 3492.615 2809.200 ;
    END
  END mprj_io[7]
  PIN mprj_io[8]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 3033.735 3492.615 3035.200 ;
    END
  END mprj_io[8]
  PIN mprj_io[9]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 3491.150 3258.735 3492.615 3260.200 ;
    END
  END mprj_io[9]
  PIN mprj_io[25]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 3995.735 33.045 3997.200 ;
    END
  END mprj_io[25]
  PIN mprj_io[35]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 1413.735 33.045 1415.200 ;
    END
  END mprj_io[35]
  PIN mprj_io[36]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 1197.735 33.045 1199.200 ;
    END
  END mprj_io[36]
  PIN mprj_io[37]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 981.735 33.045 983.200 ;
    END
  END mprj_io[37]
  PIN mprj_io[26]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 3779.735 33.045 3781.200 ;
    END
  END mprj_io[26]
  PIN mprj_io[27]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 3563.735 33.045 3565.200 ;
    END
  END mprj_io[27]
  PIN mprj_io[28]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 3347.735 33.045 3349.200 ;
    END
  END mprj_io[28]
  PIN mprj_io[29]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 3131.735 33.045 3133.200 ;
    END
  END mprj_io[29]
  PIN mprj_io[30]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 2915.735 33.045 2917.200 ;
    END
  END mprj_io[30]
  PIN mprj_io[31]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 2699.735 33.045 2701.200 ;
    END
  END mprj_io[31]
  PIN mprj_io[32]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 2061.735 33.045 2063.200 ;
    END
  END mprj_io[32]
  PIN mprj_io[33]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 1845.735 33.045 1847.200 ;
    END
  END mprj_io[33]
  PIN mprj_io[34]
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 31.580 1629.735 33.045 1631.200 ;
    END
  END mprj_io[34]
  PIN resetb
    ANTENNADIFFAREA 398.699982 ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.745 91.545 ;
    END
  END resetb
  PIN mprj_io[15]
    PORT
      LAYER met5 ;
        RECT 3142.050 5093.120 3202.890 5153.940 ;
    END
  END mprj_io[15]
  PIN mprj_io[16]
    PORT
      LAYER met5 ;
        RECT 2633.050 5093.120 2693.890 5153.940 ;
    END
  END mprj_io[16]
  PIN mprj_io[17]
    PORT
      LAYER met5 ;
        RECT 2376.050 5093.120 2436.890 5153.940 ;
    END
  END mprj_io[17]
  PIN mprj_io[14]
    PORT
      LAYER met5 ;
        RECT 3554.690 4826.465 3556.305 4828.080 ;
    END
  END mprj_io[14]
  PIN mprj_io[18]
    PORT
      LAYER met5 ;
        RECT 1931.050 5093.120 1991.890 5153.940 ;
    END
  END mprj_io[18]
  PIN vccd1_pad
    ANTENNADIFFAREA 1391.834717 ;
    PORT
      LAYER met5 ;
        RECT 3557.905 4603.265 3559.505 4604.865 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    ANTENNADIFFAREA 11026.780273 ;
    PORT
      LAYER met5 ;
        RECT 3554.690 4160.465 3556.305 4162.080 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    ANTENNADIFFAREA 11026.780273 ;
    PORT
      LAYER met5 ;
        RECT 3554.690 2587.465 3556.305 2589.080 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 14070.980469 ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.940 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 14070.980469 ;
    PORT
      LAYER met5 ;
        RECT 3554.690 2146.465 3556.305 2148.080 ;
    END
  END vssa1_pad2
  PIN vssd1_pad
    ANTENNADIFFAREA 2860.180176 ;
    PORT
      LAYER met5 ;
        RECT 3557.905 2364.265 3559.505 2365.865 ;
    END
  END vssd1_pad
  PIN mprj_io[21]
    PORT
      LAYER met5 ;
        RECT 907.050 5093.120 967.890 5153.940 ;
    END
  END mprj_io[21]
  PIN mprj_io[22]
    PORT
      LAYER met5 ;
        RECT 650.050 5093.120 710.890 5153.940 ;
    END
  END mprj_io[22]
  PIN mprj_io[23]
    PORT
      LAYER met5 ;
        RECT 393.050 5093.120 453.890 5153.940 ;
    END
  END mprj_io[23]
  PIN mprj_io[24]
    PORT
      LAYER met5 ;
        RECT 95.890 4844.465 97.505 4846.080 ;
    END
  END mprj_io[24]
  PIN mprj_io[19]
    PORT
      LAYER met5 ;
        RECT 1422.050 5093.120 1482.890 5153.940 ;
    END
  END mprj_io[19]
  PIN mprj_io[20]
    PORT
      LAYER met5 ;
        RECT 1159.050 5093.120 1219.890 5153.940 ;
    END
  END mprj_io[20]
  PIN vccd2_pad
    ANTENNADIFFAREA 1391.834717 ;
    PORT
      LAYER met5 ;
        RECT 99.105 4625.265 100.705 4626.865 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    ANTENNADIFFAREA 6809.279785 ;
    PORT
      LAYER met5 ;
        RECT 95.890 2483.465 97.505 2485.080 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    ANTENNAGATEAREA 9.750000 ;
    ANTENNADIFFAREA 7340.723145 ;
    PORT
      LAYER met5 ;
        RECT 95.890 4206.465 97.505 4208.080 ;
    END
  END vssa2_pad
  PIN vssd2_pad
    ANTENNADIFFAREA 2860.180176 ;
    PORT
      LAYER met5 ;
        RECT 99.105 2269.265 100.705 2270.865 ;
    END
  END vssd2_pad
  PIN mprj_analog[1]
    PORT
      LAYER met3 ;
        RECT 3135.455 5061.605 3144.720 5070.870 ;
    END
  END mprj_analog[1]
  PIN mprj_analog[2]
    PORT
      LAYER met3 ;
        RECT 2626.455 5061.605 2635.720 5070.870 ;
    END
  END mprj_analog[2]
  PIN mprj_analog[3]
    PORT
      LAYER met3 ;
        RECT 2369.455 5061.605 2378.720 5070.870 ;
    END
  END mprj_analog[3]
  PIN mprj_analog[0]
    PORT
      LAYER met3 ;
        RECT 3446.605 4808.280 3461.605 4823.280 ;
    END
  END mprj_analog[0]
  PIN mprj_analog[4]
    PORT
      LAYER met3 ;
        RECT 1998.290 5071.775 1999.290 5072.775 ;
    END
  END mprj_analog[4]
  PIN mprj_analog[7]
    PORT
      LAYER met3 ;
        RECT 900.455 5061.605 909.720 5070.870 ;
    END
  END mprj_analog[7]
  PIN mprj_analog[8]
    PORT
      LAYER met3 ;
        RECT 643.455 5061.605 652.720 5070.870 ;
    END
  END mprj_analog[8]
  PIN mprj_analog[9]
    PORT
      LAYER met3 ;
        RECT 386.455 5061.605 395.720 5070.870 ;
    END
  END mprj_analog[9]
  PIN mprj_analog[10]
    PORT
      LAYER met3 ;
        RECT 103.855 4818.520 117.650 4832.315 ;
    END
  END mprj_analog[10]
  PIN mprj_analog[5]
    PORT
      LAYER met3 ;
        RECT 1489.290 5071.775 1490.290 5072.775 ;
    END
  END mprj_analog[5]
  PIN mprj_analog[6]
    PORT
      LAYER met3 ;
        RECT 1226.290 5071.775 1227.290 5072.775 ;
    END
  END mprj_analog[6]
  OBS
      LAYER nwell ;
        RECT 0.000 4628.570 174.795 4630.340 ;
        RECT 0.000 4570.870 1.770 4628.570 ;
        RECT 0.000 4569.100 174.795 4570.870 ;
        RECT 0.000 4417.970 199.315 4419.430 ;
        RECT 0.000 4417.570 171.885 4417.970 ;
        RECT 0.000 4359.695 1.860 4417.570 ;
        RECT 0.000 4357.835 66.985 4359.695 ;
        RECT 0.000 4206.970 199.315 4208.430 ;
        RECT 0.000 4206.570 171.885 4206.970 ;
        RECT 0.000 4148.695 1.860 4206.570 ;
        RECT 0.000 4146.835 66.985 4148.695 ;
        RECT 0.000 4000.330 6.055 4002.000 ;
        RECT 0.000 3990.710 4.055 4000.330 ;
        RECT 0.000 3987.420 3.875 3990.710 ;
        RECT 0.000 3986.685 5.410 3987.420 ;
        RECT 0.000 3981.325 6.025 3986.685 ;
        RECT 0.000 3961.315 6.205 3979.015 ;
        RECT 0.000 3953.355 3.560 3961.315 ;
        RECT 0.000 3937.395 6.245 3953.355 ;
        RECT 0.000 3784.330 6.055 3786.000 ;
        RECT 0.000 3774.710 4.055 3784.330 ;
        RECT 0.000 3771.420 3.875 3774.710 ;
        RECT 0.000 3770.685 5.410 3771.420 ;
        RECT 0.000 3765.325 6.025 3770.685 ;
        RECT 0.000 3745.315 6.205 3763.015 ;
        RECT 0.000 3737.355 3.560 3745.315 ;
        RECT 0.000 3721.395 6.245 3737.355 ;
        RECT 0.000 3568.330 6.055 3570.000 ;
        RECT 0.000 3558.710 4.055 3568.330 ;
        RECT 0.000 3555.420 3.875 3558.710 ;
        RECT 0.000 3554.685 5.410 3555.420 ;
        RECT 0.000 3549.325 6.025 3554.685 ;
        RECT 0.000 3529.315 6.205 3547.015 ;
        RECT 0.000 3521.355 3.560 3529.315 ;
        RECT 0.000 3505.395 6.245 3521.355 ;
        RECT 0.000 3352.330 6.055 3354.000 ;
        RECT 0.000 3342.710 4.055 3352.330 ;
        RECT 0.000 3339.420 3.875 3342.710 ;
        RECT 0.000 3338.685 5.410 3339.420 ;
        RECT 0.000 3333.325 6.025 3338.685 ;
        RECT 0.000 3313.315 6.205 3331.015 ;
        RECT 0.000 3305.355 3.560 3313.315 ;
        RECT 0.000 3289.395 6.245 3305.355 ;
        RECT 0.000 3136.330 6.055 3138.000 ;
        RECT 0.000 3126.710 4.055 3136.330 ;
        RECT 0.000 3123.420 3.875 3126.710 ;
        RECT 0.000 3122.685 5.410 3123.420 ;
        RECT 0.000 3117.325 6.025 3122.685 ;
        RECT 0.000 3097.315 6.205 3115.015 ;
        RECT 0.000 3089.355 3.560 3097.315 ;
        RECT 0.000 3073.395 6.245 3089.355 ;
        RECT 0.000 2920.330 6.055 2922.000 ;
        RECT 0.000 2910.710 4.055 2920.330 ;
        RECT 0.000 2907.420 3.875 2910.710 ;
        RECT 0.000 2906.685 5.410 2907.420 ;
        RECT 0.000 2901.325 6.025 2906.685 ;
        RECT 0.000 2881.315 6.205 2899.015 ;
        RECT 0.000 2873.355 3.560 2881.315 ;
        RECT 0.000 2857.395 6.245 2873.355 ;
        RECT 0.000 2704.330 6.055 2706.000 ;
        RECT 0.000 2694.710 4.055 2704.330 ;
        RECT 0.000 2691.420 3.875 2694.710 ;
        RECT 0.000 2690.685 5.410 2691.420 ;
        RECT 0.000 2685.325 6.025 2690.685 ;
        RECT 0.000 2665.315 6.205 2683.015 ;
        RECT 0.000 2657.355 3.560 2665.315 ;
        RECT 0.000 2641.395 6.245 2657.355 ;
        RECT 0.000 2483.970 199.315 2485.430 ;
        RECT 0.000 2483.570 171.885 2483.970 ;
        RECT 0.000 2425.695 1.860 2483.570 ;
        RECT 0.000 2423.835 66.985 2425.695 ;
        RECT 0.000 2272.570 174.795 2274.340 ;
        RECT 0.000 2214.870 1.770 2272.570 ;
        RECT 0.000 2213.100 174.795 2214.870 ;
        RECT 0.000 2066.330 6.055 2068.000 ;
        RECT 0.000 2056.710 4.055 2066.330 ;
        RECT 0.000 2053.420 3.875 2056.710 ;
        RECT 0.000 2052.685 5.410 2053.420 ;
        RECT 0.000 2047.325 6.025 2052.685 ;
        RECT 0.000 2027.315 6.205 2045.015 ;
        RECT 0.000 2019.355 3.560 2027.315 ;
        RECT 0.000 2003.395 6.245 2019.355 ;
        RECT 0.000 1850.330 6.055 1852.000 ;
        RECT 0.000 1840.710 4.055 1850.330 ;
        RECT 0.000 1837.420 3.875 1840.710 ;
        RECT 0.000 1836.685 5.410 1837.420 ;
        RECT 0.000 1831.325 6.025 1836.685 ;
        RECT 0.000 1811.315 6.205 1829.015 ;
        RECT 0.000 1803.355 3.560 1811.315 ;
        RECT 0.000 1787.395 6.245 1803.355 ;
        RECT 0.000 1634.330 6.055 1636.000 ;
        RECT 0.000 1624.710 4.055 1634.330 ;
        RECT 0.000 1621.420 3.875 1624.710 ;
        RECT 0.000 1620.685 5.410 1621.420 ;
        RECT 0.000 1615.325 6.025 1620.685 ;
        RECT 0.000 1595.315 6.205 1613.015 ;
        RECT 0.000 1587.355 3.560 1595.315 ;
        RECT 0.000 1571.395 6.245 1587.355 ;
        RECT 0.000 1418.330 6.055 1420.000 ;
        RECT 0.000 1408.710 4.055 1418.330 ;
        RECT 0.000 1405.420 3.875 1408.710 ;
        RECT 0.000 1404.685 5.410 1405.420 ;
        RECT 0.000 1399.325 6.025 1404.685 ;
        RECT 0.000 1379.315 6.205 1397.015 ;
        RECT 0.000 1371.355 3.560 1379.315 ;
        RECT 0.000 1355.395 6.245 1371.355 ;
        RECT 0.000 1202.330 6.055 1204.000 ;
        RECT 0.000 1192.710 4.055 1202.330 ;
        RECT 0.000 1189.420 3.875 1192.710 ;
        RECT 0.000 1188.685 5.410 1189.420 ;
        RECT 0.000 1183.325 6.025 1188.685 ;
        RECT 0.000 1163.315 6.205 1181.015 ;
        RECT 0.000 1155.355 3.560 1163.315 ;
        RECT 0.000 1139.395 6.245 1155.355 ;
        RECT 0.000 986.330 6.055 988.000 ;
        RECT 0.000 976.710 4.055 986.330 ;
        RECT 0.000 973.420 3.875 976.710 ;
        RECT 0.000 972.685 5.410 973.420 ;
        RECT 0.000 967.325 6.025 972.685 ;
        RECT 0.000 947.315 6.205 965.015 ;
        RECT 0.000 939.355 3.560 947.315 ;
        RECT 0.000 923.395 6.245 939.355 ;
        RECT 0.000 619.970 199.315 621.430 ;
        RECT 0.000 619.570 171.885 619.970 ;
        RECT 0.000 561.695 1.860 619.570 ;
        RECT 0.000 559.835 66.985 561.695 ;
        RECT 0.000 408.570 174.795 410.340 ;
        RECT 0.000 350.870 1.770 408.570 ;
        RECT 0.000 349.100 174.795 350.870 ;
      LAYER li1 ;
        RECT 0.220 0.220 3587.780 5187.695 ;
      LAYER met1 ;
        RECT 0.000 0.000 3588.000 5187.725 ;
      LAYER met2 ;
        RECT 0.000 5016.145 3588.000 5183.075 ;
        RECT 0.000 5013.380 1207.535 5016.145 ;
        RECT 1210.300 5013.380 1470.535 5016.145 ;
        RECT 1473.300 5013.380 1979.535 5016.145 ;
        RECT 1982.300 5013.380 3588.000 5016.145 ;
        RECT 0.000 4990.845 3588.000 5013.380 ;
        RECT 0.000 4989.775 1152.215 4990.845 ;
        RECT 1153.285 4989.775 1415.215 4990.845 ;
        RECT 1416.285 4989.775 1924.215 4990.845 ;
        RECT 1925.285 4989.775 3588.000 4990.845 ;
        RECT 0.000 4390.795 3588.000 4989.775 ;
        RECT 0.000 4389.955 3376.755 4390.795 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 0.000 4388.035 3588.000 4389.955 ;
        RECT 0.000 4387.195 3376.755 4388.035 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 0.000 4384.815 3588.000 4387.195 ;
        RECT 0.000 4383.975 3376.755 4384.815 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 0.000 4381.595 3588.000 4383.975 ;
        RECT 0.000 4380.755 3376.755 4381.595 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
        RECT 0.000 4372.395 3588.000 4380.755 ;
        RECT 0.000 4371.555 3376.755 4372.395 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 0.000 4369.635 3588.000 4371.555 ;
        RECT 0.000 4368.795 3376.755 4369.635 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 0.000 4366.415 3588.000 4368.795 ;
        RECT 0.000 4365.575 3376.755 4366.415 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 0.000 4363.195 3588.000 4365.575 ;
        RECT 0.000 4362.355 3376.755 4363.195 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
        RECT 0.000 4350.775 3588.000 4362.355 ;
        RECT 0.000 4349.935 3376.755 4350.775 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 0.000 4348.015 3588.000 4349.935 ;
        RECT 0.000 4347.175 3376.755 4348.015 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 0.000 4344.795 3588.000 4347.175 ;
        RECT 0.000 4343.955 3376.755 4344.795 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 0.000 4341.575 3588.000 4343.955 ;
        RECT 0.000 4340.735 3376.755 4341.575 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 0.000 4338.815 3588.000 4340.735 ;
        RECT 0.000 4337.975 3376.755 4338.815 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 0.000 4335.595 3588.000 4337.975 ;
        RECT 0.000 4334.755 3376.755 4335.595 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 0.000 4329.615 3588.000 4334.755 ;
        RECT 0.000 4328.775 3376.755 4329.615 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 0.000 4326.395 3588.000 4328.775 ;
        RECT 0.000 4325.555 3376.755 4326.395 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 0.000 4323.175 3588.000 4325.555 ;
        RECT 0.000 4322.335 3376.755 4323.175 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
        RECT 0.000 4317.195 3588.000 4322.335 ;
        RECT 0.000 4316.355 3376.755 4317.195 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
        RECT 0.000 3997.645 3588.000 4316.355 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 211.245 3996.805 3588.000 3997.645 ;
        RECT 0.000 3991.665 3588.000 3996.805 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
        RECT 211.245 3990.825 3588.000 3991.665 ;
        RECT 0.000 3988.445 3588.000 3990.825 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 211.245 3987.605 3588.000 3988.445 ;
        RECT 0.000 3985.225 3588.000 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 211.245 3984.385 3588.000 3985.225 ;
        RECT 0.000 3979.245 3588.000 3984.385 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 211.245 3978.405 3588.000 3979.245 ;
        RECT 0.000 3976.025 3588.000 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
        RECT 211.245 3975.185 3588.000 3976.025 ;
        RECT 0.000 3973.265 3588.000 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 211.245 3972.425 3588.000 3973.265 ;
        RECT 0.000 3970.045 3588.000 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 211.245 3969.205 3588.000 3970.045 ;
        RECT 0.000 3966.825 3588.000 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 211.245 3965.985 3588.000 3966.825 ;
        RECT 0.000 3964.065 3588.000 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 211.245 3963.225 3588.000 3964.065 ;
        RECT 0.000 3951.645 3588.000 3963.225 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 211.245 3950.805 3588.000 3951.645 ;
        RECT 0.000 3948.425 3588.000 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 211.245 3947.585 3588.000 3948.425 ;
        RECT 0.000 3945.205 3588.000 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 211.245 3944.795 3588.000 3945.205 ;
        RECT 211.245 3944.365 3376.755 3944.795 ;
        RECT 0.000 3943.955 3376.755 3944.365 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 0.000 3942.445 3588.000 3943.955 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
        RECT 211.245 3942.035 3588.000 3942.445 ;
        RECT 211.245 3941.605 3376.755 3942.035 ;
        RECT 0.000 3941.195 3376.755 3941.605 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 0.000 3938.815 3588.000 3941.195 ;
        RECT 0.000 3937.975 3376.755 3938.815 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 0.000 3935.595 3588.000 3937.975 ;
        RECT 0.000 3934.755 3376.755 3935.595 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
        RECT 0.000 3933.245 3588.000 3934.755 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
        RECT 211.245 3932.405 3588.000 3933.245 ;
        RECT 0.000 3930.025 3588.000 3932.405 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 211.245 3929.185 3588.000 3930.025 ;
        RECT 0.000 3926.805 3588.000 3929.185 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 211.245 3926.395 3588.000 3926.805 ;
        RECT 211.245 3925.965 3376.755 3926.395 ;
        RECT 0.000 3925.555 3376.755 3925.965 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 0.000 3924.045 3588.000 3925.555 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
        RECT 211.245 3923.635 3588.000 3924.045 ;
        RECT 211.245 3923.205 3376.755 3923.635 ;
        RECT 0.000 3922.795 3376.755 3923.205 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 0.000 3920.415 3588.000 3922.795 ;
        RECT 0.000 3919.575 3376.755 3920.415 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 0.000 3917.195 3588.000 3919.575 ;
        RECT 0.000 3916.355 3376.755 3917.195 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
        RECT 0.000 3904.775 3588.000 3916.355 ;
        RECT 0.000 3903.935 3376.755 3904.775 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 0.000 3902.015 3588.000 3903.935 ;
        RECT 0.000 3901.175 3376.755 3902.015 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 0.000 3898.795 3588.000 3901.175 ;
        RECT 0.000 3897.955 3376.755 3898.795 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 0.000 3895.575 3588.000 3897.955 ;
        RECT 0.000 3894.735 3376.755 3895.575 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 0.000 3892.815 3588.000 3894.735 ;
        RECT 0.000 3891.975 3376.755 3892.815 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 0.000 3889.595 3588.000 3891.975 ;
        RECT 0.000 3888.755 3376.755 3889.595 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 0.000 3883.615 3588.000 3888.755 ;
        RECT 0.000 3882.775 3376.755 3883.615 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 0.000 3880.395 3588.000 3882.775 ;
        RECT 0.000 3879.555 3376.755 3880.395 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
        RECT 0.000 3877.175 3588.000 3879.555 ;
        RECT 0.000 3876.335 3376.755 3877.175 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
        RECT 0.000 3871.195 3588.000 3876.335 ;
        RECT 0.000 3870.355 3376.755 3871.195 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
        RECT 0.000 3781.645 3588.000 3870.355 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 211.245 3780.805 3588.000 3781.645 ;
        RECT 0.000 3775.665 3588.000 3780.805 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
        RECT 211.245 3774.825 3588.000 3775.665 ;
        RECT 0.000 3772.445 3588.000 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 211.245 3771.605 3588.000 3772.445 ;
        RECT 0.000 3769.225 3588.000 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 211.245 3768.385 3588.000 3769.225 ;
        RECT 0.000 3763.245 3588.000 3768.385 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 211.245 3762.405 3588.000 3763.245 ;
        RECT 0.000 3760.025 3588.000 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
        RECT 211.245 3759.185 3588.000 3760.025 ;
        RECT 0.000 3757.265 3588.000 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 211.245 3756.425 3588.000 3757.265 ;
        RECT 0.000 3754.045 3588.000 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 211.245 3753.205 3588.000 3754.045 ;
        RECT 0.000 3750.825 3588.000 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 211.245 3749.985 3588.000 3750.825 ;
        RECT 0.000 3748.065 3588.000 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 211.245 3747.225 3588.000 3748.065 ;
        RECT 0.000 3735.645 3588.000 3747.225 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
        RECT 211.245 3734.805 3588.000 3735.645 ;
        RECT 0.000 3732.425 3588.000 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 211.245 3731.585 3588.000 3732.425 ;
        RECT 0.000 3729.205 3588.000 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 211.245 3728.365 3588.000 3729.205 ;
        RECT 0.000 3726.445 3588.000 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 211.245 3725.605 3588.000 3726.445 ;
        RECT 0.000 3719.795 3588.000 3725.605 ;
        RECT 0.000 3718.955 3376.755 3719.795 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 0.000 3717.245 3588.000 3718.955 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 211.245 3717.035 3588.000 3717.245 ;
        RECT 211.245 3716.405 3376.755 3717.035 ;
        RECT 0.000 3716.195 3376.755 3716.405 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 0.000 3714.025 3588.000 3716.195 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 211.245 3713.815 3588.000 3714.025 ;
        RECT 211.245 3713.185 3376.755 3713.815 ;
        RECT 0.000 3712.975 3376.755 3713.185 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 0.000 3710.805 3588.000 3712.975 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 211.245 3710.595 3588.000 3710.805 ;
        RECT 211.245 3709.965 3376.755 3710.595 ;
        RECT 0.000 3709.755 3376.755 3709.965 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 0.000 3708.045 3588.000 3709.755 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
        RECT 211.245 3707.205 3588.000 3708.045 ;
        RECT 0.000 3701.395 3588.000 3707.205 ;
        RECT 0.000 3700.555 3376.755 3701.395 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 0.000 3698.635 3588.000 3700.555 ;
        RECT 0.000 3697.795 3376.755 3698.635 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 0.000 3695.415 3588.000 3697.795 ;
        RECT 0.000 3694.575 3376.755 3695.415 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 0.000 3692.195 3588.000 3694.575 ;
        RECT 0.000 3691.355 3376.755 3692.195 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
        RECT 0.000 3679.775 3588.000 3691.355 ;
        RECT 0.000 3678.935 3376.755 3679.775 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 0.000 3677.015 3588.000 3678.935 ;
        RECT 0.000 3676.175 3376.755 3677.015 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 0.000 3673.795 3588.000 3676.175 ;
        RECT 0.000 3672.955 3376.755 3673.795 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 0.000 3670.575 3588.000 3672.955 ;
        RECT 0.000 3669.735 3376.755 3670.575 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 0.000 3667.815 3588.000 3669.735 ;
        RECT 0.000 3666.975 3376.755 3667.815 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 0.000 3664.595 3588.000 3666.975 ;
        RECT 0.000 3663.755 3376.755 3664.595 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 0.000 3658.615 3588.000 3663.755 ;
        RECT 0.000 3657.775 3376.755 3658.615 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 0.000 3655.395 3588.000 3657.775 ;
        RECT 0.000 3654.555 3376.755 3655.395 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
        RECT 0.000 3652.175 3588.000 3654.555 ;
        RECT 0.000 3651.335 3376.755 3652.175 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
        RECT 0.000 3646.195 3588.000 3651.335 ;
        RECT 0.000 3645.355 3376.755 3646.195 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
        RECT 0.000 3565.645 3588.000 3645.355 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
        RECT 211.245 3564.805 3588.000 3565.645 ;
        RECT 0.000 3559.665 3588.000 3564.805 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
        RECT 211.245 3558.825 3588.000 3559.665 ;
        RECT 0.000 3556.445 3588.000 3558.825 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 211.245 3555.605 3588.000 3556.445 ;
        RECT 0.000 3553.225 3588.000 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 211.245 3552.385 3588.000 3553.225 ;
        RECT 0.000 3547.245 3588.000 3552.385 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 211.245 3546.405 3588.000 3547.245 ;
        RECT 0.000 3544.025 3588.000 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
        RECT 211.245 3543.185 3588.000 3544.025 ;
        RECT 0.000 3541.265 3588.000 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 211.245 3540.425 3588.000 3541.265 ;
        RECT 0.000 3538.045 3588.000 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 211.245 3537.205 3588.000 3538.045 ;
        RECT 0.000 3534.825 3588.000 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 211.245 3533.985 3588.000 3534.825 ;
        RECT 0.000 3532.065 3588.000 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
        RECT 211.245 3531.225 3588.000 3532.065 ;
        RECT 0.000 3519.645 3588.000 3531.225 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 211.245 3518.805 3588.000 3519.645 ;
        RECT 0.000 3516.425 3588.000 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 211.245 3515.585 3588.000 3516.425 ;
        RECT 0.000 3513.205 3588.000 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 211.245 3512.365 3588.000 3513.205 ;
        RECT 0.000 3510.445 3588.000 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 211.245 3509.605 3588.000 3510.445 ;
        RECT 0.000 3501.245 3588.000 3509.605 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 211.245 3500.405 3588.000 3501.245 ;
        RECT 0.000 3498.025 3588.000 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 211.245 3497.185 3588.000 3498.025 ;
        RECT 0.000 3494.805 3588.000 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 211.245 3494.795 3588.000 3494.805 ;
        RECT 211.245 3493.965 3376.755 3494.795 ;
        RECT 0.000 3493.955 3376.755 3493.965 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 0.000 3492.045 3588.000 3493.955 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
        RECT 211.245 3492.035 3588.000 3492.045 ;
        RECT 211.245 3491.205 3376.755 3492.035 ;
        RECT 0.000 3491.195 3376.755 3491.205 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 0.000 3488.815 3588.000 3491.195 ;
        RECT 0.000 3487.975 3376.755 3488.815 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 0.000 3485.595 3588.000 3487.975 ;
        RECT 0.000 3484.755 3376.755 3485.595 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
        RECT 0.000 3476.395 3588.000 3484.755 ;
        RECT 0.000 3475.555 3376.755 3476.395 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 0.000 3473.635 3588.000 3475.555 ;
        RECT 0.000 3472.795 3376.755 3473.635 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 0.000 3470.415 3588.000 3472.795 ;
        RECT 0.000 3469.575 3376.755 3470.415 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 0.000 3467.195 3588.000 3469.575 ;
        RECT 0.000 3466.355 3376.755 3467.195 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
        RECT 0.000 3454.775 3588.000 3466.355 ;
        RECT 0.000 3453.935 3376.755 3454.775 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 0.000 3452.015 3588.000 3453.935 ;
        RECT 0.000 3451.175 3376.755 3452.015 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 0.000 3448.795 3588.000 3451.175 ;
        RECT 0.000 3447.955 3376.755 3448.795 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 0.000 3445.575 3588.000 3447.955 ;
        RECT 0.000 3444.735 3376.755 3445.575 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 0.000 3442.815 3588.000 3444.735 ;
        RECT 0.000 3441.975 3376.755 3442.815 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 0.000 3439.595 3588.000 3441.975 ;
        RECT 0.000 3438.755 3376.755 3439.595 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 0.000 3433.615 3588.000 3438.755 ;
        RECT 0.000 3432.775 3376.755 3433.615 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 0.000 3430.395 3588.000 3432.775 ;
        RECT 0.000 3429.555 3376.755 3430.395 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 0.000 3427.175 3588.000 3429.555 ;
        RECT 0.000 3426.335 3376.755 3427.175 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
        RECT 0.000 3421.195 3588.000 3426.335 ;
        RECT 0.000 3420.355 3376.755 3421.195 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
        RECT 0.000 3349.645 3588.000 3420.355 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 211.245 3348.805 3588.000 3349.645 ;
        RECT 0.000 3343.665 3588.000 3348.805 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
        RECT 211.245 3342.825 3588.000 3343.665 ;
        RECT 0.000 3340.445 3588.000 3342.825 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 211.245 3339.605 3588.000 3340.445 ;
        RECT 0.000 3337.225 3588.000 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 211.245 3336.385 3588.000 3337.225 ;
        RECT 0.000 3331.245 3588.000 3336.385 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 211.245 3330.405 3588.000 3331.245 ;
        RECT 0.000 3328.025 3588.000 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
        RECT 211.245 3327.185 3588.000 3328.025 ;
        RECT 0.000 3325.265 3588.000 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 211.245 3324.425 3588.000 3325.265 ;
        RECT 0.000 3322.045 3588.000 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 211.245 3321.205 3588.000 3322.045 ;
        RECT 0.000 3318.825 3588.000 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 211.245 3317.985 3588.000 3318.825 ;
        RECT 0.000 3316.065 3588.000 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
        RECT 211.245 3315.225 3588.000 3316.065 ;
        RECT 0.000 3303.645 3588.000 3315.225 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 211.245 3302.805 3588.000 3303.645 ;
        RECT 0.000 3300.425 3588.000 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 211.245 3299.585 3588.000 3300.425 ;
        RECT 0.000 3297.205 3588.000 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 211.245 3296.365 3588.000 3297.205 ;
        RECT 0.000 3294.445 3588.000 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 211.245 3293.605 3588.000 3294.445 ;
        RECT 0.000 3285.245 3588.000 3293.605 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 211.245 3284.405 3588.000 3285.245 ;
        RECT 0.000 3282.025 3588.000 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 211.245 3281.185 3588.000 3282.025 ;
        RECT 0.000 3278.805 3588.000 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 211.245 3277.965 3588.000 3278.805 ;
        RECT 0.000 3276.045 3588.000 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
        RECT 211.245 3275.205 3588.000 3276.045 ;
        RECT 0.000 3268.795 3588.000 3275.205 ;
        RECT 0.000 3267.955 3376.755 3268.795 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 0.000 3266.035 3588.000 3267.955 ;
        RECT 0.000 3265.195 3376.755 3266.035 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 0.000 3262.815 3588.000 3265.195 ;
        RECT 0.000 3261.975 3376.755 3262.815 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 0.000 3259.595 3588.000 3261.975 ;
        RECT 0.000 3258.755 3376.755 3259.595 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
        RECT 0.000 3250.395 3588.000 3258.755 ;
        RECT 0.000 3249.555 3376.755 3250.395 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 0.000 3247.635 3588.000 3249.555 ;
        RECT 0.000 3246.795 3376.755 3247.635 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 0.000 3244.415 3588.000 3246.795 ;
        RECT 0.000 3243.575 3376.755 3244.415 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 0.000 3241.195 3588.000 3243.575 ;
        RECT 0.000 3240.355 3376.755 3241.195 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
        RECT 0.000 3228.775 3588.000 3240.355 ;
        RECT 0.000 3227.935 3376.755 3228.775 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 0.000 3226.015 3588.000 3227.935 ;
        RECT 0.000 3225.175 3376.755 3226.015 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 0.000 3222.795 3588.000 3225.175 ;
        RECT 0.000 3221.955 3376.755 3222.795 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 0.000 3219.575 3588.000 3221.955 ;
        RECT 0.000 3218.735 3376.755 3219.575 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 0.000 3216.815 3588.000 3218.735 ;
        RECT 0.000 3215.975 3376.755 3216.815 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 0.000 3213.595 3588.000 3215.975 ;
        RECT 0.000 3212.755 3376.755 3213.595 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 0.000 3207.615 3588.000 3212.755 ;
        RECT 0.000 3206.775 3376.755 3207.615 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 0.000 3204.395 3588.000 3206.775 ;
        RECT 0.000 3203.555 3376.755 3204.395 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
        RECT 0.000 3201.175 3588.000 3203.555 ;
        RECT 0.000 3200.335 3376.755 3201.175 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
        RECT 0.000 3195.195 3588.000 3200.335 ;
        RECT 0.000 3194.355 3376.755 3195.195 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
        RECT 0.000 3133.645 3588.000 3194.355 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 211.245 3132.805 3588.000 3133.645 ;
        RECT 0.000 3127.665 3588.000 3132.805 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
        RECT 211.245 3126.825 3588.000 3127.665 ;
        RECT 0.000 3124.445 3588.000 3126.825 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 211.245 3123.605 3588.000 3124.445 ;
        RECT 0.000 3121.225 3588.000 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 211.245 3120.385 3588.000 3121.225 ;
        RECT 0.000 3115.245 3588.000 3120.385 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 211.245 3114.405 3588.000 3115.245 ;
        RECT 0.000 3112.025 3588.000 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
        RECT 211.245 3111.185 3588.000 3112.025 ;
        RECT 0.000 3109.265 3588.000 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 211.245 3108.425 3588.000 3109.265 ;
        RECT 0.000 3106.045 3588.000 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 211.245 3105.205 3588.000 3106.045 ;
        RECT 0.000 3102.825 3588.000 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 211.245 3101.985 3588.000 3102.825 ;
        RECT 0.000 3100.065 3588.000 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 211.245 3099.225 3588.000 3100.065 ;
        RECT 0.000 3087.645 3588.000 3099.225 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 211.245 3086.805 3588.000 3087.645 ;
        RECT 0.000 3084.425 3588.000 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 211.245 3083.585 3588.000 3084.425 ;
        RECT 0.000 3081.205 3588.000 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 211.245 3080.365 3588.000 3081.205 ;
        RECT 0.000 3078.445 3588.000 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 211.245 3077.605 3588.000 3078.445 ;
        RECT 0.000 3069.245 3588.000 3077.605 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 211.245 3068.405 3588.000 3069.245 ;
        RECT 0.000 3066.025 3588.000 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 211.245 3065.185 3588.000 3066.025 ;
        RECT 0.000 3062.805 3588.000 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 211.245 3061.965 3588.000 3062.805 ;
        RECT 0.000 3060.045 3588.000 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
        RECT 211.245 3059.205 3588.000 3060.045 ;
        RECT 0.000 3043.795 3588.000 3059.205 ;
        RECT 0.000 3042.955 3376.755 3043.795 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 0.000 3041.035 3588.000 3042.955 ;
        RECT 0.000 3040.195 3376.755 3041.035 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 0.000 3037.815 3588.000 3040.195 ;
        RECT 0.000 3036.975 3376.755 3037.815 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 0.000 3034.595 3588.000 3036.975 ;
        RECT 0.000 3033.755 3376.755 3034.595 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
        RECT 0.000 3025.395 3588.000 3033.755 ;
        RECT 0.000 3024.555 3376.755 3025.395 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 0.000 3022.635 3588.000 3024.555 ;
        RECT 0.000 3021.795 3376.755 3022.635 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 0.000 3019.415 3588.000 3021.795 ;
        RECT 0.000 3018.575 3376.755 3019.415 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 0.000 3016.195 3588.000 3018.575 ;
        RECT 0.000 3015.355 3376.755 3016.195 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
        RECT 0.000 3003.775 3588.000 3015.355 ;
        RECT 0.000 3002.935 3376.755 3003.775 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 0.000 3001.015 3588.000 3002.935 ;
        RECT 0.000 3000.175 3376.755 3001.015 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 0.000 2997.795 3588.000 3000.175 ;
        RECT 0.000 2996.955 3376.755 2997.795 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 0.000 2994.575 3588.000 2996.955 ;
        RECT 0.000 2993.735 3376.755 2994.575 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 0.000 2991.815 3588.000 2993.735 ;
        RECT 0.000 2990.975 3376.755 2991.815 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 0.000 2988.595 3588.000 2990.975 ;
        RECT 0.000 2987.755 3376.755 2988.595 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 0.000 2982.615 3588.000 2987.755 ;
        RECT 0.000 2981.775 3376.755 2982.615 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 0.000 2979.395 3588.000 2981.775 ;
        RECT 0.000 2978.555 3376.755 2979.395 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 0.000 2976.175 3588.000 2978.555 ;
        RECT 0.000 2975.335 3376.755 2976.175 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
        RECT 0.000 2970.195 3588.000 2975.335 ;
        RECT 0.000 2969.355 3376.755 2970.195 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
        RECT 0.000 2917.645 3588.000 2969.355 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
        RECT 211.245 2916.805 3588.000 2917.645 ;
        RECT 0.000 2911.665 3588.000 2916.805 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
        RECT 211.245 2910.825 3588.000 2911.665 ;
        RECT 0.000 2908.445 3588.000 2910.825 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
        RECT 211.245 2907.605 3588.000 2908.445 ;
        RECT 0.000 2905.225 3588.000 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 211.245 2904.385 3588.000 2905.225 ;
        RECT 0.000 2899.245 3588.000 2904.385 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 211.245 2898.405 3588.000 2899.245 ;
        RECT 0.000 2896.025 3588.000 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
        RECT 211.245 2895.185 3588.000 2896.025 ;
        RECT 0.000 2893.265 3588.000 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 211.245 2892.425 3588.000 2893.265 ;
        RECT 0.000 2890.045 3588.000 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 211.245 2889.205 3588.000 2890.045 ;
        RECT 0.000 2886.825 3588.000 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 211.245 2885.985 3588.000 2886.825 ;
        RECT 0.000 2884.065 3588.000 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 211.245 2883.225 3588.000 2884.065 ;
        RECT 0.000 2871.645 3588.000 2883.225 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 211.245 2870.805 3588.000 2871.645 ;
        RECT 0.000 2868.425 3588.000 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 211.245 2867.585 3588.000 2868.425 ;
        RECT 0.000 2865.205 3588.000 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 211.245 2864.365 3588.000 2865.205 ;
        RECT 0.000 2862.445 3588.000 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 211.245 2861.605 3588.000 2862.445 ;
        RECT 0.000 2853.245 3588.000 2861.605 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 211.245 2852.405 3588.000 2853.245 ;
        RECT 0.000 2850.025 3588.000 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 211.245 2849.185 3588.000 2850.025 ;
        RECT 0.000 2846.805 3588.000 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 211.245 2845.965 3588.000 2846.805 ;
        RECT 0.000 2844.045 3588.000 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
        RECT 211.245 2843.205 3588.000 2844.045 ;
        RECT 0.000 2817.795 3588.000 2843.205 ;
        RECT 0.000 2816.955 3376.755 2817.795 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 0.000 2815.035 3588.000 2816.955 ;
        RECT 0.000 2814.195 3376.755 2815.035 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 0.000 2811.815 3588.000 2814.195 ;
        RECT 0.000 2810.975 3376.755 2811.815 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 0.000 2808.595 3588.000 2810.975 ;
        RECT 0.000 2807.755 3376.755 2808.595 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
        RECT 0.000 2799.395 3588.000 2807.755 ;
        RECT 0.000 2798.555 3376.755 2799.395 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 0.000 2796.635 3588.000 2798.555 ;
        RECT 0.000 2795.795 3376.755 2796.635 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 0.000 2793.415 3588.000 2795.795 ;
        RECT 0.000 2792.575 3376.755 2793.415 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 0.000 2790.195 3588.000 2792.575 ;
        RECT 0.000 2789.355 3376.755 2790.195 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
        RECT 0.000 2777.775 3588.000 2789.355 ;
        RECT 0.000 2776.935 3376.755 2777.775 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 0.000 2775.015 3588.000 2776.935 ;
        RECT 0.000 2774.175 3376.755 2775.015 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 0.000 2771.795 3588.000 2774.175 ;
        RECT 0.000 2770.955 3376.755 2771.795 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 0.000 2768.575 3588.000 2770.955 ;
        RECT 0.000 2767.735 3376.755 2768.575 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 0.000 2765.815 3588.000 2767.735 ;
        RECT 0.000 2764.975 3376.755 2765.815 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 0.000 2762.595 3588.000 2764.975 ;
        RECT 0.000 2761.755 3376.755 2762.595 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 0.000 2756.615 3588.000 2761.755 ;
        RECT 0.000 2755.775 3376.755 2756.615 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 0.000 2753.395 3588.000 2755.775 ;
        RECT 0.000 2752.555 3376.755 2753.395 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
        RECT 0.000 2750.175 3588.000 2752.555 ;
        RECT 0.000 2749.335 3376.755 2750.175 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 0.000 2744.195 3588.000 2749.335 ;
        RECT 0.000 2743.355 3376.755 2744.195 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
        RECT 0.000 2701.645 3588.000 2743.355 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 211.245 2700.805 3588.000 2701.645 ;
        RECT 0.000 2695.665 3588.000 2700.805 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
        RECT 211.245 2694.825 3588.000 2695.665 ;
        RECT 0.000 2692.445 3588.000 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 211.245 2691.605 3588.000 2692.445 ;
        RECT 0.000 2689.225 3588.000 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 211.245 2688.385 3588.000 2689.225 ;
        RECT 0.000 2683.245 3588.000 2688.385 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 211.245 2682.405 3588.000 2683.245 ;
        RECT 0.000 2680.025 3588.000 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
        RECT 211.245 2679.185 3588.000 2680.025 ;
        RECT 0.000 2677.265 3588.000 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 211.245 2676.425 3588.000 2677.265 ;
        RECT 0.000 2674.045 3588.000 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 211.245 2673.205 3588.000 2674.045 ;
        RECT 0.000 2670.825 3588.000 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 211.245 2669.985 3588.000 2670.825 ;
        RECT 0.000 2668.065 3588.000 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
        RECT 211.245 2667.225 3588.000 2668.065 ;
        RECT 0.000 2655.645 3588.000 2667.225 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 211.245 2654.805 3588.000 2655.645 ;
        RECT 0.000 2652.425 3588.000 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 211.245 2651.585 3588.000 2652.425 ;
        RECT 0.000 2649.205 3588.000 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 211.245 2648.365 3588.000 2649.205 ;
        RECT 0.000 2646.445 3588.000 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 211.245 2645.605 3588.000 2646.445 ;
        RECT 0.000 2637.245 3588.000 2645.605 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 211.245 2636.405 3588.000 2637.245 ;
        RECT 0.000 2634.025 3588.000 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 211.245 2633.185 3588.000 2634.025 ;
        RECT 0.000 2630.805 3588.000 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 211.245 2629.965 3588.000 2630.805 ;
        RECT 0.000 2628.045 3588.000 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
        RECT 211.245 2627.205 3588.000 2628.045 ;
        RECT 0.000 2063.645 3588.000 2627.205 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 211.245 2062.805 3588.000 2063.645 ;
        RECT 0.000 2057.665 3588.000 2062.805 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
        RECT 211.245 2056.825 3588.000 2057.665 ;
        RECT 0.000 2054.445 3588.000 2056.825 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 211.245 2053.605 3588.000 2054.445 ;
        RECT 0.000 2051.225 3588.000 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 211.245 2050.385 3588.000 2051.225 ;
        RECT 0.000 2045.245 3588.000 2050.385 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 211.245 2044.405 3588.000 2045.245 ;
        RECT 0.000 2042.025 3588.000 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
        RECT 211.245 2041.185 3588.000 2042.025 ;
        RECT 0.000 2039.265 3588.000 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 211.245 2038.425 3588.000 2039.265 ;
        RECT 0.000 2036.045 3588.000 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 211.245 2035.205 3588.000 2036.045 ;
        RECT 0.000 2032.825 3588.000 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 211.245 2031.985 3588.000 2032.825 ;
        RECT 0.000 2030.065 3588.000 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 211.245 2029.225 3588.000 2030.065 ;
        RECT 0.000 2017.645 3588.000 2029.225 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 211.245 2016.805 3588.000 2017.645 ;
        RECT 0.000 2014.425 3588.000 2016.805 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 211.245 2013.585 3588.000 2014.425 ;
        RECT 0.000 2011.205 3588.000 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 211.245 2010.365 3588.000 2011.205 ;
        RECT 0.000 2008.445 3588.000 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 211.245 2007.605 3588.000 2008.445 ;
        RECT 0.000 1999.245 3588.000 2007.605 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 211.245 1998.405 3588.000 1999.245 ;
        RECT 0.000 1996.025 3588.000 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 211.245 1995.185 3588.000 1996.025 ;
        RECT 0.000 1992.805 3588.000 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 211.245 1991.965 3588.000 1992.805 ;
        RECT 0.000 1990.045 3588.000 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
        RECT 211.245 1989.205 3588.000 1990.045 ;
        RECT 0.000 1931.795 3588.000 1989.205 ;
        RECT 0.000 1930.955 3376.755 1931.795 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 0.000 1929.035 3588.000 1930.955 ;
        RECT 0.000 1928.195 3376.755 1929.035 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 0.000 1925.815 3588.000 1928.195 ;
        RECT 0.000 1924.975 3376.755 1925.815 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 0.000 1922.595 3588.000 1924.975 ;
        RECT 0.000 1921.755 3376.755 1922.595 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 0.000 1913.395 3588.000 1921.755 ;
        RECT 0.000 1912.555 3376.755 1913.395 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 0.000 1910.635 3588.000 1912.555 ;
        RECT 0.000 1909.795 3376.755 1910.635 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 0.000 1907.415 3588.000 1909.795 ;
        RECT 0.000 1906.575 3376.755 1907.415 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 0.000 1904.195 3588.000 1906.575 ;
        RECT 0.000 1903.355 3376.755 1904.195 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 0.000 1891.775 3588.000 1903.355 ;
        RECT 0.000 1890.935 3376.755 1891.775 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 0.000 1889.015 3588.000 1890.935 ;
        RECT 0.000 1888.175 3376.755 1889.015 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 0.000 1885.795 3588.000 1888.175 ;
        RECT 0.000 1884.955 3376.755 1885.795 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 0.000 1882.575 3588.000 1884.955 ;
        RECT 0.000 1881.735 3376.755 1882.575 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 0.000 1876.595 3588.000 1881.735 ;
        RECT 0.000 1875.755 3376.755 1876.595 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 0.000 1867.395 3588.000 1875.755 ;
        RECT 0.000 1866.555 3376.755 1867.395 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 0.000 1864.175 3588.000 1866.555 ;
        RECT 0.000 1863.335 3376.755 1864.175 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
        RECT 0.000 1858.195 3588.000 1863.335 ;
        RECT 0.000 1857.355 3376.755 1858.195 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
        RECT 0.000 1847.645 3588.000 1857.355 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
        RECT 211.245 1846.805 3588.000 1847.645 ;
        RECT 0.000 1841.665 3588.000 1846.805 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
        RECT 211.245 1840.825 3588.000 1841.665 ;
        RECT 0.000 1838.445 3588.000 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 211.245 1837.605 3588.000 1838.445 ;
        RECT 0.000 1835.225 3588.000 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 211.245 1834.385 3588.000 1835.225 ;
        RECT 0.000 1829.245 3588.000 1834.385 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 211.245 1828.405 3588.000 1829.245 ;
        RECT 0.000 1826.025 3588.000 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
        RECT 211.245 1825.185 3588.000 1826.025 ;
        RECT 0.000 1823.265 3588.000 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 211.245 1822.425 3588.000 1823.265 ;
        RECT 0.000 1820.045 3588.000 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 211.245 1819.205 3588.000 1820.045 ;
        RECT 0.000 1816.825 3588.000 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 211.245 1815.985 3588.000 1816.825 ;
        RECT 0.000 1814.065 3588.000 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 211.245 1813.225 3588.000 1814.065 ;
        RECT 0.000 1801.645 3588.000 1813.225 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 211.245 1800.805 3588.000 1801.645 ;
        RECT 0.000 1798.425 3588.000 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 211.245 1797.585 3588.000 1798.425 ;
        RECT 0.000 1795.205 3588.000 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 211.245 1794.365 3588.000 1795.205 ;
        RECT 0.000 1792.445 3588.000 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 211.245 1791.605 3588.000 1792.445 ;
        RECT 0.000 1783.245 3588.000 1791.605 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 211.245 1782.405 3588.000 1783.245 ;
        RECT 0.000 1780.025 3588.000 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 211.245 1779.185 3588.000 1780.025 ;
        RECT 0.000 1776.805 3588.000 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 211.245 1775.965 3588.000 1776.805 ;
        RECT 0.000 1774.045 3588.000 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
        RECT 211.245 1773.205 3588.000 1774.045 ;
        RECT 0.000 1705.795 3588.000 1773.205 ;
        RECT 0.000 1704.955 3376.755 1705.795 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 0.000 1703.035 3588.000 1704.955 ;
        RECT 0.000 1702.195 3376.755 1703.035 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 0.000 1699.815 3588.000 1702.195 ;
        RECT 0.000 1698.975 3376.755 1699.815 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 0.000 1696.595 3588.000 1698.975 ;
        RECT 0.000 1695.755 3376.755 1696.595 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 0.000 1687.395 3588.000 1695.755 ;
        RECT 0.000 1686.555 3376.755 1687.395 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 0.000 1684.635 3588.000 1686.555 ;
        RECT 0.000 1683.795 3376.755 1684.635 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 0.000 1681.415 3588.000 1683.795 ;
        RECT 0.000 1680.575 3376.755 1681.415 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
        RECT 0.000 1678.195 3588.000 1680.575 ;
        RECT 0.000 1677.355 3376.755 1678.195 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
        RECT 0.000 1665.775 3588.000 1677.355 ;
        RECT 0.000 1664.935 3376.755 1665.775 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 0.000 1663.015 3588.000 1664.935 ;
        RECT 0.000 1662.175 3376.755 1663.015 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 0.000 1659.795 3588.000 1662.175 ;
        RECT 0.000 1658.955 3376.755 1659.795 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 0.000 1656.575 3588.000 1658.955 ;
        RECT 0.000 1655.735 3376.755 1656.575 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 0.000 1650.595 3588.000 1655.735 ;
        RECT 0.000 1649.755 3376.755 1650.595 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 0.000 1641.395 3588.000 1649.755 ;
        RECT 0.000 1640.555 3376.755 1641.395 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
        RECT 0.000 1638.175 3588.000 1640.555 ;
        RECT 0.000 1637.335 3376.755 1638.175 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 0.000 1632.195 3588.000 1637.335 ;
        RECT 0.000 1631.645 3376.755 1632.195 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 211.245 1631.355 3376.755 1631.645 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 211.245 1630.805 3588.000 1631.355 ;
        RECT 0.000 1625.665 3588.000 1630.805 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
        RECT 211.245 1624.825 3588.000 1625.665 ;
        RECT 0.000 1622.445 3588.000 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 211.245 1621.605 3588.000 1622.445 ;
        RECT 0.000 1619.225 3588.000 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 211.245 1618.385 3588.000 1619.225 ;
        RECT 0.000 1613.245 3588.000 1618.385 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 211.245 1612.405 3588.000 1613.245 ;
        RECT 0.000 1610.025 3588.000 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
        RECT 211.245 1609.185 3588.000 1610.025 ;
        RECT 0.000 1607.265 3588.000 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 211.245 1606.425 3588.000 1607.265 ;
        RECT 0.000 1604.045 3588.000 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 211.245 1603.205 3588.000 1604.045 ;
        RECT 0.000 1600.825 3588.000 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 211.245 1599.985 3588.000 1600.825 ;
        RECT 0.000 1598.065 3588.000 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
        RECT 211.245 1597.225 3588.000 1598.065 ;
        RECT 0.000 1585.645 3588.000 1597.225 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 211.245 1584.805 3588.000 1585.645 ;
        RECT 0.000 1582.425 3588.000 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 211.245 1581.585 3588.000 1582.425 ;
        RECT 0.000 1579.205 3588.000 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 211.245 1578.365 3588.000 1579.205 ;
        RECT 0.000 1576.445 3588.000 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 211.245 1575.605 3588.000 1576.445 ;
        RECT 0.000 1567.245 3588.000 1575.605 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 211.245 1566.405 3588.000 1567.245 ;
        RECT 0.000 1564.025 3588.000 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 211.245 1563.185 3588.000 1564.025 ;
        RECT 0.000 1560.805 3588.000 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 211.245 1559.965 3588.000 1560.805 ;
        RECT 0.000 1558.045 3588.000 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
        RECT 211.245 1557.205 3588.000 1558.045 ;
        RECT 0.000 1480.795 3588.000 1557.205 ;
        RECT 0.000 1479.955 3376.755 1480.795 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 0.000 1478.035 3588.000 1479.955 ;
        RECT 0.000 1477.195 3376.755 1478.035 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 0.000 1474.815 3588.000 1477.195 ;
        RECT 0.000 1473.975 3376.755 1474.815 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 0.000 1471.595 3588.000 1473.975 ;
        RECT 0.000 1470.755 3376.755 1471.595 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
        RECT 0.000 1462.395 3588.000 1470.755 ;
        RECT 0.000 1461.555 3376.755 1462.395 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 0.000 1459.635 3588.000 1461.555 ;
        RECT 0.000 1458.795 3376.755 1459.635 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 0.000 1456.415 3588.000 1458.795 ;
        RECT 0.000 1455.575 3376.755 1456.415 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 0.000 1453.195 3588.000 1455.575 ;
        RECT 0.000 1452.355 3376.755 1453.195 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 0.000 1440.775 3588.000 1452.355 ;
        RECT 0.000 1439.935 3376.755 1440.775 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 0.000 1438.015 3588.000 1439.935 ;
        RECT 0.000 1437.175 3376.755 1438.015 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 0.000 1434.795 3588.000 1437.175 ;
        RECT 0.000 1433.955 3376.755 1434.795 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 0.000 1431.575 3588.000 1433.955 ;
        RECT 0.000 1430.735 3376.755 1431.575 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 0.000 1425.595 3588.000 1430.735 ;
        RECT 0.000 1424.755 3376.755 1425.595 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 0.000 1416.395 3588.000 1424.755 ;
        RECT 0.000 1415.645 3376.755 1416.395 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 211.245 1415.555 3376.755 1415.645 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
        RECT 211.245 1414.805 3588.000 1415.555 ;
        RECT 0.000 1413.175 3588.000 1414.805 ;
        RECT 0.000 1412.335 3376.755 1413.175 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
        RECT 0.000 1409.665 3588.000 1412.335 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
        RECT 211.245 1408.825 3588.000 1409.665 ;
        RECT 0.000 1407.195 3588.000 1408.825 ;
        RECT 0.000 1406.445 3376.755 1407.195 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 211.245 1406.355 3376.755 1406.445 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
        RECT 211.245 1405.605 3588.000 1406.355 ;
        RECT 0.000 1403.225 3588.000 1405.605 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 211.245 1402.385 3588.000 1403.225 ;
        RECT 0.000 1397.245 3588.000 1402.385 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 211.245 1396.405 3588.000 1397.245 ;
        RECT 0.000 1394.025 3588.000 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
        RECT 211.245 1393.185 3588.000 1394.025 ;
        RECT 0.000 1391.265 3588.000 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 211.245 1390.425 3588.000 1391.265 ;
        RECT 0.000 1388.045 3588.000 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 211.245 1387.205 3588.000 1388.045 ;
        RECT 0.000 1384.825 3588.000 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 211.245 1383.985 3588.000 1384.825 ;
        RECT 0.000 1382.065 3588.000 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 211.245 1381.225 3588.000 1382.065 ;
        RECT 0.000 1369.645 3588.000 1381.225 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
        RECT 211.245 1368.805 3588.000 1369.645 ;
        RECT 0.000 1366.425 3588.000 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 211.245 1365.585 3588.000 1366.425 ;
        RECT 0.000 1363.205 3588.000 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 211.245 1362.365 3588.000 1363.205 ;
        RECT 0.000 1360.445 3588.000 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 211.245 1359.605 3588.000 1360.445 ;
        RECT 0.000 1351.245 3588.000 1359.605 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 211.245 1350.405 3588.000 1351.245 ;
        RECT 0.000 1348.025 3588.000 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 211.245 1347.185 3588.000 1348.025 ;
        RECT 0.000 1344.805 3588.000 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 211.245 1343.965 3588.000 1344.805 ;
        RECT 0.000 1342.045 3588.000 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
        RECT 211.245 1341.205 3588.000 1342.045 ;
        RECT 0.000 1255.795 3588.000 1341.205 ;
        RECT 0.000 1254.955 3376.755 1255.795 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 0.000 1253.035 3588.000 1254.955 ;
        RECT 0.000 1252.195 3376.755 1253.035 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 0.000 1249.815 3588.000 1252.195 ;
        RECT 0.000 1248.975 3376.755 1249.815 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 0.000 1246.595 3588.000 1248.975 ;
        RECT 0.000 1245.755 3376.755 1246.595 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 0.000 1237.395 3588.000 1245.755 ;
        RECT 0.000 1236.555 3376.755 1237.395 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 0.000 1234.635 3588.000 1236.555 ;
        RECT 0.000 1233.795 3376.755 1234.635 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 0.000 1231.415 3588.000 1233.795 ;
        RECT 0.000 1230.575 3376.755 1231.415 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 0.000 1228.195 3588.000 1230.575 ;
        RECT 0.000 1227.355 3376.755 1228.195 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 0.000 1215.775 3588.000 1227.355 ;
        RECT 0.000 1214.935 3376.755 1215.775 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 0.000 1213.015 3588.000 1214.935 ;
        RECT 0.000 1212.175 3376.755 1213.015 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 0.000 1209.795 3588.000 1212.175 ;
        RECT 0.000 1208.955 3376.755 1209.795 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 0.000 1206.575 3588.000 1208.955 ;
        RECT 0.000 1205.735 3376.755 1206.575 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 0.000 1200.595 3588.000 1205.735 ;
        RECT 0.000 1199.755 3376.755 1200.595 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 0.000 1199.645 3588.000 1199.755 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
        RECT 211.245 1198.805 3588.000 1199.645 ;
        RECT 0.000 1193.665 3588.000 1198.805 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
        RECT 211.245 1192.825 3588.000 1193.665 ;
        RECT 0.000 1191.395 3588.000 1192.825 ;
        RECT 0.000 1190.555 3376.755 1191.395 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
        RECT 0.000 1190.445 3588.000 1190.555 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
        RECT 211.245 1189.605 3588.000 1190.445 ;
        RECT 0.000 1188.175 3588.000 1189.605 ;
        RECT 0.000 1187.335 3376.755 1188.175 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
        RECT 0.000 1182.195 3588.000 1187.335 ;
        RECT 0.000 1181.355 3376.755 1182.195 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
        RECT 0.000 1181.245 3588.000 1181.355 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 211.245 1180.405 3588.000 1181.245 ;
        RECT 0.000 1175.265 3588.000 1180.405 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 211.245 1174.425 3588.000 1175.265 ;
        RECT 0.000 1172.045 3588.000 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 211.245 1171.205 3588.000 1172.045 ;
        RECT 0.000 1168.825 3588.000 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 211.245 1167.985 3588.000 1168.825 ;
        RECT 0.000 1166.065 3588.000 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 211.245 1165.225 3588.000 1166.065 ;
        RECT 0.000 1153.645 3588.000 1165.225 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 211.245 1152.805 3588.000 1153.645 ;
        RECT 0.000 1150.425 3588.000 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 211.245 1149.585 3588.000 1150.425 ;
        RECT 0.000 1147.205 3588.000 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 211.245 1146.365 3588.000 1147.205 ;
        RECT 0.000 1144.445 3588.000 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 211.245 1143.605 3588.000 1144.445 ;
        RECT 0.000 1135.245 3588.000 1143.605 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 211.245 1134.405 3588.000 1135.245 ;
        RECT 0.000 1132.025 3588.000 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 211.245 1131.185 3588.000 1132.025 ;
        RECT 0.000 1128.805 3588.000 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 211.245 1127.965 3588.000 1128.805 ;
        RECT 0.000 1126.045 3588.000 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
        RECT 211.245 1125.205 3588.000 1126.045 ;
        RECT 0.000 1029.795 3588.000 1125.205 ;
        RECT 0.000 1028.955 3376.755 1029.795 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
        RECT 0.000 1027.035 3588.000 1028.955 ;
        RECT 0.000 1026.195 3376.755 1027.035 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 0.000 1023.815 3588.000 1026.195 ;
        RECT 0.000 1022.975 3376.755 1023.815 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 0.000 1020.595 3588.000 1022.975 ;
        RECT 0.000 1019.755 3376.755 1020.595 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 0.000 1011.395 3588.000 1019.755 ;
        RECT 0.000 1010.555 3376.755 1011.395 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 0.000 1008.635 3588.000 1010.555 ;
        RECT 0.000 1007.795 3376.755 1008.635 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 0.000 1005.415 3588.000 1007.795 ;
        RECT 0.000 1004.575 3376.755 1005.415 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 0.000 1002.195 3588.000 1004.575 ;
        RECT 0.000 1001.355 3376.755 1002.195 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
        RECT 0.000 989.775 3588.000 1001.355 ;
        RECT 0.000 988.935 3376.755 989.775 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 0.000 987.015 3588.000 988.935 ;
        RECT 0.000 986.175 3376.755 987.015 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 0.000 983.795 3588.000 986.175 ;
        RECT 0.000 983.645 3376.755 983.795 ;
        RECT 0.000 982.805 208.285 983.645 ;
        RECT 211.245 982.955 3376.755 983.645 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 211.245 982.805 3588.000 982.955 ;
        RECT 0.000 980.575 3588.000 982.805 ;
        RECT 0.000 979.735 3376.755 980.575 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 0.000 977.665 3588.000 979.735 ;
        RECT 0.000 976.825 208.285 977.665 ;
        RECT 211.245 976.825 3588.000 977.665 ;
        RECT 0.000 974.595 3588.000 976.825 ;
        RECT 0.000 974.445 3376.755 974.595 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 211.245 973.755 3376.755 974.445 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 211.245 973.605 3588.000 973.755 ;
        RECT 0.000 965.395 3588.000 973.605 ;
        RECT 0.000 965.245 3376.755 965.395 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 211.245 964.555 3376.755 965.245 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 211.245 964.405 3588.000 964.555 ;
        RECT 0.000 962.175 3588.000 964.405 ;
        RECT 0.000 961.335 3376.755 962.175 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
        RECT 0.000 959.265 3588.000 961.335 ;
        RECT 0.000 958.425 208.285 959.265 ;
        RECT 211.245 958.425 3588.000 959.265 ;
        RECT 0.000 956.195 3588.000 958.425 ;
        RECT 0.000 956.045 3376.755 956.195 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 211.245 955.355 3376.755 956.045 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 211.245 955.205 3588.000 955.355 ;
        RECT 0.000 952.825 3588.000 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
        RECT 211.245 951.985 3588.000 952.825 ;
        RECT 0.000 950.065 3588.000 951.985 ;
        RECT 0.000 949.225 208.285 950.065 ;
        RECT 211.245 949.225 3588.000 950.065 ;
        RECT 0.000 937.645 3588.000 949.225 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 211.245 936.805 3588.000 937.645 ;
        RECT 0.000 934.425 3588.000 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 211.245 933.585 3588.000 934.425 ;
        RECT 0.000 931.205 3588.000 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 211.245 930.365 3588.000 931.205 ;
        RECT 0.000 928.445 3588.000 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 211.245 927.605 3588.000 928.445 ;
        RECT 0.000 919.245 3588.000 927.605 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 211.245 918.405 3588.000 919.245 ;
        RECT 0.000 916.025 3588.000 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 211.245 915.185 3588.000 916.025 ;
        RECT 0.000 912.805 3588.000 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 211.245 911.965 3588.000 912.805 ;
        RECT 0.000 910.045 3588.000 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
        RECT 211.245 909.205 3588.000 910.045 ;
        RECT 0.000 804.795 3588.000 909.205 ;
        RECT 0.000 803.955 3376.755 804.795 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 0.000 802.035 3588.000 803.955 ;
        RECT 0.000 801.195 3376.755 802.035 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 0.000 798.815 3588.000 801.195 ;
        RECT 0.000 797.975 3376.755 798.815 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 0.000 795.595 3588.000 797.975 ;
        RECT 0.000 794.755 3376.755 795.595 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
        RECT 0.000 786.395 3588.000 794.755 ;
        RECT 0.000 785.555 3376.755 786.395 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 0.000 783.635 3588.000 785.555 ;
        RECT 0.000 782.795 3376.755 783.635 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 0.000 780.415 3588.000 782.795 ;
        RECT 0.000 779.575 3376.755 780.415 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 0.000 777.195 3588.000 779.575 ;
        RECT 0.000 776.355 3376.755 777.195 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
        RECT 0.000 764.775 3588.000 776.355 ;
        RECT 0.000 763.935 3376.755 764.775 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 0.000 762.015 3588.000 763.935 ;
        RECT 0.000 761.175 3376.755 762.015 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 0.000 758.795 3588.000 761.175 ;
        RECT 0.000 757.955 3376.755 758.795 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 0.000 755.575 3588.000 757.955 ;
        RECT 0.000 754.735 3376.755 755.575 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 0.000 749.595 3588.000 754.735 ;
        RECT 0.000 748.755 3376.755 749.595 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 0.000 740.395 3588.000 748.755 ;
        RECT 0.000 739.555 3376.755 740.395 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 0.000 737.175 3588.000 739.555 ;
        RECT 0.000 736.335 3376.755 737.175 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
        RECT 0.000 731.195 3588.000 736.335 ;
        RECT 0.000 730.355 3376.755 731.195 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
        RECT 0.000 578.795 3588.000 730.355 ;
        RECT 0.000 577.955 3376.755 578.795 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 0.000 576.035 3588.000 577.955 ;
        RECT 0.000 575.195 3376.755 576.035 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 0.000 572.815 3588.000 575.195 ;
        RECT 0.000 571.975 3376.755 572.815 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 0.000 569.595 3588.000 571.975 ;
        RECT 0.000 568.755 3376.755 569.595 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 0.000 560.395 3588.000 568.755 ;
        RECT 0.000 559.555 3376.755 560.395 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 0.000 557.635 3588.000 559.555 ;
        RECT 0.000 556.795 3376.755 557.635 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 0.000 554.415 3588.000 556.795 ;
        RECT 0.000 553.575 3376.755 554.415 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 0.000 551.195 3588.000 553.575 ;
        RECT 0.000 550.355 3376.755 551.195 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 0.000 538.775 3588.000 550.355 ;
        RECT 0.000 537.935 3376.755 538.775 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 0.000 536.015 3588.000 537.935 ;
        RECT 0.000 535.175 3376.755 536.015 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 0.000 532.795 3588.000 535.175 ;
        RECT 0.000 531.955 3376.755 532.795 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 0.000 529.575 3588.000 531.955 ;
        RECT 0.000 528.735 3376.755 529.575 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 0.000 523.595 3588.000 528.735 ;
        RECT 0.000 522.755 3376.755 523.595 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 0.000 514.395 3588.000 522.755 ;
        RECT 0.000 513.555 3376.755 514.395 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 0.000 511.175 3588.000 513.555 ;
        RECT 0.000 510.335 3376.755 511.175 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
        RECT 0.000 505.195 3588.000 510.335 ;
        RECT 0.000 504.355 3376.755 505.195 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
        RECT 0.000 211.410 3588.000 504.355 ;
        RECT 0.000 211.245 1540.995 211.410 ;
        RECT 0.000 208.285 936.355 211.245 ;
        RECT 937.195 208.285 969.935 211.245 ;
        RECT 970.775 208.285 1534.555 211.245 ;
        RECT 1535.395 208.450 1540.995 211.245 ;
        RECT 1541.835 211.245 2624.575 211.410 ;
        RECT 1541.835 208.450 1808.555 211.245 ;
        RECT 1535.395 208.285 1808.555 208.450 ;
        RECT 1809.395 208.285 2027.355 211.245 ;
        RECT 2028.195 208.285 2060.935 211.245 ;
        RECT 2061.775 208.285 2082.555 211.245 ;
        RECT 2083.395 208.285 2098.195 211.245 ;
        RECT 2099.035 208.285 2301.355 211.245 ;
        RECT 2302.195 208.285 2334.935 211.245 ;
        RECT 2335.775 208.285 2356.555 211.245 ;
        RECT 2357.395 208.285 2372.195 211.245 ;
        RECT 2373.035 208.285 2575.355 211.245 ;
        RECT 2576.195 208.285 2602.955 211.245 ;
        RECT 2603.795 208.285 2608.935 211.245 ;
        RECT 2609.775 208.450 2624.575 211.245 ;
        RECT 2625.415 211.245 3588.000 211.410 ;
        RECT 2625.415 208.450 2630.555 211.245 ;
        RECT 2609.775 208.285 2630.555 208.450 ;
        RECT 2631.395 208.285 3588.000 211.245 ;
        RECT 0.000 200.280 3588.000 208.285 ;
        RECT 0.000 199.390 708.055 200.280 ;
        RECT 709.345 199.390 3588.000 200.280 ;
        RECT 0.000 195.905 3588.000 199.390 ;
        RECT 0.000 195.245 1551.015 195.905 ;
        RECT 1551.675 195.245 1825.015 195.905 ;
        RECT 1825.675 195.245 2647.015 195.905 ;
        RECT 2647.675 195.245 3588.000 195.905 ;
        RECT 0.000 0.000 3588.000 195.245 ;
      LAYER met3 ;
        RECT 0.000 5073.175 3588.000 5188.000 ;
        RECT 0.000 5071.375 1225.890 5073.175 ;
        RECT 1227.690 5071.375 1488.890 5073.175 ;
        RECT 1490.690 5071.375 1997.890 5073.175 ;
        RECT 1999.690 5071.375 3588.000 5073.175 ;
        RECT 0.000 5071.270 3588.000 5071.375 ;
        RECT 0.000 5061.205 386.055 5071.270 ;
        RECT 396.120 5061.205 643.055 5071.270 ;
        RECT 653.120 5061.205 900.055 5071.270 ;
        RECT 910.120 5061.205 2369.055 5071.270 ;
        RECT 2379.120 5061.205 2626.055 5071.270 ;
        RECT 2636.120 5061.205 3135.055 5071.270 ;
        RECT 3145.120 5061.205 3588.000 5071.270 ;
        RECT 0.000 4832.715 3588.000 5061.205 ;
        RECT 0.000 4818.120 103.455 4832.715 ;
        RECT 118.050 4823.680 3588.000 4832.715 ;
        RECT 118.050 4818.120 3446.205 4823.680 ;
        RECT 0.000 4807.880 3446.205 4818.120 ;
        RECT 3462.005 4807.880 3588.000 4823.680 ;
        RECT 0.000 0.000 3588.000 4807.880 ;
      LAYER met4 ;
        RECT 0.000 2374.400 3588.000 5188.000 ;
        RECT 0.000 2300.360 3444.005 2374.400 ;
        RECT 0.000 2298.600 3402.535 2300.360 ;
        RECT 3406.785 2298.600 3444.005 2300.360 ;
        RECT 3445.135 2298.600 3588.000 2374.400 ;
        RECT 0.000 2280.870 3588.000 2298.600 ;
        RECT 0.000 2280.515 0.335 2280.870 ;
        RECT 0.000 2280.470 24.215 2280.515 ;
        RECT 24.615 2279.400 3588.000 2280.870 ;
        RECT 0.000 2277.825 0.175 2278.225 ;
        RECT 24.615 2277.825 142.865 2279.400 ;
        RECT 0.000 2203.600 142.865 2277.825 ;
        RECT 143.995 2277.330 164.265 2279.400 ;
        RECT 168.515 2279.395 192.115 2279.400 ;
        RECT 168.515 2277.635 181.215 2279.395 ;
        RECT 185.465 2277.635 192.115 2279.395 ;
        RECT 168.515 2277.330 192.115 2277.635 ;
        RECT 198.365 2277.330 3588.000 2279.400 ;
        RECT 143.995 2203.600 3588.000 2277.330 ;
        RECT 0.000 187.460 3588.000 2203.600 ;
        RECT 0.000 184.665 191.760 187.460 ;
        RECT 194.555 184.665 3588.000 187.460 ;
        RECT 0.000 158.815 3588.000 184.665 ;
        RECT 0.000 153.365 662.600 158.815 ;
        RECT 664.670 153.365 3588.000 158.815 ;
        RECT 0.000 144.295 3588.000 153.365 ;
        RECT 0.000 143.195 176.265 144.295 ;
        RECT 177.365 143.195 3588.000 144.295 ;
        RECT 0.000 0.000 3588.000 143.195 ;
      LAYER met5 ;
        RECT 0.000 5155.540 3588.000 5188.000 ;
        RECT 0.000 5091.520 391.450 5155.540 ;
        RECT 455.490 5091.520 648.450 5155.540 ;
        RECT 712.490 5091.520 905.450 5155.540 ;
        RECT 969.490 5091.520 1157.450 5155.540 ;
        RECT 1221.490 5091.520 1420.450 5155.540 ;
        RECT 1484.490 5091.520 1672.450 5155.540 ;
        RECT 1736.490 5091.520 1929.450 5155.540 ;
        RECT 1993.490 5091.520 2374.450 5155.540 ;
        RECT 2438.490 5091.520 2631.450 5155.540 ;
        RECT 2695.490 5091.520 2883.450 5155.540 ;
        RECT 2947.490 5091.520 3140.450 5155.540 ;
        RECT 3204.490 5091.520 3588.000 5155.540 ;
        RECT 0.000 4847.680 3588.000 5091.520 ;
        RECT 0.000 4842.865 94.290 4847.680 ;
        RECT 99.105 4842.865 3588.000 4847.680 ;
        RECT 0.000 4829.680 3588.000 4842.865 ;
        RECT 0.000 4824.865 3553.090 4829.680 ;
        RECT 3557.905 4824.865 3588.000 4829.680 ;
        RECT 0.000 4628.465 3588.000 4824.865 ;
        RECT 0.000 4623.665 97.505 4628.465 ;
        RECT 102.305 4623.665 3588.000 4628.465 ;
        RECT 0.000 4606.465 3588.000 4623.665 ;
        RECT 0.000 4601.665 3556.305 4606.465 ;
        RECT 3561.105 4601.665 3588.000 4606.465 ;
        RECT 0.000 4420.680 3588.000 4601.665 ;
        RECT 0.000 4415.865 94.290 4420.680 ;
        RECT 99.105 4415.865 3588.000 4420.680 ;
        RECT 0.000 4383.800 3588.000 4415.865 ;
        RECT 0.000 4379.135 3489.550 4383.800 ;
        RECT 3494.215 4379.135 3588.000 4383.800 ;
        RECT 0.000 4209.680 3588.000 4379.135 ;
        RECT 0.000 4204.865 94.290 4209.680 ;
        RECT 99.105 4204.865 3588.000 4209.680 ;
        RECT 0.000 4163.680 3588.000 4204.865 ;
        RECT 0.000 4158.865 3553.090 4163.680 ;
        RECT 3557.905 4158.865 3588.000 4163.680 ;
        RECT 0.000 3998.800 3588.000 4158.865 ;
        RECT 0.000 3994.135 29.980 3998.800 ;
        RECT 34.645 3994.135 3588.000 3998.800 ;
        RECT 0.000 3937.800 3588.000 3994.135 ;
        RECT 0.000 3933.135 3489.550 3937.800 ;
        RECT 3494.215 3933.135 3588.000 3937.800 ;
        RECT 0.000 3782.800 3588.000 3933.135 ;
        RECT 0.000 3778.135 29.980 3782.800 ;
        RECT 34.645 3778.135 3588.000 3782.800 ;
        RECT 0.000 3712.800 3588.000 3778.135 ;
        RECT 0.000 3708.135 3489.550 3712.800 ;
        RECT 3494.215 3708.135 3588.000 3712.800 ;
        RECT 0.000 3566.800 3588.000 3708.135 ;
        RECT 0.000 3562.135 29.980 3566.800 ;
        RECT 34.645 3562.135 3588.000 3566.800 ;
        RECT 0.000 3487.800 3588.000 3562.135 ;
        RECT 0.000 3483.135 3489.550 3487.800 ;
        RECT 3494.215 3483.135 3588.000 3487.800 ;
        RECT 0.000 3350.800 3588.000 3483.135 ;
        RECT 0.000 3346.135 29.980 3350.800 ;
        RECT 34.645 3346.135 3588.000 3350.800 ;
        RECT 0.000 3261.800 3588.000 3346.135 ;
        RECT 0.000 3257.135 3489.550 3261.800 ;
        RECT 3494.215 3257.135 3588.000 3261.800 ;
        RECT 0.000 3134.800 3588.000 3257.135 ;
        RECT 0.000 3130.135 29.980 3134.800 ;
        RECT 34.645 3130.135 3588.000 3134.800 ;
        RECT 0.000 3036.800 3588.000 3130.135 ;
        RECT 0.000 3032.135 3489.550 3036.800 ;
        RECT 3494.215 3032.135 3588.000 3036.800 ;
        RECT 0.000 2918.800 3588.000 3032.135 ;
        RECT 0.000 2914.135 29.980 2918.800 ;
        RECT 34.645 2914.135 3588.000 2918.800 ;
        RECT 0.000 2810.800 3588.000 2914.135 ;
        RECT 0.000 2806.135 3489.550 2810.800 ;
        RECT 3494.215 2806.135 3588.000 2810.800 ;
        RECT 0.000 2702.800 3588.000 2806.135 ;
        RECT 0.000 2698.135 29.980 2702.800 ;
        RECT 34.645 2698.135 3588.000 2702.800 ;
        RECT 0.000 2590.680 3588.000 2698.135 ;
        RECT 0.000 2585.865 3553.090 2590.680 ;
        RECT 3557.905 2585.865 3588.000 2590.680 ;
        RECT 0.000 2486.680 3588.000 2585.865 ;
        RECT 0.000 2481.865 94.290 2486.680 ;
        RECT 99.105 2481.865 3588.000 2486.680 ;
        RECT 0.000 2367.465 3588.000 2481.865 ;
        RECT 0.000 2362.665 3556.305 2367.465 ;
        RECT 3561.105 2362.665 3588.000 2367.465 ;
        RECT 0.000 2272.465 3588.000 2362.665 ;
        RECT 0.000 2267.665 97.505 2272.465 ;
        RECT 102.305 2267.665 3588.000 2272.465 ;
        RECT 0.000 2149.680 3588.000 2267.665 ;
        RECT 0.000 2144.865 3553.090 2149.680 ;
        RECT 3557.905 2144.865 3588.000 2149.680 ;
        RECT 0.000 2064.800 3588.000 2144.865 ;
        RECT 0.000 2060.135 29.980 2064.800 ;
        RECT 34.645 2060.135 3588.000 2064.800 ;
        RECT 0.000 1924.800 3588.000 2060.135 ;
        RECT 0.000 1920.135 3489.550 1924.800 ;
        RECT 3494.215 1920.135 3588.000 1924.800 ;
        RECT 0.000 1848.800 3588.000 1920.135 ;
        RECT 0.000 1844.135 29.980 1848.800 ;
        RECT 34.645 1844.135 3588.000 1848.800 ;
        RECT 0.000 1698.800 3588.000 1844.135 ;
        RECT 0.000 1694.135 3489.550 1698.800 ;
        RECT 3494.215 1694.135 3588.000 1698.800 ;
        RECT 0.000 1632.800 3588.000 1694.135 ;
        RECT 0.000 1628.135 29.980 1632.800 ;
        RECT 34.645 1628.135 3588.000 1632.800 ;
        RECT 0.000 1473.800 3588.000 1628.135 ;
        RECT 0.000 1469.135 3489.550 1473.800 ;
        RECT 3494.215 1469.135 3588.000 1473.800 ;
        RECT 0.000 1416.800 3588.000 1469.135 ;
        RECT 0.000 1412.135 29.980 1416.800 ;
        RECT 34.645 1412.135 3588.000 1416.800 ;
        RECT 0.000 1248.800 3588.000 1412.135 ;
        RECT 0.000 1244.135 3489.550 1248.800 ;
        RECT 3494.215 1244.135 3588.000 1248.800 ;
        RECT 0.000 1200.800 3588.000 1244.135 ;
        RECT 0.000 1196.135 29.980 1200.800 ;
        RECT 34.645 1196.135 3588.000 1200.800 ;
        RECT 0.000 1022.800 3588.000 1196.135 ;
        RECT 0.000 1018.135 3489.550 1022.800 ;
        RECT 3494.215 1018.135 3588.000 1022.800 ;
        RECT 0.000 984.800 3588.000 1018.135 ;
        RECT 0.000 980.135 29.980 984.800 ;
        RECT 34.645 980.135 3588.000 984.800 ;
        RECT 0.000 797.800 3588.000 980.135 ;
        RECT 0.000 793.135 3489.550 797.800 ;
        RECT 3494.215 793.135 3588.000 797.800 ;
        RECT 0.000 622.680 3588.000 793.135 ;
        RECT 0.000 617.865 94.290 622.680 ;
        RECT 99.105 617.865 3588.000 622.680 ;
        RECT 0.000 571.800 3588.000 617.865 ;
        RECT 0.000 567.135 3489.550 571.800 ;
        RECT 3494.215 567.135 3588.000 571.800 ;
        RECT 0.000 408.465 3588.000 567.135 ;
        RECT 0.000 403.665 97.505 408.465 ;
        RECT 102.305 403.665 3588.000 408.465 ;
        RECT 0.000 101.970 3588.000 403.665 ;
        RECT 0.000 98.655 1270.000 101.970 ;
        RECT 0.000 96.475 935.255 98.655 ;
        RECT 0.000 32.455 399.510 96.475 ;
        RECT 463.550 93.840 935.255 96.475 ;
        RECT 940.070 97.170 1270.000 98.655 ;
        RECT 1274.800 98.655 3588.000 101.970 ;
        RECT 1274.800 97.170 1478.255 98.655 ;
        RECT 940.070 93.840 1478.255 97.170 ;
        RECT 1483.070 93.840 1752.255 98.655 ;
        RECT 1757.070 93.840 2026.255 98.655 ;
        RECT 2031.070 93.840 2300.255 98.655 ;
        RECT 2305.070 93.840 2574.255 98.655 ;
        RECT 2579.070 96.475 3588.000 98.655 ;
        RECT 2579.070 93.840 2850.510 96.475 ;
        RECT 463.550 93.145 2850.510 93.840 ;
        RECT 463.550 34.115 681.965 93.145 ;
        RECT 722.345 34.115 2850.510 93.145 ;
        RECT 463.550 32.455 2850.510 34.115 ;
        RECT 2914.550 32.455 3119.510 96.475 ;
        RECT 3183.550 32.455 3588.000 96.475 ;
        RECT 0.000 0.000 3588.000 32.455 ;
  END
END chip_io_alt
END LIBRARY

