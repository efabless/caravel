VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_power_routing
  CLASS BLOCK ;
  FOREIGN caravel_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  OBS
      LAYER met1 ;
        RECT 3240.520 232.950 3250.800 235.940 ;
      LAYER met2 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
      LAYER met3 ;
        RECT 30.110 169.500 3559.070 5158.480 ;
      LAYER met4 ;
        RECT 30.530 169.790 3558.650 5158.060 ;
      LAYER met5 ;
        RECT 30.170 213.940 3558.940 5158.390 ;
  END
END caravel_power_routing
END LIBRARY

