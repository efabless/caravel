magic
tech sky130A
magscale 1 2
timestamp 1665711229
<< locali >>
rect 416588 996667 416806 996673
rect 662589 996585 662807 996591
rect 663785 996585 664003 996591
rect 664981 996585 665199 996591
rect 666177 996585 666395 996591
rect 167978 996342 168196 996348
rect 169174 996342 169392 996348
rect 170370 996342 170588 996348
rect 40596 891200 40602 891418
rect 40596 890004 40602 890222
rect 40596 888808 40602 889026
rect 40596 887612 40602 887830
rect 40596 886416 40602 886634
rect 676932 714240 676938 714458
rect 676932 713044 676938 713262
rect 676932 711848 676938 712066
rect 676932 710652 676938 710870
rect 676932 709456 676938 709674
rect 676932 708260 676938 708478
rect 40621 610554 40627 610772
rect 40621 609358 40627 609576
rect 40621 608162 40627 608380
rect 40621 606966 40627 607184
rect 40621 605770 40627 605988
rect 40621 604574 40627 604792
rect 40621 603378 40627 603596
rect 40621 602182 40627 602400
rect 40621 600986 40627 601204
rect 40621 599790 40627 600008
rect 40621 598594 40627 598812
rect 676932 453416 676938 453634
rect 676932 452220 676938 452438
rect 676932 451024 676938 451242
rect 676932 449828 676938 450046
rect 676932 448632 676938 448850
rect 676932 447436 676938 447654
rect 676932 446240 676938 446458
rect 676932 445044 676938 445262
rect 676932 443848 676938 444066
rect 676932 442652 676938 442870
rect 676932 441456 676938 441674
rect 676932 440260 676938 440478
rect 40643 352373 40649 352591
rect 40643 351177 40649 351395
rect 40643 349981 40649 350199
rect 40643 348785 40649 349003
rect 40643 347589 40649 347807
rect 40643 346393 40649 346611
rect 40643 345197 40649 345415
rect 40643 344001 40649 344219
rect 40643 342805 40649 343023
rect 40643 341609 40649 341827
rect 40643 340413 40649 340631
rect 40643 339217 40649 339435
rect 40643 338021 40649 338239
rect 40643 336825 40649 337043
rect 40643 335629 40649 335847
rect 134848 223204 135066 223210
rect 136044 223204 136262 223210
rect 137240 223204 137458 223210
rect 138436 223204 138654 223210
rect 139632 223204 139850 223210
rect 140828 223204 141046 223210
rect 142024 223204 142242 223210
rect 143220 223204 143438 223210
rect 144416 223204 144634 223210
rect 145612 223204 145830 223210
rect 146808 223204 147026 223210
rect 148004 223204 148222 223210
rect 149200 223204 149418 223210
rect 150396 223204 150614 223210
rect 151592 223204 151810 223210
rect 152788 223204 153006 223210
rect 153984 223204 154202 223210
rect 155180 223204 155398 223210
rect 156376 223204 156594 223210
rect 157572 223204 157790 223210
rect 158768 223204 158986 223210
rect 394848 223204 395066 223210
rect 396044 223204 396262 223210
rect 397240 223204 397458 223210
rect 398436 223204 398654 223210
rect 399632 223204 399850 223210
rect 400828 223204 401046 223210
rect 402024 223204 402242 223210
rect 403220 223204 403438 223210
rect 404416 223204 404634 223210
rect 405612 223204 405830 223210
rect 406808 223204 407026 223210
rect 408004 223204 408222 223210
rect 409200 223204 409418 223210
rect 410396 223204 410614 223210
rect 411592 223204 411810 223210
rect 412788 223204 413006 223210
rect 413984 223204 414202 223210
rect 415180 223204 415398 223210
rect 416376 223204 416594 223210
rect 417572 223204 417790 223210
rect 418768 223204 418986 223210
<< viali >>
rect 416870 997217 416904 997387
rect 417514 997285 417732 997319
rect 662871 997135 662905 997305
rect 663515 997203 663733 997237
rect 664067 997135 664101 997305
rect 664711 997203 664929 997237
rect 665263 997135 665297 997305
rect 665907 997203 666125 997237
rect 666459 997135 666493 997305
rect 667103 997203 667321 997237
rect 167052 996960 167270 996994
rect 167880 996892 167914 997062
rect 168248 996960 168466 996994
rect 169076 996892 169110 997062
rect 169444 996960 169662 996994
rect 170272 996892 170306 997062
rect 416588 996673 416806 996707
rect 417516 996605 417550 996775
rect 662589 996591 662807 996625
rect 663517 996523 663551 996693
rect 663785 996591 664003 996625
rect 664713 996523 664747 996693
rect 664981 996591 665199 996625
rect 665909 996523 665943 996693
rect 666177 996591 666395 996625
rect 667105 996523 667139 996693
rect 167234 996280 167268 996450
rect 167978 996348 168196 996382
rect 168430 996280 168464 996450
rect 169174 996348 169392 996382
rect 169626 996280 169660 996450
rect 170370 996348 170588 996382
rect 40562 891200 40596 891418
rect 39882 891102 40052 891136
rect 39950 890274 39984 890492
rect 40494 890456 40664 890490
rect 40562 890004 40596 890222
rect 39882 889906 40052 889940
rect 39950 889078 39984 889296
rect 40494 889260 40664 889294
rect 40562 888808 40596 889026
rect 39882 888710 40052 888744
rect 39950 887882 39984 888100
rect 40494 888064 40664 888098
rect 40562 887612 40596 887830
rect 39882 887514 40052 887548
rect 39950 886686 39984 886904
rect 40494 886868 40664 886902
rect 40562 886416 40596 886634
rect 39882 886318 40052 886352
rect 39950 885490 39984 885708
rect 40494 885672 40664 885706
rect 676938 714240 676972 714458
rect 677482 714142 677652 714176
rect 676870 713496 677040 713530
rect 677550 713314 677584 713532
rect 676938 713044 676972 713262
rect 677482 712946 677652 712980
rect 676870 712300 677040 712334
rect 677550 712118 677584 712336
rect 676938 711848 676972 712066
rect 677482 711750 677652 711784
rect 676870 711104 677040 711138
rect 677550 710922 677584 711140
rect 676938 710652 676972 710870
rect 677482 710554 677652 710588
rect 676870 709908 677040 709942
rect 677550 709726 677584 709944
rect 676938 709456 676972 709674
rect 677482 709358 677652 709392
rect 676870 708712 677040 708746
rect 677550 708530 677584 708748
rect 676938 708260 676972 708478
rect 677482 708162 677652 708196
rect 676870 707516 677040 707550
rect 677550 707334 677584 707552
rect 40587 610554 40621 610772
rect 39907 610456 40077 610490
rect 39975 609628 40009 609846
rect 40519 609810 40689 609844
rect 40587 609358 40621 609576
rect 39907 609260 40077 609294
rect 39975 608432 40009 608650
rect 40519 608614 40689 608648
rect 40587 608162 40621 608380
rect 39907 608064 40077 608098
rect 39975 607236 40009 607454
rect 40519 607418 40689 607452
rect 40587 606966 40621 607184
rect 39907 606868 40077 606902
rect 39975 606040 40009 606258
rect 40519 606222 40689 606256
rect 40587 605770 40621 605988
rect 39907 605672 40077 605706
rect 39975 604844 40009 605062
rect 40519 605026 40689 605060
rect 40587 604574 40621 604792
rect 39907 604476 40077 604510
rect 39975 603648 40009 603866
rect 40519 603830 40689 603864
rect 40587 603378 40621 603596
rect 39907 603280 40077 603314
rect 39975 602452 40009 602670
rect 40519 602634 40689 602668
rect 40587 602182 40621 602400
rect 39907 602084 40077 602118
rect 39975 601256 40009 601474
rect 40519 601438 40689 601472
rect 40587 600986 40621 601204
rect 39907 600888 40077 600922
rect 39975 600060 40009 600278
rect 40519 600242 40689 600276
rect 40587 599790 40621 600008
rect 39907 599692 40077 599726
rect 39975 598864 40009 599082
rect 40519 599046 40689 599080
rect 40587 598594 40621 598812
rect 39907 598496 40077 598530
rect 39975 597668 40009 597886
rect 40519 597850 40689 597884
rect 676938 453416 676972 453634
rect 677482 453318 677652 453352
rect 676870 452672 677040 452706
rect 677550 452490 677584 452708
rect 676938 452220 676972 452438
rect 677482 452122 677652 452156
rect 676870 451476 677040 451510
rect 677550 451294 677584 451512
rect 676938 451024 676972 451242
rect 677482 450926 677652 450960
rect 676870 450280 677040 450314
rect 677550 450098 677584 450316
rect 676938 449828 676972 450046
rect 677482 449730 677652 449764
rect 676870 449084 677040 449118
rect 677550 448902 677584 449120
rect 676938 448632 676972 448850
rect 677482 448534 677652 448568
rect 676870 447888 677040 447922
rect 677550 447706 677584 447924
rect 676938 447436 676972 447654
rect 677482 447338 677652 447372
rect 676870 446692 677040 446726
rect 677550 446510 677584 446728
rect 676938 446240 676972 446458
rect 677482 446142 677652 446176
rect 676870 445496 677040 445530
rect 677550 445314 677584 445532
rect 676938 445044 676972 445262
rect 677482 444946 677652 444980
rect 676870 444300 677040 444334
rect 677550 444118 677584 444336
rect 676938 443848 676972 444066
rect 677482 443750 677652 443784
rect 676870 443104 677040 443138
rect 677550 442922 677584 443140
rect 676938 442652 676972 442870
rect 677482 442554 677652 442588
rect 676870 441908 677040 441942
rect 677550 441726 677584 441944
rect 676938 441456 676972 441674
rect 677482 441358 677652 441392
rect 676870 440712 677040 440746
rect 677550 440530 677584 440748
rect 676938 440260 676972 440478
rect 677482 440162 677652 440196
rect 676870 439516 677040 439550
rect 677550 439334 677584 439552
rect 40609 352373 40643 352591
rect 39929 352275 40099 352309
rect 39997 351447 40031 351665
rect 40541 351629 40711 351663
rect 40609 351177 40643 351395
rect 39929 351079 40099 351113
rect 39997 350251 40031 350469
rect 40541 350433 40711 350467
rect 40609 349981 40643 350199
rect 39929 349883 40099 349917
rect 39997 349055 40031 349273
rect 40541 349237 40711 349271
rect 40609 348785 40643 349003
rect 39929 348687 40099 348721
rect 39997 347859 40031 348077
rect 40541 348041 40711 348075
rect 40609 347589 40643 347807
rect 39929 347491 40099 347525
rect 39997 346663 40031 346881
rect 40541 346845 40711 346879
rect 40609 346393 40643 346611
rect 39929 346295 40099 346329
rect 39997 345467 40031 345685
rect 40541 345649 40711 345683
rect 40609 345197 40643 345415
rect 39929 345099 40099 345133
rect 39997 344271 40031 344489
rect 40541 344453 40711 344487
rect 40609 344001 40643 344219
rect 39929 343903 40099 343937
rect 39997 343075 40031 343293
rect 40541 343257 40711 343291
rect 40609 342805 40643 343023
rect 39929 342707 40099 342741
rect 39997 341879 40031 342097
rect 40541 342061 40711 342095
rect 40609 341609 40643 341827
rect 39929 341511 40099 341545
rect 39997 340683 40031 340901
rect 40541 340865 40711 340899
rect 40609 340413 40643 340631
rect 39929 340315 40099 340349
rect 39997 339487 40031 339705
rect 40541 339669 40711 339703
rect 40609 339217 40643 339435
rect 39929 339119 40099 339153
rect 39997 338291 40031 338509
rect 40541 338473 40711 338507
rect 40609 338021 40643 338239
rect 39929 337923 40099 337957
rect 39997 337095 40031 337313
rect 40541 337277 40711 337311
rect 40609 336825 40643 337043
rect 39929 336727 40099 336761
rect 39997 335899 40031 336117
rect 40541 336081 40711 336115
rect 40609 335629 40643 335847
rect 39929 335531 40099 335565
rect 39997 334703 40031 334921
rect 40541 334885 40711 334919
rect 134104 223102 134138 223272
rect 134848 223170 135066 223204
rect 135300 223102 135334 223272
rect 136044 223170 136262 223204
rect 136496 223102 136530 223272
rect 137240 223170 137458 223204
rect 137692 223102 137726 223272
rect 138436 223170 138654 223204
rect 138888 223102 138922 223272
rect 139632 223170 139850 223204
rect 140084 223102 140118 223272
rect 140828 223170 141046 223204
rect 141280 223102 141314 223272
rect 142024 223170 142242 223204
rect 142476 223102 142510 223272
rect 143220 223170 143438 223204
rect 143672 223102 143706 223272
rect 144416 223170 144634 223204
rect 144868 223102 144902 223272
rect 145612 223170 145830 223204
rect 146064 223102 146098 223272
rect 146808 223170 147026 223204
rect 147260 223102 147294 223272
rect 148004 223170 148222 223204
rect 148456 223102 148490 223272
rect 149200 223170 149418 223204
rect 149652 223102 149686 223272
rect 150396 223170 150614 223204
rect 150848 223102 150882 223272
rect 151592 223170 151810 223204
rect 152044 223102 152078 223272
rect 152788 223170 153006 223204
rect 153240 223102 153274 223272
rect 153984 223170 154202 223204
rect 154436 223102 154470 223272
rect 155180 223170 155398 223204
rect 155632 223102 155666 223272
rect 156376 223170 156594 223204
rect 156828 223102 156862 223272
rect 157572 223170 157790 223204
rect 158024 223102 158058 223272
rect 158768 223170 158986 223204
rect 394104 223102 394138 223272
rect 394848 223170 395066 223204
rect 395300 223102 395334 223272
rect 396044 223170 396262 223204
rect 396496 223102 396530 223272
rect 397240 223170 397458 223204
rect 397692 223102 397726 223272
rect 398436 223170 398654 223204
rect 398888 223102 398922 223272
rect 399632 223170 399850 223204
rect 400084 223102 400118 223272
rect 400828 223170 401046 223204
rect 401280 223102 401314 223272
rect 402024 223170 402242 223204
rect 402476 223102 402510 223272
rect 403220 223170 403438 223204
rect 403672 223102 403706 223272
rect 404416 223170 404634 223204
rect 404868 223102 404902 223272
rect 405612 223170 405830 223204
rect 406064 223102 406098 223272
rect 406808 223170 407026 223204
rect 407260 223102 407294 223272
rect 408004 223170 408222 223204
rect 408456 223102 408490 223272
rect 409200 223170 409418 223204
rect 409652 223102 409686 223272
rect 410396 223170 410614 223204
rect 410848 223102 410882 223272
rect 411592 223170 411810 223204
rect 412044 223102 412078 223272
rect 412788 223170 413006 223204
rect 413240 223102 413274 223272
rect 413984 223170 414202 223204
rect 414436 223102 414470 223272
rect 415180 223170 415398 223204
rect 415632 223102 415666 223272
rect 416376 223170 416594 223204
rect 416828 223102 416862 223272
rect 417572 223170 417790 223204
rect 418024 223102 418058 223272
rect 418768 223170 418986 223204
rect 135118 222558 135336 222592
rect 135946 222490 135980 222660
rect 136314 222558 136532 222592
rect 137142 222490 137176 222660
rect 137510 222558 137728 222592
rect 138338 222490 138372 222660
rect 138706 222558 138924 222592
rect 139534 222490 139568 222660
rect 139902 222558 140120 222592
rect 140730 222490 140764 222660
rect 141098 222558 141316 222592
rect 141926 222490 141960 222660
rect 142294 222558 142512 222592
rect 143122 222490 143156 222660
rect 143490 222558 143708 222592
rect 144318 222490 144352 222660
rect 144686 222558 144904 222592
rect 145514 222490 145548 222660
rect 145882 222558 146100 222592
rect 146710 222490 146744 222660
rect 147078 222558 147296 222592
rect 147906 222490 147940 222660
rect 148274 222558 148492 222592
rect 149102 222490 149136 222660
rect 149470 222558 149688 222592
rect 150298 222490 150332 222660
rect 150666 222558 150884 222592
rect 151494 222490 151528 222660
rect 151862 222558 152080 222592
rect 152690 222490 152724 222660
rect 153058 222558 153276 222592
rect 153886 222490 153920 222660
rect 154254 222558 154472 222592
rect 155082 222490 155116 222660
rect 155450 222558 155668 222592
rect 156278 222490 156312 222660
rect 156646 222558 156864 222592
rect 157474 222490 157508 222660
rect 158024 222490 158058 222660
rect 158668 222558 158886 222592
rect 395118 222558 395336 222592
rect 395946 222490 395980 222660
rect 396314 222558 396532 222592
rect 397142 222490 397176 222660
rect 397510 222558 397728 222592
rect 398338 222490 398372 222660
rect 398706 222558 398924 222592
rect 399534 222490 399568 222660
rect 399902 222558 400120 222592
rect 400730 222490 400764 222660
rect 401098 222558 401316 222592
rect 401926 222490 401960 222660
rect 402294 222558 402512 222592
rect 403122 222490 403156 222660
rect 403490 222558 403708 222592
rect 404318 222490 404352 222660
rect 404686 222558 404904 222592
rect 405514 222490 405548 222660
rect 405882 222558 406100 222592
rect 406710 222490 406744 222660
rect 407078 222558 407296 222592
rect 407906 222490 407940 222660
rect 408274 222558 408492 222592
rect 409102 222490 409136 222660
rect 409470 222558 409688 222592
rect 410298 222490 410332 222660
rect 410666 222558 410884 222592
rect 411494 222490 411528 222660
rect 411862 222558 412080 222592
rect 412690 222490 412724 222660
rect 413058 222558 413276 222592
rect 413886 222490 413920 222660
rect 414254 222558 414472 222592
rect 415082 222490 415116 222660
rect 415450 222558 415668 222592
rect 416278 222490 416312 222660
rect 416646 222558 416864 222592
rect 417474 222490 417508 222660
rect 418024 222490 418058 222660
rect 418668 222558 418886 222592
<< metal1 >>
rect 416862 997387 416914 997399
rect 417502 997275 417514 997327
rect 417732 997275 417744 997327
rect 662863 997305 662915 997317
rect 416862 997205 416914 997217
rect 664059 997305 664111 997317
rect 663503 997193 663515 997245
rect 663733 997193 663745 997245
rect 662863 997123 662915 997135
rect 665255 997305 665307 997317
rect 664699 997193 664711 997245
rect 664929 997193 664941 997245
rect 664059 997123 664111 997135
rect 666451 997305 666503 997317
rect 665895 997193 665907 997245
rect 666125 997193 666137 997245
rect 665255 997123 665307 997135
rect 667091 997193 667103 997245
rect 667321 997193 667333 997245
rect 666451 997123 666503 997135
rect 167870 997062 167922 997074
rect 167040 996950 167052 997002
rect 167270 996950 167282 997002
rect 169066 997062 169118 997074
rect 168236 996950 168248 997002
rect 168466 996950 168478 997002
rect 167870 996880 167922 996892
rect 170262 997062 170314 997074
rect 169432 996950 169444 997002
rect 169662 996950 169674 997002
rect 169066 996880 169118 996892
rect 417844 997026 418598 997044
rect 417844 996966 418223 997026
rect 418580 996966 418598 997026
rect 417844 996948 418598 996966
rect 170262 996880 170314 996892
rect 417508 996775 417560 996787
rect 416576 996663 416588 996715
rect 416806 996663 416818 996715
rect 663509 996693 663561 996705
rect 417508 996593 417560 996605
rect 662577 996581 662589 996633
rect 662807 996581 662819 996633
rect 664705 996693 664757 996705
rect 663773 996581 663785 996633
rect 664003 996581 664015 996633
rect 663509 996511 663561 996523
rect 665901 996693 665953 996705
rect 664969 996581 664981 996633
rect 665199 996581 665211 996633
rect 664705 996511 664757 996523
rect 667097 996693 667149 996705
rect 666165 996581 666177 996633
rect 666395 996581 666407 996633
rect 665901 996511 665953 996523
rect 667097 996511 667149 996523
rect 167224 996450 167276 996462
rect 168420 996450 168472 996462
rect 167966 996338 167978 996390
rect 168196 996338 168208 996390
rect 167224 996268 167276 996280
rect 169616 996450 169668 996462
rect 169162 996338 169174 996390
rect 169392 996338 169404 996390
rect 168420 996268 168472 996280
rect 170358 996338 170370 996390
rect 170588 996338 170600 996390
rect 169616 996268 169668 996280
rect 42491 995429 169626 995457
rect 40554 891418 40606 891430
rect 42491 891357 42519 995429
rect 169620 995405 169626 995429
rect 169678 995405 169684 995457
rect 170463 995401 170469 995453
rect 170521 995429 170527 995453
rect 170521 995401 172109 995429
rect 42467 891351 42519 891357
rect 42467 891293 42519 891299
rect 42547 995373 169502 995401
rect 40554 891188 40606 891200
rect 42547 891163 42575 995373
rect 169496 995349 169502 995373
rect 169554 995349 169560 995401
rect 170269 995345 170275 995397
rect 170327 995373 170333 995397
rect 170327 995345 171909 995373
rect 42523 891157 42575 891163
rect 39870 891092 39882 891144
rect 40052 891092 40064 891144
rect 42523 891099 42575 891105
rect 42603 995317 168430 995345
rect 42463 890508 42515 890514
rect 39942 890492 39994 890504
rect 40482 890446 40494 890498
rect 40664 890446 40676 890498
rect 42463 890450 42515 890456
rect 39942 890262 39994 890274
rect 40554 890222 40606 890234
rect 40554 889992 40606 890004
rect 39870 889896 39882 889948
rect 40052 889896 40064 889948
rect 39942 889296 39994 889308
rect 40482 889250 40494 889302
rect 40664 889250 40676 889302
rect 39942 889066 39994 889078
rect 40554 889026 40606 889038
rect 40554 888796 40606 888808
rect 39870 888700 39882 888752
rect 40052 888700 40064 888752
rect 39942 888100 39994 888112
rect 40482 888054 40494 888106
rect 40664 888054 40676 888106
rect 39942 887870 39994 887882
rect 40554 887830 40606 887842
rect 40554 887600 40606 887612
rect 39870 887504 39882 887556
rect 40052 887504 40064 887556
rect 39942 886904 39994 886916
rect 40482 886858 40494 886910
rect 40664 886858 40676 886910
rect 39942 886674 39994 886686
rect 40554 886634 40606 886646
rect 40554 886404 40606 886416
rect 39870 886308 39882 886360
rect 40052 886308 40064 886360
rect 39942 885708 39994 885720
rect 40482 885662 40494 885714
rect 40664 885662 40676 885714
rect 39942 885478 39994 885490
rect 40579 610772 40631 610784
rect 42463 610711 42491 890450
rect 42439 610705 42491 610711
rect 42439 610647 42491 610653
rect 42519 890384 42571 890390
rect 42519 890326 42571 890332
rect 40579 610542 40631 610554
rect 42519 610517 42547 890326
rect 42603 890137 42631 995317
rect 168424 995293 168430 995317
rect 168482 995293 168488 995345
rect 169243 995289 169249 995341
rect 169301 995317 169307 995341
rect 169301 995289 171711 995317
rect 42579 890131 42631 890137
rect 42579 890073 42631 890079
rect 42659 995261 168306 995289
rect 42659 889967 42687 995261
rect 168300 995237 168306 995261
rect 168358 995237 168364 995289
rect 169073 995233 169079 995285
rect 169131 995261 169137 995285
rect 169131 995233 171511 995261
rect 416649 995247 416655 995271
rect 42635 889961 42687 889967
rect 42635 889903 42687 889909
rect 42715 995205 167234 995233
rect 42495 610511 42547 610517
rect 39895 610446 39907 610498
rect 40077 610446 40089 610498
rect 42495 610453 42547 610459
rect 42575 889312 42627 889318
rect 42575 889254 42627 889260
rect 42435 609862 42487 609868
rect 39967 609846 40019 609858
rect 40507 609800 40519 609852
rect 40689 609800 40701 609852
rect 42435 609804 42487 609810
rect 39967 609616 40019 609628
rect 40579 609576 40631 609588
rect 40579 609346 40631 609358
rect 39895 609250 39907 609302
rect 40077 609250 40089 609302
rect 39967 608650 40019 608662
rect 40507 608604 40519 608656
rect 40689 608604 40701 608656
rect 39967 608420 40019 608432
rect 40579 608380 40631 608392
rect 40579 608150 40631 608162
rect 39895 608054 39907 608106
rect 40077 608054 40089 608106
rect 39967 607454 40019 607466
rect 40507 607408 40519 607460
rect 40689 607408 40701 607460
rect 39967 607224 40019 607236
rect 40579 607184 40631 607196
rect 40579 606954 40631 606966
rect 39895 606858 39907 606910
rect 40077 606858 40089 606910
rect 39967 606258 40019 606270
rect 40507 606212 40519 606264
rect 40689 606212 40701 606264
rect 39967 606028 40019 606040
rect 40579 605988 40631 606000
rect 40579 605758 40631 605770
rect 39895 605662 39907 605714
rect 40077 605662 40089 605714
rect 39967 605062 40019 605074
rect 40507 605016 40519 605068
rect 40689 605016 40701 605068
rect 39967 604832 40019 604844
rect 40579 604792 40631 604804
rect 40579 604562 40631 604574
rect 39895 604466 39907 604518
rect 40077 604466 40089 604518
rect 39967 603866 40019 603878
rect 40507 603820 40519 603872
rect 40689 603820 40701 603872
rect 39967 603636 40019 603648
rect 40579 603596 40631 603608
rect 40579 603366 40631 603378
rect 39895 603270 39907 603322
rect 40077 603270 40089 603322
rect 39967 602670 40019 602682
rect 40507 602624 40519 602676
rect 40689 602624 40701 602676
rect 39967 602440 40019 602452
rect 40579 602400 40631 602412
rect 40579 602170 40631 602182
rect 39895 602074 39907 602126
rect 40077 602074 40089 602126
rect 39967 601474 40019 601486
rect 40507 601428 40519 601480
rect 40689 601428 40701 601480
rect 39967 601244 40019 601256
rect 40579 601204 40631 601216
rect 40579 600974 40631 600986
rect 39895 600878 39907 600930
rect 40077 600878 40089 600930
rect 39967 600278 40019 600290
rect 40507 600232 40519 600284
rect 40689 600232 40701 600284
rect 39967 600048 40019 600060
rect 40579 600008 40631 600020
rect 40579 599778 40631 599790
rect 39895 599682 39907 599734
rect 40077 599682 40089 599734
rect 39967 599082 40019 599094
rect 40507 599036 40519 599088
rect 40689 599036 40701 599088
rect 39967 598852 40019 598864
rect 40579 598812 40631 598824
rect 40579 598582 40631 598594
rect 39895 598486 39907 598538
rect 40077 598486 40089 598538
rect 39967 597886 40019 597898
rect 40507 597840 40519 597892
rect 40689 597840 40701 597892
rect 39967 597656 40019 597668
rect 40601 352591 40653 352603
rect 42435 352530 42463 609804
rect 42411 352524 42463 352530
rect 42411 352466 42463 352472
rect 42491 609738 42543 609744
rect 42491 609680 42543 609686
rect 40601 352361 40653 352373
rect 42491 352336 42519 609680
rect 42575 609491 42603 889254
rect 42551 609485 42603 609491
rect 42551 609427 42603 609433
rect 42631 889188 42683 889194
rect 42631 889130 42683 889136
rect 42631 609321 42659 889130
rect 42715 888965 42743 995205
rect 167228 995181 167234 995205
rect 167286 995181 167292 995233
rect 168071 995177 168077 995229
rect 168129 995205 168135 995229
rect 415907 995219 416655 995247
rect 416707 995219 416713 995271
rect 417492 995223 417498 995275
rect 417550 995247 661880 995275
rect 662650 995247 662656 995271
rect 417550 995223 417556 995247
rect 661842 995219 662656 995247
rect 662708 995219 662714 995271
rect 663493 995223 663499 995275
rect 663551 995247 675148 995275
rect 663551 995223 663557 995247
rect 168129 995177 171310 995205
rect 416843 995191 416849 995215
rect 42691 888959 42743 888965
rect 42691 888901 42743 888907
rect 42771 995149 167110 995177
rect 42771 888771 42799 995149
rect 167104 995125 167110 995149
rect 167162 995125 167168 995177
rect 167877 995121 167883 995173
rect 167935 995149 167941 995173
rect 416107 995163 416849 995191
rect 416901 995163 416907 995215
rect 417611 995191 417622 995219
rect 417616 995167 417622 995191
rect 417674 995191 661762 995219
rect 662844 995191 662850 995215
rect 417674 995167 417680 995191
rect 661725 995163 662850 995191
rect 662902 995163 662908 995215
rect 663617 995167 663623 995219
rect 663675 995191 675092 995219
rect 663675 995167 663681 995191
rect 167935 995121 171110 995149
rect 663846 995135 663852 995159
rect 660923 995107 663852 995135
rect 663904 995107 663910 995159
rect 664689 995111 664695 995163
rect 664747 995135 675036 995163
rect 664747 995111 664753 995135
rect 664040 995079 664046 995103
rect 661123 995051 664046 995079
rect 664098 995051 664104 995103
rect 664813 995055 664819 995107
rect 664871 995079 674980 995107
rect 664871 995055 664877 995079
rect 665042 995023 665048 995047
rect 661323 994995 665048 995023
rect 665100 994995 665106 995047
rect 665885 994999 665891 995051
rect 665943 995023 674924 995051
rect 665943 994999 665949 995023
rect 665236 994967 665242 994991
rect 661523 994939 665242 994967
rect 665294 994939 665300 994991
rect 666009 994943 666015 994995
rect 666067 994967 674868 994995
rect 666067 994943 666073 994967
rect 666238 994911 666244 994935
rect 661723 994883 666244 994911
rect 666296 994883 666302 994935
rect 667081 994887 667087 994939
rect 667139 994911 674812 994939
rect 667139 994887 667145 994911
rect 666432 994855 666438 994879
rect 661923 994827 666438 994855
rect 666490 994827 666496 994879
rect 667200 994855 667211 994883
rect 667205 994831 667211 994855
rect 667263 994855 674756 994883
rect 667263 994831 667269 994855
rect 42747 888765 42799 888771
rect 42747 888707 42799 888713
rect 42607 609315 42659 609321
rect 42607 609257 42659 609263
rect 42687 888116 42739 888122
rect 42687 888058 42739 888064
rect 42467 352330 42519 352336
rect 39917 352265 39929 352317
rect 40099 352265 40111 352317
rect 42467 352272 42519 352278
rect 42547 608666 42599 608672
rect 42547 608608 42599 608614
rect 42407 351681 42459 351687
rect 39989 351665 40041 351677
rect 40529 351619 40541 351671
rect 40711 351619 40723 351671
rect 42407 351623 42459 351629
rect 39989 351435 40041 351447
rect 40601 351395 40653 351407
rect 40601 351165 40653 351177
rect 39917 351069 39929 351121
rect 40099 351069 40111 351121
rect 39989 350469 40041 350481
rect 40529 350423 40541 350475
rect 40711 350423 40723 350475
rect 39989 350239 40041 350251
rect 40601 350199 40653 350211
rect 40601 349969 40653 349981
rect 39917 349873 39929 349925
rect 40099 349873 40111 349925
rect 39989 349273 40041 349285
rect 40529 349227 40541 349279
rect 40711 349227 40723 349279
rect 39989 349043 40041 349055
rect 40601 349003 40653 349015
rect 40601 348773 40653 348785
rect 39917 348677 39929 348729
rect 40099 348677 40111 348729
rect 39989 348077 40041 348089
rect 40529 348031 40541 348083
rect 40711 348031 40723 348083
rect 39989 347847 40041 347859
rect 40601 347807 40653 347819
rect 40601 347577 40653 347589
rect 39917 347481 39929 347533
rect 40099 347481 40111 347533
rect 39989 346881 40041 346893
rect 40529 346835 40541 346887
rect 40711 346835 40723 346887
rect 39989 346651 40041 346663
rect 40601 346611 40653 346623
rect 40601 346381 40653 346393
rect 39917 346285 39929 346337
rect 40099 346285 40111 346337
rect 39989 345685 40041 345697
rect 40529 345639 40541 345691
rect 40711 345639 40723 345691
rect 39989 345455 40041 345467
rect 40601 345415 40653 345427
rect 40601 345185 40653 345197
rect 39917 345089 39929 345141
rect 40099 345089 40111 345141
rect 39989 344489 40041 344501
rect 40529 344443 40541 344495
rect 40711 344443 40723 344495
rect 39989 344259 40041 344271
rect 40601 344219 40653 344231
rect 40601 343989 40653 344001
rect 39917 343893 39929 343945
rect 40099 343893 40111 343945
rect 39989 343293 40041 343305
rect 40529 343247 40541 343299
rect 40711 343247 40723 343299
rect 39989 343063 40041 343075
rect 40601 343023 40653 343035
rect 40601 342793 40653 342805
rect 39917 342697 39929 342749
rect 40099 342697 40111 342749
rect 39989 342097 40041 342109
rect 40529 342051 40541 342103
rect 40711 342051 40723 342103
rect 39989 341867 40041 341879
rect 40601 341827 40653 341839
rect 40601 341597 40653 341609
rect 39917 341501 39929 341553
rect 40099 341501 40111 341553
rect 39989 340901 40041 340913
rect 40529 340855 40541 340907
rect 40711 340855 40723 340907
rect 39989 340671 40041 340683
rect 40601 340631 40653 340643
rect 40601 340401 40653 340413
rect 39917 340305 39929 340357
rect 40099 340305 40111 340357
rect 39989 339705 40041 339717
rect 40529 339659 40541 339711
rect 40711 339659 40723 339711
rect 39989 339475 40041 339487
rect 40601 339435 40653 339447
rect 40601 339205 40653 339217
rect 39917 339109 39929 339161
rect 40099 339109 40111 339161
rect 39989 338509 40041 338521
rect 40529 338463 40541 338515
rect 40711 338463 40723 338515
rect 39989 338279 40041 338291
rect 40601 338239 40653 338251
rect 40601 338009 40653 338021
rect 39917 337913 39929 337965
rect 40099 337913 40111 337965
rect 39989 337313 40041 337325
rect 40529 337267 40541 337319
rect 40711 337267 40723 337319
rect 39989 337083 40041 337095
rect 40601 337043 40653 337055
rect 40601 336813 40653 336825
rect 39917 336717 39929 336769
rect 40099 336717 40111 336769
rect 39989 336117 40041 336129
rect 40529 336071 40541 336123
rect 40711 336071 40723 336123
rect 39989 335887 40041 335899
rect 40601 335847 40653 335859
rect 40601 335617 40653 335629
rect 39917 335521 39929 335573
rect 40099 335521 40111 335573
rect 39989 334921 40041 334933
rect 40529 334875 40541 334927
rect 40711 334875 40723 334927
rect 39989 334691 40041 334703
rect 42407 224252 42435 351623
rect 42463 351557 42515 351563
rect 42463 351499 42515 351505
rect 42463 224308 42491 351499
rect 42547 351310 42575 608608
rect 42523 351304 42575 351310
rect 42523 351246 42575 351252
rect 42603 608542 42655 608548
rect 42603 608484 42655 608490
rect 42603 351140 42631 608484
rect 42687 608319 42715 888058
rect 42663 608313 42715 608319
rect 42663 608255 42715 608261
rect 42743 887992 42795 887998
rect 42743 887934 42795 887940
rect 42743 608125 42771 887934
rect 42827 887745 42855 892517
rect 42803 887739 42855 887745
rect 42803 887681 42855 887687
rect 42883 887575 42911 892317
rect 42859 887569 42911 887575
rect 42859 887511 42911 887517
rect 42719 608119 42771 608125
rect 42719 608061 42771 608067
rect 42799 886920 42851 886926
rect 42799 886862 42851 886868
rect 42579 351134 42631 351140
rect 42579 351076 42631 351082
rect 42659 607470 42711 607476
rect 42659 607412 42711 607418
rect 42519 350485 42571 350491
rect 42519 350427 42571 350433
rect 42519 224364 42547 350427
rect 42575 350361 42627 350367
rect 42575 350303 42627 350309
rect 42575 224420 42603 350303
rect 42659 350138 42687 607412
rect 42635 350132 42687 350138
rect 42635 350074 42687 350080
rect 42715 607346 42767 607352
rect 42715 607288 42767 607294
rect 42715 349944 42743 607288
rect 42799 607099 42827 886862
rect 42775 607093 42827 607099
rect 42775 607035 42827 607041
rect 42855 886796 42907 886802
rect 42855 886738 42907 886744
rect 42855 606929 42883 886738
rect 42939 886573 42967 892117
rect 42915 886567 42967 886573
rect 42915 886509 42967 886515
rect 42995 886379 43023 891917
rect 42971 886373 43023 886379
rect 42971 886315 43023 886321
rect 42831 606923 42883 606929
rect 42831 606865 42883 606871
rect 42911 885724 42963 885730
rect 42911 885666 42963 885672
rect 42691 349938 42743 349944
rect 42691 349880 42743 349886
rect 42771 606274 42823 606280
rect 42771 606216 42823 606222
rect 42631 349289 42683 349295
rect 42631 349231 42683 349237
rect 42631 224476 42659 349231
rect 42687 349165 42739 349171
rect 42687 349107 42739 349113
rect 42687 224532 42715 349107
rect 42771 348918 42799 606216
rect 42747 348912 42799 348918
rect 42747 348854 42799 348860
rect 42827 606150 42879 606156
rect 42827 606092 42879 606098
rect 42827 348748 42855 606092
rect 42911 605927 42939 885666
rect 42887 605921 42939 605927
rect 42887 605863 42939 605869
rect 42967 885600 43019 885606
rect 42967 885542 43019 885548
rect 42967 605733 42995 885542
rect 674728 715999 674756 994855
rect 674700 715963 674756 715999
rect 674476 708223 674504 714921
rect 674532 708417 674560 715121
rect 674588 709419 674616 715321
rect 674644 709613 674672 715521
rect 674700 710615 674728 715963
rect 674784 715872 674812 994911
rect 674756 715836 674812 715872
rect 674756 710809 674784 715836
rect 674840 715738 674868 994967
rect 674812 715703 674868 715738
rect 674812 711811 674840 715703
rect 674896 715598 674924 995023
rect 674868 715562 674924 715598
rect 674868 712005 674896 715562
rect 674952 715461 674980 995079
rect 674924 715425 674980 715461
rect 674924 713007 674952 715425
rect 675008 715315 675036 995135
rect 674980 715278 675036 715315
rect 674980 713201 675008 715278
rect 675064 715186 675092 995191
rect 675036 715151 675092 715186
rect 675036 714203 675064 715151
rect 675120 715077 675148 995247
rect 675092 715042 675148 715077
rect 675092 714373 675120 715042
rect 676928 714458 676980 714470
rect 675092 714367 675144 714373
rect 675092 714309 675144 714315
rect 676928 714228 676980 714240
rect 675036 714197 675088 714203
rect 675036 714139 675088 714145
rect 677470 714132 677482 714184
rect 677652 714132 677664 714184
rect 675096 713548 675148 713554
rect 675096 713490 675148 713496
rect 675040 713424 675092 713430
rect 675040 713366 675092 713372
rect 674980 713195 675032 713201
rect 674980 713137 675032 713143
rect 674924 713001 674976 713007
rect 674924 712943 674976 712949
rect 674984 712352 675036 712358
rect 674984 712294 675036 712300
rect 674928 712228 674980 712234
rect 674928 712170 674980 712176
rect 674868 711999 674920 712005
rect 674868 711941 674920 711947
rect 674812 711805 674864 711811
rect 674812 711747 674864 711753
rect 674872 711156 674924 711162
rect 674872 711098 674924 711104
rect 674816 711032 674868 711038
rect 674816 710974 674868 710980
rect 674756 710803 674808 710809
rect 674756 710745 674808 710751
rect 674700 710609 674752 710615
rect 674700 710551 674752 710557
rect 674760 709960 674812 709966
rect 674760 709902 674812 709908
rect 674704 709836 674756 709842
rect 674704 709778 674756 709784
rect 674644 709607 674696 709613
rect 674644 709549 674696 709555
rect 674588 709413 674640 709419
rect 674588 709355 674640 709361
rect 674648 708764 674700 708770
rect 674648 708706 674700 708712
rect 674592 708640 674644 708646
rect 674592 708582 674644 708588
rect 674532 708411 674584 708417
rect 674532 708353 674584 708359
rect 674476 708217 674528 708223
rect 674476 708159 674528 708165
rect 674536 707568 674588 707574
rect 674536 707510 674588 707516
rect 674504 707450 674532 707455
rect 674480 707444 674532 707450
rect 674480 707386 674532 707392
rect 42943 605727 42995 605733
rect 42943 605669 42995 605675
rect 42803 348742 42855 348748
rect 42803 348684 42855 348690
rect 42883 605078 42935 605084
rect 42883 605020 42935 605026
rect 42743 348093 42795 348099
rect 42743 348035 42795 348041
rect 42743 224588 42771 348035
rect 42799 347969 42851 347975
rect 42799 347911 42851 347917
rect 42799 224644 42827 347911
rect 42883 347746 42911 605020
rect 42859 347740 42911 347746
rect 42859 347682 42911 347688
rect 42939 604954 42991 604960
rect 42939 604896 42991 604902
rect 42939 347552 42967 604896
rect 43023 604731 43051 613556
rect 42999 604725 43051 604731
rect 42999 604667 43051 604673
rect 43079 604537 43107 613356
rect 43055 604531 43107 604537
rect 43055 604473 43107 604479
rect 42915 347546 42967 347552
rect 42915 347488 42967 347494
rect 42995 603882 43047 603888
rect 42995 603824 43047 603830
rect 42855 346897 42907 346903
rect 42855 346839 42907 346845
rect 42855 224700 42883 346839
rect 42911 346773 42963 346779
rect 42911 346715 42963 346721
rect 42911 224756 42939 346715
rect 42995 346550 43023 603824
rect 42971 346544 43023 346550
rect 42971 346486 43023 346492
rect 43051 603758 43103 603764
rect 43051 603700 43103 603706
rect 43051 346356 43079 603700
rect 43135 603535 43163 613156
rect 43111 603529 43163 603535
rect 43111 603471 43163 603477
rect 43191 603341 43219 612956
rect 43167 603335 43219 603341
rect 43167 603277 43219 603283
rect 43027 346350 43079 346356
rect 43027 346292 43079 346298
rect 43107 602686 43159 602692
rect 43107 602628 43159 602634
rect 42967 345701 43019 345707
rect 42967 345643 43019 345649
rect 42967 224812 42995 345643
rect 43023 345577 43075 345583
rect 43023 345519 43075 345525
rect 43023 224868 43051 345519
rect 43107 345354 43135 602628
rect 43083 345348 43135 345354
rect 43083 345290 43135 345296
rect 43163 602562 43215 602568
rect 43163 602504 43215 602510
rect 43163 345160 43191 602504
rect 43247 602339 43275 612756
rect 43223 602333 43275 602339
rect 43223 602275 43275 602281
rect 43303 602145 43331 612556
rect 43279 602139 43331 602145
rect 43279 602081 43331 602087
rect 43139 345154 43191 345160
rect 43139 345096 43191 345102
rect 43219 601490 43271 601496
rect 43219 601432 43271 601438
rect 43079 344505 43131 344511
rect 43079 344447 43131 344453
rect 43079 224924 43107 344447
rect 43135 344381 43187 344387
rect 43135 344323 43187 344329
rect 43135 224980 43163 344323
rect 43219 344158 43247 601432
rect 43195 344152 43247 344158
rect 43195 344094 43247 344100
rect 43275 601366 43327 601372
rect 43275 601308 43327 601314
rect 43275 343964 43303 601308
rect 43359 601143 43387 612356
rect 43335 601137 43387 601143
rect 43335 601079 43387 601085
rect 43415 600949 43443 612156
rect 43391 600943 43443 600949
rect 43391 600885 43443 600891
rect 43251 343958 43303 343964
rect 43251 343900 43303 343906
rect 43331 600294 43383 600300
rect 43331 600236 43383 600242
rect 43191 343309 43243 343315
rect 43191 343251 43243 343257
rect 43191 225036 43219 343251
rect 43247 343185 43299 343191
rect 43247 343127 43299 343133
rect 43247 225092 43275 343127
rect 43331 342962 43359 600236
rect 43307 342956 43359 342962
rect 43307 342898 43359 342904
rect 43387 600170 43439 600176
rect 43387 600112 43439 600118
rect 43387 342768 43415 600112
rect 43471 599947 43499 611956
rect 43447 599941 43499 599947
rect 43447 599883 43499 599889
rect 43527 599753 43555 611756
rect 43503 599747 43555 599753
rect 43503 599689 43555 599695
rect 43363 342762 43415 342768
rect 43363 342704 43415 342710
rect 43443 599098 43495 599104
rect 43443 599040 43495 599046
rect 43303 342113 43355 342119
rect 43303 342055 43355 342061
rect 43303 225148 43331 342055
rect 43359 341989 43411 341995
rect 43359 341931 43411 341937
rect 43359 225204 43387 341931
rect 43443 341766 43471 599040
rect 43419 341760 43471 341766
rect 43419 341702 43471 341708
rect 43499 598974 43551 598980
rect 43499 598916 43551 598922
rect 43499 341572 43527 598916
rect 43583 598751 43611 611556
rect 43559 598745 43611 598751
rect 43559 598687 43611 598693
rect 43639 598557 43667 611356
rect 43615 598551 43667 598557
rect 43615 598493 43667 598499
rect 43475 341566 43527 341572
rect 43475 341508 43527 341514
rect 43555 597902 43607 597908
rect 43555 597844 43607 597850
rect 43415 340917 43467 340923
rect 43415 340859 43467 340865
rect 43415 225260 43443 340859
rect 43471 340793 43523 340799
rect 43471 340735 43523 340741
rect 43471 225316 43499 340735
rect 43555 340570 43583 597844
rect 43531 340564 43583 340570
rect 43531 340506 43583 340512
rect 43611 597778 43663 597784
rect 43611 597720 43663 597726
rect 43611 340376 43639 597720
rect 673804 440223 673832 454055
rect 673860 440417 673888 454255
rect 673916 441419 673944 454455
rect 673972 441613 674000 454655
rect 674028 442615 674056 454855
rect 674084 442809 674112 455055
rect 674140 443811 674168 455255
rect 674196 444005 674224 455455
rect 674252 445007 674280 455655
rect 674308 445201 674336 455855
rect 674364 446203 674392 456055
rect 674420 446397 674448 456255
rect 674504 455108 674532 707386
rect 674476 455079 674532 455108
rect 674476 447399 674504 455079
rect 674560 455050 674588 707510
rect 674532 455020 674588 455050
rect 674532 447593 674560 455020
rect 674616 454991 674644 708582
rect 674588 454963 674644 454991
rect 674588 448595 674616 454963
rect 674672 454931 674700 708706
rect 674644 454898 674700 454931
rect 674644 448789 674672 454898
rect 674728 454866 674756 709778
rect 674700 454836 674756 454866
rect 674700 449791 674728 454836
rect 674784 454805 674812 709902
rect 674756 454769 674812 454805
rect 674756 449961 674784 454769
rect 674840 454733 674868 710974
rect 674812 454699 674868 454733
rect 674812 450987 674840 454699
rect 674896 454666 674924 711098
rect 674868 454635 674924 454666
rect 674868 451181 674896 454635
rect 674952 454606 674980 712170
rect 674924 454573 674980 454606
rect 674924 452183 674952 454573
rect 675008 454544 675036 712294
rect 674980 454501 675036 454544
rect 674980 452353 675008 454501
rect 675064 454472 675092 713366
rect 675036 454432 675092 454472
rect 675036 453379 675064 454432
rect 675120 454403 675148 713490
rect 676858 713486 676870 713538
rect 677040 713486 677052 713538
rect 677540 713532 677592 713544
rect 677540 713302 677592 713314
rect 676928 713262 676980 713274
rect 676928 713032 676980 713044
rect 677470 712936 677482 712988
rect 677652 712936 677664 712988
rect 676858 712290 676870 712342
rect 677040 712290 677052 712342
rect 677540 712336 677592 712348
rect 677540 712106 677592 712118
rect 676928 712066 676980 712078
rect 676928 711836 676980 711848
rect 677470 711740 677482 711792
rect 677652 711740 677664 711792
rect 676858 711094 676870 711146
rect 677040 711094 677052 711146
rect 677540 711140 677592 711152
rect 677540 710910 677592 710922
rect 676928 710870 676980 710882
rect 676928 710640 676980 710652
rect 677470 710544 677482 710596
rect 677652 710544 677664 710596
rect 676858 709898 676870 709950
rect 677040 709898 677052 709950
rect 677540 709944 677592 709956
rect 677540 709714 677592 709726
rect 676928 709674 676980 709686
rect 676928 709444 676980 709456
rect 677470 709348 677482 709400
rect 677652 709348 677664 709400
rect 676858 708702 676870 708754
rect 677040 708702 677052 708754
rect 677540 708748 677592 708760
rect 677540 708518 677592 708530
rect 676928 708478 676980 708490
rect 676928 708248 676980 708260
rect 677470 708152 677482 708204
rect 677652 708152 677664 708204
rect 676858 707506 676870 707558
rect 677040 707506 677052 707558
rect 677540 707552 677592 707564
rect 677540 707322 677592 707334
rect 675092 454365 675148 454403
rect 675092 453573 675120 454365
rect 676928 453634 676980 453646
rect 675092 453567 675144 453573
rect 675092 453509 675144 453515
rect 676928 453404 676980 453416
rect 675036 453373 675088 453379
rect 675036 453315 675088 453321
rect 677470 453308 677482 453360
rect 677652 453308 677664 453360
rect 675096 452724 675148 452730
rect 675096 452666 675148 452672
rect 675040 452600 675092 452606
rect 675040 452542 675092 452548
rect 674980 452347 675032 452353
rect 674980 452289 675032 452295
rect 674924 452177 674976 452183
rect 674924 452119 674976 452125
rect 674984 451528 675036 451534
rect 674984 451470 675036 451476
rect 674928 451404 674980 451410
rect 674928 451346 674980 451352
rect 674868 451175 674920 451181
rect 674868 451117 674920 451123
rect 674812 450981 674864 450987
rect 674812 450923 674864 450929
rect 674872 450332 674924 450338
rect 674872 450274 674924 450280
rect 674816 450208 674868 450214
rect 674816 450150 674868 450156
rect 674756 449955 674808 449961
rect 674756 449897 674808 449903
rect 674700 449785 674752 449791
rect 674700 449727 674752 449733
rect 674760 449136 674812 449142
rect 674760 449078 674812 449084
rect 674704 449012 674756 449018
rect 674704 448954 674756 448960
rect 674644 448783 674696 448789
rect 674644 448725 674696 448731
rect 674588 448589 674640 448595
rect 674588 448531 674640 448537
rect 674648 447940 674700 447946
rect 674648 447882 674700 447888
rect 674592 447816 674644 447822
rect 674592 447758 674644 447764
rect 674532 447587 674584 447593
rect 674532 447529 674584 447535
rect 674476 447393 674528 447399
rect 674476 447335 674528 447341
rect 674536 446744 674588 446750
rect 674536 446686 674588 446692
rect 674480 446620 674532 446626
rect 674480 446562 674532 446568
rect 674420 446391 674472 446397
rect 674420 446333 674472 446339
rect 674364 446197 674416 446203
rect 674364 446139 674416 446145
rect 674424 445548 674476 445554
rect 674424 445490 674476 445496
rect 674368 445424 674420 445430
rect 674368 445366 674420 445372
rect 674308 445195 674360 445201
rect 674308 445137 674360 445143
rect 674252 445001 674304 445007
rect 674252 444943 674304 444949
rect 674312 444352 674364 444358
rect 674312 444294 674364 444300
rect 674256 444228 674308 444234
rect 674256 444170 674308 444176
rect 674196 443999 674248 444005
rect 674196 443941 674248 443947
rect 674140 443805 674192 443811
rect 674140 443747 674192 443753
rect 674200 443156 674252 443162
rect 674200 443098 674252 443104
rect 674144 443032 674196 443038
rect 674144 442974 674196 442980
rect 674084 442803 674136 442809
rect 674084 442745 674136 442751
rect 674028 442609 674080 442615
rect 674028 442551 674080 442557
rect 674088 441960 674140 441966
rect 674088 441902 674140 441908
rect 674032 441836 674084 441842
rect 674032 441778 674084 441784
rect 673972 441607 674024 441613
rect 673972 441549 674024 441555
rect 673916 441413 673968 441419
rect 673916 441355 673968 441361
rect 673976 440764 674028 440770
rect 673976 440706 674028 440712
rect 673920 440640 673972 440646
rect 673920 440582 673972 440588
rect 673860 440411 673912 440417
rect 673860 440353 673912 440359
rect 673804 440217 673856 440223
rect 673804 440159 673856 440165
rect 673864 439568 673916 439574
rect 673864 439510 673916 439516
rect 673808 439444 673860 439450
rect 673808 439386 673860 439392
rect 43587 340370 43639 340376
rect 43587 340312 43639 340318
rect 43527 339721 43579 339727
rect 43527 339663 43579 339669
rect 43527 225372 43555 339663
rect 43583 339597 43635 339603
rect 43583 339539 43635 339545
rect 43583 225428 43611 339539
rect 43667 339374 43695 354730
rect 43643 339368 43695 339374
rect 43643 339310 43695 339316
rect 43723 339180 43751 354530
rect 43699 339174 43751 339180
rect 43699 339116 43751 339122
rect 43639 338525 43691 338531
rect 43639 338467 43691 338473
rect 43639 225484 43667 338467
rect 43695 338401 43747 338407
rect 43695 338343 43747 338349
rect 43695 225540 43723 338343
rect 43779 338178 43807 354330
rect 43755 338172 43807 338178
rect 43755 338114 43807 338120
rect 43835 337984 43863 354130
rect 43811 337978 43863 337984
rect 43811 337920 43863 337926
rect 43751 337329 43803 337335
rect 43751 337271 43803 337277
rect 43751 225596 43779 337271
rect 43807 337205 43859 337211
rect 43807 337147 43859 337153
rect 43807 225652 43835 337147
rect 43891 336958 43919 353930
rect 43867 336952 43919 336958
rect 43867 336894 43919 336900
rect 43947 336788 43975 353730
rect 43923 336782 43975 336788
rect 43923 336724 43975 336730
rect 43863 336133 43915 336139
rect 43863 336075 43915 336081
rect 43863 225708 43891 336075
rect 43919 336009 43971 336015
rect 43919 335951 43971 335957
rect 43919 225764 43947 335951
rect 44003 335786 44031 353530
rect 43979 335780 44031 335786
rect 43979 335722 44031 335728
rect 44059 335592 44087 353330
rect 44035 335586 44087 335592
rect 44035 335528 44087 335534
rect 43975 334937 44027 334943
rect 43975 334879 44027 334885
rect 43975 225820 44003 334879
rect 44031 334813 44083 334819
rect 44031 334755 44083 334761
rect 44031 225876 44059 334755
rect 394098 225904 394104 225928
rect 134098 225876 134104 225900
rect 44031 225848 134104 225876
rect 134156 225848 134162 225900
rect 134941 225852 134947 225904
rect 134999 225876 394104 225904
rect 394156 225876 394162 225928
rect 394941 225880 394947 225932
rect 394999 225904 673748 225932
rect 394999 225880 395005 225904
rect 134999 225852 135005 225876
rect 395170 225848 395176 225872
rect 135170 225820 135176 225844
rect 43975 225792 135176 225820
rect 135228 225792 135234 225844
rect 135943 225796 135949 225848
rect 136001 225820 395176 225848
rect 395228 225820 395234 225872
rect 395943 225824 395949 225876
rect 396001 225848 673692 225876
rect 396001 225824 396007 225848
rect 136001 225796 136007 225820
rect 395294 225792 395300 225816
rect 135294 225764 135300 225788
rect 43919 225736 135300 225764
rect 135352 225736 135358 225788
rect 136137 225740 136143 225792
rect 136195 225764 395300 225792
rect 395352 225764 395358 225816
rect 396137 225768 396143 225820
rect 396195 225792 673636 225820
rect 396195 225768 396201 225792
rect 136195 225740 136201 225764
rect 396366 225736 396372 225760
rect 136366 225708 136372 225732
rect 43863 225680 136372 225708
rect 136424 225680 136430 225732
rect 137139 225684 137145 225736
rect 137197 225708 396372 225736
rect 396424 225708 396430 225760
rect 397139 225712 397145 225764
rect 397197 225736 673580 225764
rect 397197 225712 397203 225736
rect 137197 225684 137203 225708
rect 396490 225680 396496 225704
rect 136490 225652 136496 225676
rect 43807 225624 136496 225652
rect 136548 225624 136554 225676
rect 137333 225628 137339 225680
rect 137391 225652 396496 225680
rect 396548 225652 396554 225704
rect 397333 225656 397339 225708
rect 397391 225680 673524 225708
rect 397391 225656 397397 225680
rect 137391 225628 137397 225652
rect 397562 225624 397568 225648
rect 137562 225596 137568 225620
rect 43751 225568 137568 225596
rect 137620 225568 137626 225620
rect 138335 225572 138341 225624
rect 138393 225596 397568 225624
rect 397620 225596 397626 225648
rect 398335 225600 398341 225652
rect 398393 225624 673468 225652
rect 398393 225600 398399 225624
rect 138393 225572 138399 225596
rect 397686 225568 397692 225592
rect 137686 225540 137692 225564
rect 43695 225512 137692 225540
rect 137744 225512 137750 225564
rect 138529 225516 138535 225568
rect 138587 225540 397692 225568
rect 397744 225540 397750 225592
rect 398529 225544 398535 225596
rect 398587 225568 673412 225596
rect 398587 225544 398593 225568
rect 138587 225516 138593 225540
rect 398758 225512 398764 225536
rect 138758 225484 138764 225508
rect 43639 225456 138764 225484
rect 138816 225456 138822 225508
rect 139531 225460 139537 225512
rect 139589 225484 398764 225512
rect 398816 225484 398822 225536
rect 399531 225488 399537 225540
rect 399589 225512 673356 225540
rect 399589 225488 399595 225512
rect 139589 225460 139595 225484
rect 398882 225456 398888 225480
rect 138882 225428 138888 225452
rect 43583 225400 138888 225428
rect 138940 225400 138946 225452
rect 139725 225404 139731 225456
rect 139783 225428 398888 225456
rect 398940 225428 398946 225480
rect 399725 225432 399731 225484
rect 399783 225456 673300 225484
rect 399783 225432 399789 225456
rect 139783 225404 139789 225428
rect 399954 225400 399960 225424
rect 139954 225372 139960 225396
rect 43527 225344 139960 225372
rect 140012 225344 140018 225396
rect 140727 225348 140733 225400
rect 140785 225372 399960 225400
rect 400012 225372 400018 225424
rect 400727 225376 400733 225428
rect 400785 225400 673244 225428
rect 400785 225376 400791 225400
rect 140785 225348 140791 225372
rect 400078 225344 400084 225368
rect 140078 225316 140084 225340
rect 43471 225288 140084 225316
rect 140136 225288 140142 225340
rect 140897 225292 140903 225344
rect 140955 225316 400084 225344
rect 400136 225316 400142 225368
rect 400897 225320 400903 225372
rect 400955 225344 673188 225372
rect 400955 225320 400961 225344
rect 140955 225292 140961 225316
rect 401150 225288 401156 225312
rect 141150 225260 141156 225284
rect 43415 225232 141156 225260
rect 141208 225232 141214 225284
rect 141923 225236 141929 225288
rect 141981 225260 401156 225288
rect 401208 225260 401214 225312
rect 401923 225264 401929 225316
rect 401981 225288 673132 225316
rect 401981 225264 401987 225288
rect 141981 225236 141987 225260
rect 401274 225232 401280 225256
rect 141274 225204 141280 225228
rect 43359 225176 141280 225204
rect 141332 225176 141338 225228
rect 142117 225180 142123 225232
rect 142175 225204 401280 225232
rect 401332 225204 401338 225256
rect 402117 225208 402123 225260
rect 402175 225232 673076 225260
rect 402175 225208 402181 225232
rect 142175 225180 142181 225204
rect 402346 225176 402352 225200
rect 142346 225148 142352 225172
rect 43303 225120 142352 225148
rect 142404 225120 142410 225172
rect 143119 225124 143125 225176
rect 143177 225148 402352 225176
rect 402404 225148 402410 225200
rect 403119 225152 403125 225204
rect 403177 225176 673020 225204
rect 403177 225152 403183 225176
rect 143177 225124 143183 225148
rect 402470 225120 402476 225144
rect 142470 225092 142476 225116
rect 43247 225064 142476 225092
rect 142528 225064 142534 225116
rect 143289 225068 143295 225120
rect 143347 225092 402476 225120
rect 402528 225092 402534 225144
rect 403289 225096 403295 225148
rect 403347 225120 672964 225148
rect 403347 225096 403353 225120
rect 143347 225068 143353 225092
rect 403542 225064 403548 225088
rect 143542 225036 143548 225060
rect 43191 225008 143548 225036
rect 143600 225008 143606 225060
rect 144315 225012 144321 225064
rect 144373 225036 403548 225064
rect 403600 225036 403606 225088
rect 404315 225040 404321 225092
rect 404373 225064 672908 225092
rect 404373 225040 404379 225064
rect 144373 225012 144379 225036
rect 403666 225008 403672 225032
rect 143666 224980 143672 225004
rect 43135 224952 143672 224980
rect 143724 224952 143730 225004
rect 144509 224956 144515 225008
rect 144567 224980 403672 225008
rect 403724 224980 403730 225032
rect 404509 224984 404515 225036
rect 404567 225008 672852 225036
rect 404567 224984 404573 225008
rect 144567 224956 144573 224980
rect 404738 224952 404744 224976
rect 144738 224924 144744 224948
rect 43079 224896 144744 224924
rect 144796 224896 144802 224948
rect 145511 224900 145517 224952
rect 145569 224924 404744 224952
rect 404796 224924 404802 224976
rect 405511 224928 405517 224980
rect 405569 224952 672796 224980
rect 405569 224928 405575 224952
rect 145569 224900 145575 224924
rect 404862 224896 404868 224920
rect 144862 224868 144868 224892
rect 43023 224840 144868 224868
rect 144920 224840 144926 224892
rect 145705 224844 145711 224896
rect 145763 224868 404868 224896
rect 404920 224868 404926 224920
rect 405705 224872 405711 224924
rect 405763 224896 672740 224924
rect 405763 224872 405769 224896
rect 145763 224844 145769 224868
rect 405934 224840 405940 224864
rect 145934 224812 145940 224836
rect 42967 224784 145940 224812
rect 145992 224784 145998 224836
rect 146707 224788 146713 224840
rect 146765 224812 405940 224840
rect 405992 224812 405998 224864
rect 406707 224816 406713 224868
rect 406765 224840 672684 224868
rect 406765 224816 406771 224840
rect 146765 224788 146771 224812
rect 406058 224784 406064 224808
rect 146058 224756 146064 224780
rect 42911 224728 146064 224756
rect 146116 224728 146122 224780
rect 146901 224732 146907 224784
rect 146959 224756 406064 224784
rect 406116 224756 406122 224808
rect 406901 224760 406907 224812
rect 406959 224784 672628 224812
rect 406959 224760 406965 224784
rect 146959 224732 146965 224756
rect 407130 224728 407136 224752
rect 147130 224700 147136 224724
rect 42855 224672 147136 224700
rect 147188 224672 147194 224724
rect 147903 224676 147909 224728
rect 147961 224700 407136 224728
rect 407188 224700 407194 224752
rect 407903 224704 407909 224756
rect 407961 224728 672572 224756
rect 407961 224704 407967 224728
rect 147961 224676 147967 224700
rect 407254 224672 407260 224696
rect 147254 224644 147260 224668
rect 42799 224616 147260 224644
rect 147312 224616 147318 224668
rect 148097 224620 148103 224672
rect 148155 224644 407260 224672
rect 407312 224644 407318 224696
rect 408097 224648 408103 224700
rect 408155 224672 672516 224700
rect 408155 224648 408161 224672
rect 148155 224620 148161 224644
rect 408326 224616 408332 224640
rect 148326 224588 148332 224612
rect 42743 224560 148332 224588
rect 148384 224560 148390 224612
rect 149099 224564 149105 224616
rect 149157 224588 408332 224616
rect 408384 224588 408390 224640
rect 409099 224592 409105 224644
rect 409157 224616 672460 224644
rect 409157 224592 409163 224616
rect 149157 224564 149163 224588
rect 408450 224560 408456 224584
rect 148450 224532 148456 224556
rect 42687 224504 148456 224532
rect 148508 224504 148514 224556
rect 149293 224508 149299 224560
rect 149351 224532 408456 224560
rect 408508 224532 408514 224584
rect 409293 224536 409299 224588
rect 409351 224560 672404 224588
rect 409351 224536 409357 224560
rect 149351 224508 149357 224532
rect 409522 224504 409528 224528
rect 149522 224476 149528 224500
rect 42631 224448 149528 224476
rect 149580 224448 149586 224500
rect 150295 224452 150301 224504
rect 150353 224476 409528 224504
rect 409580 224476 409586 224528
rect 410295 224480 410301 224532
rect 410353 224504 672348 224532
rect 410353 224480 410359 224504
rect 150353 224452 150359 224476
rect 409646 224448 409652 224472
rect 149646 224420 149652 224444
rect 42575 224392 149652 224420
rect 149704 224392 149710 224444
rect 150489 224396 150495 224448
rect 150547 224420 409652 224448
rect 409704 224420 409710 224472
rect 410489 224424 410495 224476
rect 410547 224448 672292 224476
rect 410547 224424 410553 224448
rect 150547 224396 150553 224420
rect 410718 224392 410724 224416
rect 150718 224364 150724 224388
rect 42519 224336 150724 224364
rect 150776 224336 150782 224388
rect 151491 224340 151497 224392
rect 151549 224364 410724 224392
rect 410776 224364 410782 224416
rect 411491 224368 411497 224420
rect 411549 224392 672236 224420
rect 411549 224368 411555 224392
rect 151549 224340 151555 224364
rect 410842 224336 410848 224360
rect 150842 224308 150848 224332
rect 42463 224280 150848 224308
rect 150900 224280 150906 224332
rect 151685 224284 151691 224336
rect 151743 224308 410848 224336
rect 410900 224308 410906 224360
rect 411685 224312 411691 224364
rect 411743 224336 672180 224364
rect 411743 224312 411749 224336
rect 151743 224284 151749 224308
rect 411914 224280 411920 224304
rect 151914 224252 151920 224276
rect 42407 224224 151920 224252
rect 151972 224224 151978 224276
rect 152687 224228 152693 224280
rect 152745 224252 411920 224280
rect 411972 224252 411978 224304
rect 412687 224256 412693 224308
rect 412745 224280 672124 224308
rect 412745 224256 412751 224280
rect 152745 224228 152751 224252
rect 412038 224224 412044 224248
rect 152038 224196 152044 224220
rect 131123 224168 152044 224196
rect 152096 224168 152102 224220
rect 152881 224172 152887 224224
rect 152939 224196 412044 224224
rect 412096 224196 412102 224248
rect 412881 224200 412887 224252
rect 412939 224224 672068 224252
rect 412939 224200 412945 224224
rect 152939 224172 152945 224196
rect 413110 224168 413116 224192
rect 153110 224140 153116 224164
rect 131323 224112 153116 224140
rect 153168 224112 153174 224164
rect 153883 224116 153889 224168
rect 153941 224140 413116 224168
rect 413168 224140 413174 224192
rect 413883 224144 413889 224196
rect 413941 224168 672012 224196
rect 413941 224144 413947 224168
rect 153941 224116 153947 224140
rect 413234 224112 413240 224136
rect 153234 224084 153240 224108
rect 131523 224056 153240 224084
rect 153292 224056 153298 224108
rect 154077 224060 154083 224112
rect 154135 224084 413240 224112
rect 413292 224084 413298 224136
rect 414077 224088 414083 224140
rect 414135 224112 671956 224140
rect 414135 224088 414141 224112
rect 154135 224060 154141 224084
rect 414306 224056 414312 224080
rect 154306 224028 154312 224052
rect 131723 224000 154312 224028
rect 154364 224000 154370 224052
rect 155079 224004 155085 224056
rect 155137 224028 414312 224056
rect 414364 224028 414370 224080
rect 415079 224032 415085 224084
rect 415137 224056 671900 224084
rect 415137 224032 415143 224056
rect 155137 224004 155143 224028
rect 414430 224000 414436 224024
rect 154430 223972 154436 223996
rect 131923 223944 154436 223972
rect 154488 223944 154494 223996
rect 155249 223948 155255 224000
rect 155307 223972 414436 224000
rect 414488 223972 414494 224024
rect 415249 223976 415255 224028
rect 415307 224000 671844 224028
rect 415307 223976 415313 224000
rect 155307 223948 155313 223972
rect 415502 223944 415508 223968
rect 155502 223916 155508 223940
rect 132123 223888 155508 223916
rect 155560 223888 155566 223940
rect 156275 223892 156281 223944
rect 156333 223916 415508 223944
rect 415560 223916 415566 223968
rect 416275 223920 416281 223972
rect 416333 223944 671788 223972
rect 416333 223920 416339 223944
rect 156333 223892 156339 223916
rect 415626 223888 415632 223912
rect 155626 223860 155632 223884
rect 132323 223832 155632 223860
rect 155684 223832 155690 223884
rect 156469 223836 156475 223888
rect 156527 223860 415632 223888
rect 415684 223860 415690 223912
rect 416469 223864 416475 223916
rect 416527 223888 671732 223916
rect 416527 223864 416533 223888
rect 156527 223836 156533 223860
rect 416698 223832 416704 223856
rect 156698 223804 156704 223828
rect 132523 223776 156704 223804
rect 156756 223776 156762 223828
rect 157471 223780 157477 223832
rect 157529 223804 416704 223832
rect 416756 223804 416762 223856
rect 417471 223808 417477 223860
rect 417529 223832 671676 223860
rect 417529 223808 417535 223832
rect 157529 223780 157535 223804
rect 416822 223776 416828 223800
rect 156822 223748 156828 223772
rect 132723 223720 156828 223748
rect 156880 223720 156886 223772
rect 157641 223724 157647 223776
rect 157699 223748 416828 223776
rect 416880 223748 416886 223800
rect 417641 223752 417647 223804
rect 417699 223776 671620 223804
rect 417699 223752 417705 223776
rect 157699 223724 157705 223748
rect 417894 223720 417900 223744
rect 157894 223692 157900 223716
rect 132923 223664 157900 223692
rect 157952 223664 157958 223716
rect 158667 223668 158673 223720
rect 158725 223692 417900 223720
rect 417952 223692 417958 223744
rect 418667 223696 418673 223748
rect 418725 223720 671564 223748
rect 418725 223696 418731 223720
rect 158725 223668 158731 223692
rect 418018 223664 418024 223688
rect 158018 223636 158024 223660
rect 133123 223608 158024 223636
rect 158076 223608 158082 223660
rect 158861 223612 158867 223664
rect 158919 223636 418024 223664
rect 418076 223636 418082 223688
rect 418861 223640 418867 223692
rect 418919 223664 671508 223692
rect 418919 223640 418925 223664
rect 158919 223612 158925 223636
rect 134094 223272 134146 223284
rect 135290 223272 135342 223284
rect 134836 223162 134848 223214
rect 135066 223162 135078 223214
rect 134094 223090 134146 223102
rect 136486 223272 136538 223284
rect 136032 223162 136044 223214
rect 136262 223162 136274 223214
rect 135290 223090 135342 223102
rect 137682 223272 137734 223284
rect 137228 223162 137240 223214
rect 137458 223162 137470 223214
rect 136486 223090 136538 223102
rect 138878 223272 138930 223284
rect 138424 223162 138436 223214
rect 138654 223162 138666 223214
rect 137682 223090 137734 223102
rect 140074 223272 140126 223284
rect 139620 223162 139632 223214
rect 139850 223162 139862 223214
rect 138878 223090 138930 223102
rect 141270 223272 141322 223284
rect 140816 223162 140828 223214
rect 141046 223162 141058 223214
rect 140074 223090 140126 223102
rect 142466 223272 142518 223284
rect 142012 223162 142024 223214
rect 142242 223162 142254 223214
rect 141270 223090 141322 223102
rect 143662 223272 143714 223284
rect 143208 223162 143220 223214
rect 143438 223162 143450 223214
rect 142466 223090 142518 223102
rect 144858 223272 144910 223284
rect 144404 223162 144416 223214
rect 144634 223162 144646 223214
rect 143662 223090 143714 223102
rect 146054 223272 146106 223284
rect 145600 223162 145612 223214
rect 145830 223162 145842 223214
rect 144858 223090 144910 223102
rect 147250 223272 147302 223284
rect 146796 223162 146808 223214
rect 147026 223162 147038 223214
rect 146054 223090 146106 223102
rect 148446 223272 148498 223284
rect 147992 223162 148004 223214
rect 148222 223162 148234 223214
rect 147250 223090 147302 223102
rect 149642 223272 149694 223284
rect 149188 223162 149200 223214
rect 149418 223162 149430 223214
rect 148446 223090 148498 223102
rect 150838 223272 150890 223284
rect 150384 223162 150396 223214
rect 150614 223162 150626 223214
rect 149642 223090 149694 223102
rect 152034 223272 152086 223284
rect 151580 223162 151592 223214
rect 151810 223162 151822 223214
rect 150838 223090 150890 223102
rect 153230 223272 153282 223284
rect 152776 223162 152788 223214
rect 153006 223162 153018 223214
rect 152034 223090 152086 223102
rect 154426 223272 154478 223284
rect 153972 223162 153984 223214
rect 154202 223162 154214 223214
rect 153230 223090 153282 223102
rect 155622 223272 155674 223284
rect 155168 223162 155180 223214
rect 155398 223162 155410 223214
rect 154426 223090 154478 223102
rect 156818 223272 156870 223284
rect 156364 223162 156376 223214
rect 156594 223162 156606 223214
rect 155622 223090 155674 223102
rect 158014 223272 158066 223284
rect 157560 223162 157572 223214
rect 157790 223162 157802 223214
rect 156818 223090 156870 223102
rect 394094 223272 394146 223284
rect 158756 223162 158768 223214
rect 158986 223162 158998 223214
rect 158014 223090 158066 223102
rect 395290 223272 395342 223284
rect 394836 223162 394848 223214
rect 395066 223162 395078 223214
rect 394094 223090 394146 223102
rect 396486 223272 396538 223284
rect 396032 223162 396044 223214
rect 396262 223162 396274 223214
rect 395290 223090 395342 223102
rect 397682 223272 397734 223284
rect 397228 223162 397240 223214
rect 397458 223162 397470 223214
rect 396486 223090 396538 223102
rect 398878 223272 398930 223284
rect 398424 223162 398436 223214
rect 398654 223162 398666 223214
rect 397682 223090 397734 223102
rect 400074 223272 400126 223284
rect 399620 223162 399632 223214
rect 399850 223162 399862 223214
rect 398878 223090 398930 223102
rect 401270 223272 401322 223284
rect 400816 223162 400828 223214
rect 401046 223162 401058 223214
rect 400074 223090 400126 223102
rect 402466 223272 402518 223284
rect 402012 223162 402024 223214
rect 402242 223162 402254 223214
rect 401270 223090 401322 223102
rect 403662 223272 403714 223284
rect 403208 223162 403220 223214
rect 403438 223162 403450 223214
rect 402466 223090 402518 223102
rect 404858 223272 404910 223284
rect 404404 223162 404416 223214
rect 404634 223162 404646 223214
rect 403662 223090 403714 223102
rect 406054 223272 406106 223284
rect 405600 223162 405612 223214
rect 405830 223162 405842 223214
rect 404858 223090 404910 223102
rect 407250 223272 407302 223284
rect 406796 223162 406808 223214
rect 407026 223162 407038 223214
rect 406054 223090 406106 223102
rect 408446 223272 408498 223284
rect 407992 223162 408004 223214
rect 408222 223162 408234 223214
rect 407250 223090 407302 223102
rect 409642 223272 409694 223284
rect 409188 223162 409200 223214
rect 409418 223162 409430 223214
rect 408446 223090 408498 223102
rect 410838 223272 410890 223284
rect 410384 223162 410396 223214
rect 410614 223162 410626 223214
rect 409642 223090 409694 223102
rect 412034 223272 412086 223284
rect 411580 223162 411592 223214
rect 411810 223162 411822 223214
rect 410838 223090 410890 223102
rect 413230 223272 413282 223284
rect 412776 223162 412788 223214
rect 413006 223162 413018 223214
rect 412034 223090 412086 223102
rect 414426 223272 414478 223284
rect 413972 223162 413984 223214
rect 414202 223162 414214 223214
rect 413230 223090 413282 223102
rect 415622 223272 415674 223284
rect 415168 223162 415180 223214
rect 415398 223162 415410 223214
rect 414426 223090 414478 223102
rect 416818 223272 416870 223284
rect 416364 223162 416376 223214
rect 416594 223162 416606 223214
rect 415622 223090 415674 223102
rect 418014 223272 418066 223284
rect 417560 223162 417572 223214
rect 417790 223162 417802 223214
rect 416818 223090 416870 223102
rect 418756 223162 418768 223214
rect 418986 223162 418998 223214
rect 418014 223090 418066 223102
rect 671480 223050 671508 223664
rect 671536 222850 671564 223720
rect 135936 222660 135988 222672
rect 135106 222550 135118 222602
rect 135336 222550 135348 222602
rect 137132 222660 137184 222672
rect 136302 222550 136314 222602
rect 136532 222550 136544 222602
rect 135936 222478 135988 222490
rect 138328 222660 138380 222672
rect 137498 222550 137510 222602
rect 137728 222550 137740 222602
rect 137132 222478 137184 222490
rect 139524 222660 139576 222672
rect 138694 222550 138706 222602
rect 138924 222550 138936 222602
rect 138328 222478 138380 222490
rect 140720 222660 140772 222672
rect 139890 222550 139902 222602
rect 140120 222550 140132 222602
rect 139524 222478 139576 222490
rect 141916 222660 141968 222672
rect 141086 222550 141098 222602
rect 141316 222550 141328 222602
rect 140720 222478 140772 222490
rect 143112 222660 143164 222672
rect 142282 222550 142294 222602
rect 142512 222550 142524 222602
rect 141916 222478 141968 222490
rect 144308 222660 144360 222672
rect 143478 222550 143490 222602
rect 143708 222550 143720 222602
rect 143112 222478 143164 222490
rect 145504 222660 145556 222672
rect 144674 222550 144686 222602
rect 144904 222550 144916 222602
rect 144308 222478 144360 222490
rect 146700 222660 146752 222672
rect 145870 222550 145882 222602
rect 146100 222550 146112 222602
rect 145504 222478 145556 222490
rect 147896 222660 147948 222672
rect 147066 222550 147078 222602
rect 147296 222550 147308 222602
rect 146700 222478 146752 222490
rect 149092 222660 149144 222672
rect 148262 222550 148274 222602
rect 148492 222550 148504 222602
rect 147896 222478 147948 222490
rect 150288 222660 150340 222672
rect 149458 222550 149470 222602
rect 149688 222550 149700 222602
rect 149092 222478 149144 222490
rect 151484 222660 151536 222672
rect 150654 222550 150666 222602
rect 150884 222550 150896 222602
rect 150288 222478 150340 222490
rect 152680 222660 152732 222672
rect 151850 222550 151862 222602
rect 152080 222550 152092 222602
rect 151484 222478 151536 222490
rect 153876 222660 153928 222672
rect 153046 222550 153058 222602
rect 153276 222550 153288 222602
rect 152680 222478 152732 222490
rect 155072 222660 155124 222672
rect 154242 222550 154254 222602
rect 154472 222550 154484 222602
rect 153876 222478 153928 222490
rect 156268 222660 156320 222672
rect 155438 222550 155450 222602
rect 155668 222550 155680 222602
rect 155072 222478 155124 222490
rect 157464 222660 157516 222672
rect 156634 222550 156646 222602
rect 156864 222550 156876 222602
rect 156268 222478 156320 222490
rect 157464 222478 157516 222490
rect 158016 222660 158068 222672
rect 395936 222660 395988 222672
rect 158656 222550 158668 222602
rect 158886 222550 158898 222602
rect 395106 222550 395118 222602
rect 395336 222550 395348 222602
rect 158016 222478 158068 222490
rect 397132 222660 397184 222672
rect 396302 222550 396314 222602
rect 396532 222550 396544 222602
rect 395936 222478 395988 222490
rect 398328 222660 398380 222672
rect 397498 222550 397510 222602
rect 397728 222550 397740 222602
rect 397132 222478 397184 222490
rect 399524 222660 399576 222672
rect 398694 222550 398706 222602
rect 398924 222550 398936 222602
rect 398328 222478 398380 222490
rect 400720 222660 400772 222672
rect 399890 222550 399902 222602
rect 400120 222550 400132 222602
rect 399524 222478 399576 222490
rect 401916 222660 401968 222672
rect 401086 222550 401098 222602
rect 401316 222550 401328 222602
rect 400720 222478 400772 222490
rect 403112 222660 403164 222672
rect 402282 222550 402294 222602
rect 402512 222550 402524 222602
rect 401916 222478 401968 222490
rect 404308 222660 404360 222672
rect 403478 222550 403490 222602
rect 403708 222550 403720 222602
rect 403112 222478 403164 222490
rect 405504 222660 405556 222672
rect 404674 222550 404686 222602
rect 404904 222550 404916 222602
rect 404308 222478 404360 222490
rect 406700 222660 406752 222672
rect 405870 222550 405882 222602
rect 406100 222550 406112 222602
rect 405504 222478 405556 222490
rect 407896 222660 407948 222672
rect 407066 222550 407078 222602
rect 407296 222550 407308 222602
rect 406700 222478 406752 222490
rect 409092 222660 409144 222672
rect 408262 222550 408274 222602
rect 408492 222550 408504 222602
rect 407896 222478 407948 222490
rect 410288 222660 410340 222672
rect 409458 222550 409470 222602
rect 409688 222550 409700 222602
rect 409092 222478 409144 222490
rect 411484 222660 411536 222672
rect 410654 222550 410666 222602
rect 410884 222550 410896 222602
rect 410288 222478 410340 222490
rect 412680 222660 412732 222672
rect 411850 222550 411862 222602
rect 412080 222550 412092 222602
rect 411484 222478 411536 222490
rect 413876 222660 413928 222672
rect 413046 222550 413058 222602
rect 413276 222550 413288 222602
rect 412680 222478 412732 222490
rect 415072 222660 415124 222672
rect 414242 222550 414254 222602
rect 414472 222550 414484 222602
rect 413876 222478 413928 222490
rect 416268 222660 416320 222672
rect 415438 222550 415450 222602
rect 415668 222550 415680 222602
rect 415072 222478 415124 222490
rect 417464 222660 417516 222672
rect 416634 222550 416646 222602
rect 416864 222550 416876 222602
rect 416268 222478 416320 222490
rect 417464 222478 417516 222490
rect 418016 222660 418068 222672
rect 671592 222650 671620 223776
rect 418656 222550 418668 222602
rect 418886 222550 418898 222602
rect 418016 222478 418068 222490
rect 671648 222450 671676 223832
rect 671704 222250 671732 223888
rect 671760 222050 671788 223944
rect 671816 221850 671844 224000
rect 671872 221650 671900 224056
rect 671928 221450 671956 224112
rect 671984 221250 672012 224168
rect 672040 221050 672068 224224
rect 672096 220850 672124 224280
rect 672152 220650 672180 224336
rect 672208 220450 672236 224392
rect 672264 220250 672292 224448
rect 672320 220050 672348 224504
rect 672376 219850 672404 224560
rect 672432 219650 672460 224616
rect 672488 219450 672516 224672
rect 672544 219250 672572 224728
rect 672600 219050 672628 224784
rect 672656 218850 672684 224840
rect 672712 218650 672740 224896
rect 672768 218450 672796 224952
rect 672824 218250 672852 225008
rect 672880 218050 672908 225064
rect 672936 217850 672964 225120
rect 672992 217650 673020 225176
rect 673048 217450 673076 225232
rect 673104 217250 673132 225288
rect 673160 217050 673188 225344
rect 673216 216850 673244 225400
rect 673272 216650 673300 225456
rect 673328 216450 673356 225512
rect 673384 216250 673412 225568
rect 673440 216050 673468 225624
rect 673496 215850 673524 225680
rect 673552 215650 673580 225736
rect 673608 215450 673636 225792
rect 673664 215250 673692 225848
rect 673720 215050 673748 225904
rect 673832 215050 673860 439386
rect 673888 214850 673916 439510
rect 673944 214650 673972 440582
rect 674000 214450 674028 440706
rect 674056 214250 674084 441778
rect 674112 214050 674140 441902
rect 674168 213850 674196 442974
rect 674224 213650 674252 443098
rect 674280 213450 674308 444170
rect 674336 213250 674364 444294
rect 674392 213050 674420 445366
rect 674448 212850 674476 445490
rect 674504 212650 674532 446562
rect 674560 212450 674588 446686
rect 674616 212250 674644 447758
rect 674672 212050 674700 447882
rect 674728 211850 674756 448954
rect 674784 211650 674812 449078
rect 674840 211450 674868 450150
rect 674896 211250 674924 450274
rect 674952 211050 674980 451346
rect 675008 210850 675036 451470
rect 675064 210650 675092 452542
rect 675120 210450 675148 452666
rect 676858 452662 676870 452714
rect 677040 452662 677052 452714
rect 677540 452708 677592 452720
rect 677540 452478 677592 452490
rect 676928 452438 676980 452450
rect 676928 452208 676980 452220
rect 677470 452112 677482 452164
rect 677652 452112 677664 452164
rect 676858 451466 676870 451518
rect 677040 451466 677052 451518
rect 677540 451512 677592 451524
rect 677540 451282 677592 451294
rect 676928 451242 676980 451254
rect 676928 451012 676980 451024
rect 677470 450916 677482 450968
rect 677652 450916 677664 450968
rect 676858 450270 676870 450322
rect 677040 450270 677052 450322
rect 677540 450316 677592 450328
rect 677540 450086 677592 450098
rect 676928 450046 676980 450058
rect 676928 449816 676980 449828
rect 677470 449720 677482 449772
rect 677652 449720 677664 449772
rect 676858 449074 676870 449126
rect 677040 449074 677052 449126
rect 677540 449120 677592 449132
rect 677540 448890 677592 448902
rect 676928 448850 676980 448862
rect 676928 448620 676980 448632
rect 677470 448524 677482 448576
rect 677652 448524 677664 448576
rect 676858 447878 676870 447930
rect 677040 447878 677052 447930
rect 677540 447924 677592 447936
rect 677540 447694 677592 447706
rect 676928 447654 676980 447666
rect 676928 447424 676980 447436
rect 677470 447328 677482 447380
rect 677652 447328 677664 447380
rect 676858 446682 676870 446734
rect 677040 446682 677052 446734
rect 677540 446728 677592 446740
rect 677540 446498 677592 446510
rect 676928 446458 676980 446470
rect 676928 446228 676980 446240
rect 677470 446132 677482 446184
rect 677652 446132 677664 446184
rect 676858 445486 676870 445538
rect 677040 445486 677052 445538
rect 677540 445532 677592 445544
rect 677540 445302 677592 445314
rect 676928 445262 676980 445274
rect 676928 445032 676980 445044
rect 677470 444936 677482 444988
rect 677652 444936 677664 444988
rect 676858 444290 676870 444342
rect 677040 444290 677052 444342
rect 677540 444336 677592 444348
rect 677540 444106 677592 444118
rect 676928 444066 676980 444078
rect 676928 443836 676980 443848
rect 677470 443740 677482 443792
rect 677652 443740 677664 443792
rect 676858 443094 676870 443146
rect 677040 443094 677052 443146
rect 677540 443140 677592 443152
rect 677540 442910 677592 442922
rect 676928 442870 676980 442882
rect 676928 442640 676980 442652
rect 677470 442544 677482 442596
rect 677652 442544 677664 442596
rect 676858 441898 676870 441950
rect 677040 441898 677052 441950
rect 677540 441944 677592 441956
rect 677540 441714 677592 441726
rect 676928 441674 676980 441686
rect 676928 441444 676980 441456
rect 677470 441348 677482 441400
rect 677652 441348 677664 441400
rect 676858 440702 676870 440754
rect 677040 440702 677052 440754
rect 677540 440748 677592 440760
rect 677540 440518 677592 440530
rect 676928 440478 676980 440490
rect 676928 440248 676980 440260
rect 677470 440152 677482 440204
rect 677652 440152 677664 440204
rect 676858 439506 676870 439558
rect 677040 439506 677052 439558
rect 677540 439552 677592 439564
rect 677540 439322 677592 439334
<< via1 >>
rect 417027 997507 417384 997567
rect 664237 997425 664594 997485
rect 168590 997178 168947 997238
rect 416862 997217 416870 997387
rect 416870 997217 416904 997387
rect 416904 997217 416914 997387
rect 417514 997319 417732 997327
rect 417514 997285 417732 997319
rect 417514 997275 417732 997285
rect 662863 997135 662871 997305
rect 662871 997135 662905 997305
rect 662905 997135 662915 997305
rect 663515 997237 663733 997245
rect 663515 997203 663733 997237
rect 663515 997193 663733 997203
rect 664059 997135 664067 997305
rect 664067 997135 664101 997305
rect 664101 997135 664111 997305
rect 664711 997237 664929 997245
rect 664711 997203 664929 997237
rect 664711 997193 664929 997203
rect 665255 997135 665263 997305
rect 665263 997135 665297 997305
rect 665297 997135 665307 997305
rect 665907 997237 666125 997245
rect 665907 997203 666125 997237
rect 665907 997193 666125 997203
rect 666451 997135 666459 997305
rect 666459 997135 666493 997305
rect 666493 997135 666503 997305
rect 667103 997237 667321 997245
rect 667103 997203 667321 997237
rect 667103 997193 667321 997203
rect 167052 996994 167270 997002
rect 167052 996960 167270 996994
rect 167052 996950 167270 996960
rect 167870 996892 167880 997062
rect 167880 996892 167914 997062
rect 167914 996892 167922 997062
rect 168248 996994 168466 997002
rect 168248 996960 168466 996994
rect 168248 996950 168466 996960
rect 169066 996892 169076 997062
rect 169076 996892 169110 997062
rect 169110 996892 169118 997062
rect 169444 996994 169662 997002
rect 169444 996960 169662 996994
rect 169444 996950 169662 996960
rect 170262 996892 170272 997062
rect 170272 996892 170306 997062
rect 170306 996892 170314 997062
rect 418223 996966 418580 997026
rect 665433 996884 665790 996944
rect 169786 996637 170143 996697
rect 416588 996707 416806 996715
rect 416588 996673 416806 996707
rect 416588 996663 416806 996673
rect 417508 996605 417516 996775
rect 417516 996605 417550 996775
rect 417550 996605 417560 996775
rect 662589 996625 662807 996633
rect 662589 996591 662807 996625
rect 662589 996581 662807 996591
rect 663509 996523 663517 996693
rect 663517 996523 663551 996693
rect 663551 996523 663561 996693
rect 663785 996625 664003 996633
rect 663785 996591 664003 996625
rect 663785 996581 664003 996591
rect 664705 996523 664713 996693
rect 664713 996523 664747 996693
rect 664747 996523 664757 996693
rect 664981 996625 665199 996633
rect 664981 996591 665199 996625
rect 664981 996581 665199 996591
rect 665901 996523 665909 996693
rect 665909 996523 665943 996693
rect 665943 996523 665953 996693
rect 666177 996625 666395 996633
rect 666177 996591 666395 996625
rect 666177 996581 666395 996591
rect 667097 996523 667105 996693
rect 667105 996523 667139 996693
rect 667139 996523 667149 996693
rect 167224 996280 167234 996450
rect 167234 996280 167268 996450
rect 167268 996280 167276 996450
rect 167978 996382 168196 996390
rect 167978 996348 168196 996382
rect 167978 996338 168196 996348
rect 168420 996280 168430 996450
rect 168430 996280 168464 996450
rect 168464 996280 168472 996450
rect 169174 996382 169392 996390
rect 169174 996348 169392 996382
rect 169174 996338 169392 996348
rect 169616 996280 169626 996450
rect 169626 996280 169660 996450
rect 169660 996280 169668 996450
rect 417027 996425 417384 996485
rect 170370 996382 170588 996390
rect 170370 996348 170588 996382
rect 170370 996338 170588 996348
rect 664237 996343 664594 996403
rect 168590 996096 168947 996156
rect 40554 891200 40562 891418
rect 40562 891200 40596 891418
rect 40596 891200 40606 891418
rect 169626 995405 169678 995457
rect 170469 995401 170521 995453
rect 42467 891299 42519 891351
rect 169502 995349 169554 995401
rect 170275 995345 170327 995397
rect 39882 891136 40052 891144
rect 39882 891102 40052 891136
rect 39882 891092 40052 891102
rect 42523 891105 42575 891157
rect 39942 890274 39950 890492
rect 39950 890274 39984 890492
rect 39984 890274 39994 890492
rect 40494 890490 40664 890498
rect 40494 890456 40664 890490
rect 40494 890446 40664 890456
rect 42463 890456 42515 890508
rect 40554 890004 40562 890222
rect 40562 890004 40596 890222
rect 40596 890004 40606 890222
rect 39882 889940 40052 889948
rect 39882 889906 40052 889940
rect 39882 889896 40052 889906
rect 40241 889384 40301 889741
rect 39942 889078 39950 889296
rect 39950 889078 39984 889296
rect 39984 889078 39994 889296
rect 40494 889294 40664 889302
rect 40494 889260 40664 889294
rect 40494 889250 40664 889260
rect 40554 888808 40562 889026
rect 40562 888808 40596 889026
rect 40596 888808 40606 889026
rect 39882 888744 40052 888752
rect 39882 888710 40052 888744
rect 39882 888700 40052 888710
rect 39700 888188 39760 888545
rect 40782 888188 40842 888545
rect 39942 887882 39950 888100
rect 39950 887882 39984 888100
rect 39984 887882 39994 888100
rect 40494 888098 40664 888106
rect 40494 888064 40664 888098
rect 40494 888054 40664 888064
rect 40554 887612 40562 887830
rect 40562 887612 40596 887830
rect 40596 887612 40606 887830
rect 39882 887548 40052 887556
rect 39882 887514 40052 887548
rect 39882 887504 40052 887514
rect 39942 886686 39950 886904
rect 39950 886686 39984 886904
rect 39984 886686 39994 886904
rect 40494 886902 40664 886910
rect 40494 886868 40664 886902
rect 40494 886858 40664 886868
rect 40554 886416 40562 886634
rect 40562 886416 40596 886634
rect 40596 886416 40606 886634
rect 39882 886352 40052 886360
rect 39882 886318 40052 886352
rect 39882 886308 40052 886318
rect 39942 885490 39950 885708
rect 39950 885490 39984 885708
rect 39984 885490 39994 885708
rect 40494 885706 40664 885714
rect 40494 885672 40664 885706
rect 40494 885662 40664 885672
rect 40579 610554 40587 610772
rect 40587 610554 40621 610772
rect 40621 610554 40631 610772
rect 42439 610653 42491 610705
rect 42519 890332 42571 890384
rect 168430 995293 168482 995345
rect 169249 995289 169301 995341
rect 42579 890079 42631 890131
rect 168306 995237 168358 995289
rect 169079 995233 169131 995285
rect 42635 889909 42687 889961
rect 39907 610490 40077 610498
rect 39907 610456 40077 610490
rect 39907 610446 40077 610456
rect 42495 610459 42547 610511
rect 42575 889260 42627 889312
rect 39967 609628 39975 609846
rect 39975 609628 40009 609846
rect 40009 609628 40019 609846
rect 40519 609844 40689 609852
rect 40519 609810 40689 609844
rect 40519 609800 40689 609810
rect 42435 609810 42487 609862
rect 40579 609358 40587 609576
rect 40587 609358 40621 609576
rect 40621 609358 40631 609576
rect 39907 609294 40077 609302
rect 39907 609260 40077 609294
rect 39907 609250 40077 609260
rect 39967 608432 39975 608650
rect 39975 608432 40009 608650
rect 40009 608432 40019 608650
rect 40519 608648 40689 608656
rect 40519 608614 40689 608648
rect 40519 608604 40689 608614
rect 40579 608162 40587 608380
rect 40587 608162 40621 608380
rect 40621 608162 40631 608380
rect 39907 608098 40077 608106
rect 39907 608064 40077 608098
rect 39907 608054 40077 608064
rect 39967 607236 39975 607454
rect 39975 607236 40009 607454
rect 40009 607236 40019 607454
rect 40519 607452 40689 607460
rect 40519 607418 40689 607452
rect 40519 607408 40689 607418
rect 40579 606966 40587 607184
rect 40587 606966 40621 607184
rect 40621 606966 40631 607184
rect 39907 606902 40077 606910
rect 39907 606868 40077 606902
rect 39907 606858 40077 606868
rect 39967 606040 39975 606258
rect 39975 606040 40009 606258
rect 40009 606040 40019 606258
rect 40519 606256 40689 606264
rect 40519 606222 40689 606256
rect 40519 606212 40689 606222
rect 40579 605770 40587 605988
rect 40587 605770 40621 605988
rect 40621 605770 40631 605988
rect 39907 605706 40077 605714
rect 39907 605672 40077 605706
rect 39907 605662 40077 605672
rect 40272 605210 40332 605567
rect 39967 604844 39975 605062
rect 39975 604844 40009 605062
rect 40009 604844 40019 605062
rect 40519 605060 40689 605068
rect 40519 605026 40689 605060
rect 40519 605016 40689 605026
rect 40579 604574 40587 604792
rect 40587 604574 40621 604792
rect 40621 604574 40631 604792
rect 39907 604510 40077 604518
rect 39907 604476 40077 604510
rect 39907 604466 40077 604476
rect 39731 604014 39791 604371
rect 40813 604014 40873 604371
rect 39967 603648 39975 603866
rect 39975 603648 40009 603866
rect 40009 603648 40019 603866
rect 40519 603864 40689 603872
rect 40519 603830 40689 603864
rect 40519 603820 40689 603830
rect 40579 603378 40587 603596
rect 40587 603378 40621 603596
rect 40621 603378 40631 603596
rect 39907 603314 40077 603322
rect 39907 603280 40077 603314
rect 39907 603270 40077 603280
rect 39967 602452 39975 602670
rect 39975 602452 40009 602670
rect 40009 602452 40019 602670
rect 40519 602668 40689 602676
rect 40519 602634 40689 602668
rect 40519 602624 40689 602634
rect 40579 602182 40587 602400
rect 40587 602182 40621 602400
rect 40621 602182 40631 602400
rect 39907 602118 40077 602126
rect 39907 602084 40077 602118
rect 39907 602074 40077 602084
rect 39967 601256 39975 601474
rect 39975 601256 40009 601474
rect 40009 601256 40019 601474
rect 40519 601472 40689 601480
rect 40519 601438 40689 601472
rect 40519 601428 40689 601438
rect 40579 600986 40587 601204
rect 40587 600986 40621 601204
rect 40621 600986 40631 601204
rect 39907 600922 40077 600930
rect 39907 600888 40077 600922
rect 39907 600878 40077 600888
rect 39967 600060 39975 600278
rect 39975 600060 40009 600278
rect 40009 600060 40019 600278
rect 40519 600276 40689 600284
rect 40519 600242 40689 600276
rect 40519 600232 40689 600242
rect 40579 599790 40587 600008
rect 40587 599790 40621 600008
rect 40621 599790 40631 600008
rect 39907 599726 40077 599734
rect 39907 599692 40077 599726
rect 39907 599682 40077 599692
rect 39967 598864 39975 599082
rect 39975 598864 40009 599082
rect 40009 598864 40019 599082
rect 40519 599080 40689 599088
rect 40519 599046 40689 599080
rect 40519 599036 40689 599046
rect 40579 598594 40587 598812
rect 40587 598594 40621 598812
rect 40621 598594 40631 598812
rect 39907 598530 40077 598538
rect 39907 598496 40077 598530
rect 39907 598486 40077 598496
rect 39967 597668 39975 597886
rect 39975 597668 40009 597886
rect 40009 597668 40019 597886
rect 40519 597884 40689 597892
rect 40519 597850 40689 597884
rect 40519 597840 40689 597850
rect 40601 352373 40609 352591
rect 40609 352373 40643 352591
rect 40643 352373 40653 352591
rect 42411 352472 42463 352524
rect 42491 609686 42543 609738
rect 42551 609433 42603 609485
rect 42631 889136 42683 889188
rect 167234 995181 167286 995233
rect 168077 995177 168129 995229
rect 416655 995219 416707 995271
rect 417498 995223 417550 995275
rect 662656 995219 662708 995271
rect 663499 995223 663551 995275
rect 42691 888907 42743 888959
rect 167110 995125 167162 995177
rect 167883 995121 167935 995173
rect 416849 995163 416901 995215
rect 417622 995167 417674 995219
rect 662850 995163 662902 995215
rect 663623 995167 663675 995219
rect 663852 995107 663904 995159
rect 664695 995111 664747 995163
rect 664046 995051 664098 995103
rect 664819 995055 664871 995107
rect 665048 994995 665100 995047
rect 665891 994999 665943 995051
rect 665242 994939 665294 994991
rect 666015 994943 666067 994995
rect 666244 994883 666296 994935
rect 667087 994887 667139 994939
rect 666438 994827 666490 994879
rect 667211 994831 667263 994883
rect 42747 888713 42799 888765
rect 42607 609263 42659 609315
rect 42687 888064 42739 888116
rect 39929 352309 40099 352317
rect 39929 352275 40099 352309
rect 39929 352265 40099 352275
rect 42467 352278 42519 352330
rect 42547 608614 42599 608666
rect 39989 351447 39997 351665
rect 39997 351447 40031 351665
rect 40031 351447 40041 351665
rect 40541 351663 40711 351671
rect 40541 351629 40711 351663
rect 40541 351619 40711 351629
rect 42407 351629 42459 351681
rect 40601 351177 40609 351395
rect 40609 351177 40643 351395
rect 40643 351177 40653 351395
rect 39929 351113 40099 351121
rect 39929 351079 40099 351113
rect 39929 351069 40099 351079
rect 39989 350251 39997 350469
rect 39997 350251 40031 350469
rect 40031 350251 40041 350469
rect 40541 350467 40711 350475
rect 40541 350433 40711 350467
rect 40541 350423 40711 350433
rect 40601 349981 40609 350199
rect 40609 349981 40643 350199
rect 40643 349981 40653 350199
rect 39929 349917 40099 349925
rect 39929 349883 40099 349917
rect 39929 349873 40099 349883
rect 39989 349055 39997 349273
rect 39997 349055 40031 349273
rect 40031 349055 40041 349273
rect 40541 349271 40711 349279
rect 40541 349237 40711 349271
rect 40541 349227 40711 349237
rect 40601 348785 40609 349003
rect 40609 348785 40643 349003
rect 40643 348785 40653 349003
rect 39929 348721 40099 348729
rect 39929 348687 40099 348721
rect 39929 348677 40099 348687
rect 39989 347859 39997 348077
rect 39997 347859 40031 348077
rect 40031 347859 40041 348077
rect 40541 348075 40711 348083
rect 40541 348041 40711 348075
rect 40541 348031 40711 348041
rect 40601 347589 40609 347807
rect 40609 347589 40643 347807
rect 40643 347589 40653 347807
rect 39929 347525 40099 347533
rect 39929 347491 40099 347525
rect 39929 347481 40099 347491
rect 39989 346663 39997 346881
rect 39997 346663 40031 346881
rect 40031 346663 40041 346881
rect 40541 346879 40711 346887
rect 40541 346845 40711 346879
rect 40541 346835 40711 346845
rect 40601 346393 40609 346611
rect 40609 346393 40643 346611
rect 40643 346393 40653 346611
rect 39929 346329 40099 346337
rect 39929 346295 40099 346329
rect 39929 346285 40099 346295
rect 39989 345467 39997 345685
rect 39997 345467 40031 345685
rect 40031 345467 40041 345685
rect 40541 345683 40711 345691
rect 40541 345649 40711 345683
rect 40541 345639 40711 345649
rect 40601 345197 40609 345415
rect 40609 345197 40643 345415
rect 40643 345197 40653 345415
rect 39929 345133 40099 345141
rect 39929 345099 40099 345133
rect 39929 345089 40099 345099
rect 39989 344271 39997 344489
rect 39997 344271 40031 344489
rect 40031 344271 40041 344489
rect 40541 344487 40711 344495
rect 40541 344453 40711 344487
rect 40541 344443 40711 344453
rect 40601 344001 40609 344219
rect 40609 344001 40643 344219
rect 40643 344001 40653 344219
rect 39929 343937 40099 343945
rect 39929 343903 40099 343937
rect 39929 343893 40099 343903
rect 40291 343371 40351 343728
rect 39989 343075 39997 343293
rect 39997 343075 40031 343293
rect 40031 343075 40041 343293
rect 40541 343291 40711 343299
rect 40541 343257 40711 343291
rect 40541 343247 40711 343257
rect 40601 342805 40609 343023
rect 40609 342805 40643 343023
rect 40643 342805 40653 343023
rect 39929 342741 40099 342749
rect 39929 342707 40099 342741
rect 39929 342697 40099 342707
rect 39750 342175 39810 342532
rect 40832 342175 40892 342532
rect 39989 341879 39997 342097
rect 39997 341879 40031 342097
rect 40031 341879 40041 342097
rect 40541 342095 40711 342103
rect 40541 342061 40711 342095
rect 40541 342051 40711 342061
rect 40601 341609 40609 341827
rect 40609 341609 40643 341827
rect 40643 341609 40653 341827
rect 39929 341545 40099 341553
rect 39929 341511 40099 341545
rect 39929 341501 40099 341511
rect 39989 340683 39997 340901
rect 39997 340683 40031 340901
rect 40031 340683 40041 340901
rect 40541 340899 40711 340907
rect 40541 340865 40711 340899
rect 40541 340855 40711 340865
rect 40601 340413 40609 340631
rect 40609 340413 40643 340631
rect 40643 340413 40653 340631
rect 39929 340349 40099 340357
rect 39929 340315 40099 340349
rect 39929 340305 40099 340315
rect 39989 339487 39997 339705
rect 39997 339487 40031 339705
rect 40031 339487 40041 339705
rect 40541 339703 40711 339711
rect 40541 339669 40711 339703
rect 40541 339659 40711 339669
rect 40601 339217 40609 339435
rect 40609 339217 40643 339435
rect 40643 339217 40653 339435
rect 39929 339153 40099 339161
rect 39929 339119 40099 339153
rect 39929 339109 40099 339119
rect 39989 338291 39997 338509
rect 39997 338291 40031 338509
rect 40031 338291 40041 338509
rect 40541 338507 40711 338515
rect 40541 338473 40711 338507
rect 40541 338463 40711 338473
rect 40601 338021 40609 338239
rect 40609 338021 40643 338239
rect 40643 338021 40653 338239
rect 39929 337957 40099 337965
rect 39929 337923 40099 337957
rect 39929 337913 40099 337923
rect 39989 337095 39997 337313
rect 39997 337095 40031 337313
rect 40031 337095 40041 337313
rect 40541 337311 40711 337319
rect 40541 337277 40711 337311
rect 40541 337267 40711 337277
rect 40601 336825 40609 337043
rect 40609 336825 40643 337043
rect 40643 336825 40653 337043
rect 39929 336761 40099 336769
rect 39929 336727 40099 336761
rect 39929 336717 40099 336727
rect 39989 335899 39997 336117
rect 39997 335899 40031 336117
rect 40031 335899 40041 336117
rect 40541 336115 40711 336123
rect 40541 336081 40711 336115
rect 40541 336071 40711 336081
rect 40601 335629 40609 335847
rect 40609 335629 40643 335847
rect 40643 335629 40653 335847
rect 39929 335565 40099 335573
rect 39929 335531 40099 335565
rect 39929 335521 40099 335531
rect 39989 334703 39997 334921
rect 39997 334703 40031 334921
rect 40031 334703 40041 334921
rect 40541 334919 40711 334927
rect 40541 334885 40711 334919
rect 40541 334875 40711 334885
rect 42463 351505 42515 351557
rect 42523 351252 42575 351304
rect 42603 608490 42655 608542
rect 42663 608261 42715 608313
rect 42743 887940 42795 887992
rect 42803 887687 42855 887739
rect 42859 887517 42911 887569
rect 42719 608067 42771 608119
rect 42799 886868 42851 886920
rect 42579 351082 42631 351134
rect 42659 607418 42711 607470
rect 42519 350433 42571 350485
rect 42575 350309 42627 350361
rect 42635 350080 42687 350132
rect 42715 607294 42767 607346
rect 42775 607041 42827 607093
rect 42855 886744 42907 886796
rect 42915 886515 42967 886567
rect 42971 886321 43023 886373
rect 42831 606871 42883 606923
rect 42911 885672 42963 885724
rect 42691 349886 42743 349938
rect 42771 606222 42823 606274
rect 42631 349237 42683 349289
rect 42687 349113 42739 349165
rect 42747 348860 42799 348912
rect 42827 606098 42879 606150
rect 42887 605869 42939 605921
rect 42967 885548 43019 885600
rect 675092 714315 675144 714367
rect 676928 714240 676938 714458
rect 676938 714240 676972 714458
rect 676972 714240 676980 714458
rect 675036 714145 675088 714197
rect 677482 714176 677652 714184
rect 677482 714142 677652 714176
rect 677482 714132 677652 714142
rect 675096 713496 675148 713548
rect 675040 713372 675092 713424
rect 674980 713143 675032 713195
rect 674924 712949 674976 713001
rect 674984 712300 675036 712352
rect 674928 712176 674980 712228
rect 674868 711947 674920 711999
rect 674812 711753 674864 711805
rect 674872 711104 674924 711156
rect 674816 710980 674868 711032
rect 674756 710751 674808 710803
rect 674700 710557 674752 710609
rect 674760 709908 674812 709960
rect 674704 709784 674756 709836
rect 674644 709555 674696 709607
rect 674588 709361 674640 709413
rect 674648 708712 674700 708764
rect 674592 708588 674644 708640
rect 674532 708359 674584 708411
rect 674476 708165 674528 708217
rect 674536 707516 674588 707568
rect 674480 707392 674532 707444
rect 42943 605675 42995 605727
rect 42803 348690 42855 348742
rect 42883 605026 42935 605078
rect 42743 348041 42795 348093
rect 42799 347917 42851 347969
rect 42859 347688 42911 347740
rect 42939 604902 42991 604954
rect 42999 604673 43051 604725
rect 43055 604479 43107 604531
rect 42915 347494 42967 347546
rect 42995 603830 43047 603882
rect 42855 346845 42907 346897
rect 42911 346721 42963 346773
rect 42971 346492 43023 346544
rect 43051 603706 43103 603758
rect 43111 603477 43163 603529
rect 43167 603283 43219 603335
rect 43027 346298 43079 346350
rect 43107 602634 43159 602686
rect 42967 345649 43019 345701
rect 43023 345525 43075 345577
rect 43083 345296 43135 345348
rect 43163 602510 43215 602562
rect 43223 602281 43275 602333
rect 43279 602087 43331 602139
rect 43139 345102 43191 345154
rect 43219 601438 43271 601490
rect 43079 344453 43131 344505
rect 43135 344329 43187 344381
rect 43195 344100 43247 344152
rect 43275 601314 43327 601366
rect 43335 601085 43387 601137
rect 43391 600891 43443 600943
rect 43251 343906 43303 343958
rect 43331 600242 43383 600294
rect 43191 343257 43243 343309
rect 43247 343133 43299 343185
rect 43307 342904 43359 342956
rect 43387 600118 43439 600170
rect 43447 599889 43499 599941
rect 43503 599695 43555 599747
rect 43363 342710 43415 342762
rect 43443 599046 43495 599098
rect 43303 342061 43355 342113
rect 43359 341937 43411 341989
rect 43419 341708 43471 341760
rect 43499 598922 43551 598974
rect 43559 598693 43611 598745
rect 43615 598499 43667 598551
rect 43475 341514 43527 341566
rect 43555 597850 43607 597902
rect 43415 340865 43467 340917
rect 43471 340741 43523 340793
rect 43531 340512 43583 340564
rect 43611 597726 43663 597778
rect 676870 713530 677040 713538
rect 676870 713496 677040 713530
rect 676870 713486 677040 713496
rect 677540 713314 677550 713532
rect 677550 713314 677584 713532
rect 677584 713314 677592 713532
rect 676928 713044 676938 713262
rect 676938 713044 676972 713262
rect 676972 713044 676980 713262
rect 677482 712980 677652 712988
rect 677482 712946 677652 712980
rect 677482 712936 677652 712946
rect 676870 712334 677040 712342
rect 676870 712300 677040 712334
rect 676870 712290 677040 712300
rect 677540 712118 677550 712336
rect 677550 712118 677584 712336
rect 677584 712118 677592 712336
rect 676928 711848 676938 712066
rect 676938 711848 676972 712066
rect 676972 711848 676980 712066
rect 677482 711784 677652 711792
rect 677482 711750 677652 711784
rect 677482 711740 677652 711750
rect 676693 711296 676753 711653
rect 677775 711296 677835 711653
rect 676870 711138 677040 711146
rect 676870 711104 677040 711138
rect 676870 711094 677040 711104
rect 677540 710922 677550 711140
rect 677550 710922 677584 711140
rect 677584 710922 677592 711140
rect 676928 710652 676938 710870
rect 676938 710652 676972 710870
rect 676972 710652 676980 710870
rect 677482 710588 677652 710596
rect 677482 710554 677652 710588
rect 677482 710544 677652 710554
rect 677234 710100 677294 710457
rect 676870 709942 677040 709950
rect 676870 709908 677040 709942
rect 676870 709898 677040 709908
rect 677540 709726 677550 709944
rect 677550 709726 677584 709944
rect 677584 709726 677592 709944
rect 676928 709456 676938 709674
rect 676938 709456 676972 709674
rect 676972 709456 676980 709674
rect 677482 709392 677652 709400
rect 677482 709358 677652 709392
rect 677482 709348 677652 709358
rect 676870 708746 677040 708754
rect 676870 708712 677040 708746
rect 676870 708702 677040 708712
rect 677540 708530 677550 708748
rect 677550 708530 677584 708748
rect 677584 708530 677592 708748
rect 676928 708260 676938 708478
rect 676938 708260 676972 708478
rect 676972 708260 676980 708478
rect 677482 708196 677652 708204
rect 677482 708162 677652 708196
rect 677482 708152 677652 708162
rect 676870 707550 677040 707558
rect 676870 707516 677040 707550
rect 676870 707506 677040 707516
rect 677540 707334 677550 707552
rect 677550 707334 677584 707552
rect 677584 707334 677592 707552
rect 675092 453515 675144 453567
rect 676928 453416 676938 453634
rect 676938 453416 676972 453634
rect 676972 453416 676980 453634
rect 675036 453321 675088 453373
rect 677482 453352 677652 453360
rect 677482 453318 677652 453352
rect 677482 453308 677652 453318
rect 675096 452672 675148 452724
rect 675040 452548 675092 452600
rect 674980 452295 675032 452347
rect 674924 452125 674976 452177
rect 674984 451476 675036 451528
rect 674928 451352 674980 451404
rect 674868 451123 674920 451175
rect 674812 450929 674864 450981
rect 674872 450280 674924 450332
rect 674816 450156 674868 450208
rect 674756 449903 674808 449955
rect 674700 449733 674752 449785
rect 674760 449084 674812 449136
rect 674704 448960 674756 449012
rect 674644 448731 674696 448783
rect 674588 448537 674640 448589
rect 674648 447888 674700 447940
rect 674592 447764 674644 447816
rect 674532 447535 674584 447587
rect 674476 447341 674528 447393
rect 674536 446692 674588 446744
rect 674480 446568 674532 446620
rect 674420 446339 674472 446391
rect 674364 446145 674416 446197
rect 674424 445496 674476 445548
rect 674368 445372 674420 445424
rect 674308 445143 674360 445195
rect 674252 444949 674304 445001
rect 674312 444300 674364 444352
rect 674256 444176 674308 444228
rect 674196 443947 674248 443999
rect 674140 443753 674192 443805
rect 674200 443104 674252 443156
rect 674144 442980 674196 443032
rect 674084 442751 674136 442803
rect 674028 442557 674080 442609
rect 674088 441908 674140 441960
rect 674032 441784 674084 441836
rect 673972 441555 674024 441607
rect 673916 441361 673968 441413
rect 673976 440712 674028 440764
rect 673920 440588 673972 440640
rect 673860 440359 673912 440411
rect 673804 440165 673856 440217
rect 673864 439516 673916 439568
rect 673808 439392 673860 439444
rect 43587 340318 43639 340370
rect 43527 339669 43579 339721
rect 43583 339545 43635 339597
rect 43643 339316 43695 339368
rect 43699 339122 43751 339174
rect 43639 338473 43691 338525
rect 43695 338349 43747 338401
rect 43755 338120 43807 338172
rect 43811 337926 43863 337978
rect 43751 337277 43803 337329
rect 43807 337153 43859 337205
rect 43867 336900 43919 336952
rect 43923 336730 43975 336782
rect 43863 336081 43915 336133
rect 43919 335957 43971 336009
rect 43979 335728 44031 335780
rect 44035 335534 44087 335586
rect 43975 334885 44027 334937
rect 44031 334761 44083 334813
rect 134104 225848 134156 225900
rect 134947 225852 134999 225904
rect 394104 225876 394156 225928
rect 394947 225880 394999 225932
rect 135176 225792 135228 225844
rect 135949 225796 136001 225848
rect 395176 225820 395228 225872
rect 395949 225824 396001 225876
rect 135300 225736 135352 225788
rect 136143 225740 136195 225792
rect 395300 225764 395352 225816
rect 396143 225768 396195 225820
rect 136372 225680 136424 225732
rect 137145 225684 137197 225736
rect 396372 225708 396424 225760
rect 397145 225712 397197 225764
rect 136496 225624 136548 225676
rect 137339 225628 137391 225680
rect 396496 225652 396548 225704
rect 397339 225656 397391 225708
rect 137568 225568 137620 225620
rect 138341 225572 138393 225624
rect 397568 225596 397620 225648
rect 398341 225600 398393 225652
rect 137692 225512 137744 225564
rect 138535 225516 138587 225568
rect 397692 225540 397744 225592
rect 398535 225544 398587 225596
rect 138764 225456 138816 225508
rect 139537 225460 139589 225512
rect 398764 225484 398816 225536
rect 399537 225488 399589 225540
rect 138888 225400 138940 225452
rect 139731 225404 139783 225456
rect 398888 225428 398940 225480
rect 399731 225432 399783 225484
rect 139960 225344 140012 225396
rect 140733 225348 140785 225400
rect 399960 225372 400012 225424
rect 400733 225376 400785 225428
rect 140084 225288 140136 225340
rect 140903 225292 140955 225344
rect 400084 225316 400136 225368
rect 400903 225320 400955 225372
rect 141156 225232 141208 225284
rect 141929 225236 141981 225288
rect 401156 225260 401208 225312
rect 401929 225264 401981 225316
rect 141280 225176 141332 225228
rect 142123 225180 142175 225232
rect 401280 225204 401332 225256
rect 402123 225208 402175 225260
rect 142352 225120 142404 225172
rect 143125 225124 143177 225176
rect 402352 225148 402404 225200
rect 403125 225152 403177 225204
rect 142476 225064 142528 225116
rect 143295 225068 143347 225120
rect 402476 225092 402528 225144
rect 403295 225096 403347 225148
rect 143548 225008 143600 225060
rect 144321 225012 144373 225064
rect 403548 225036 403600 225088
rect 404321 225040 404373 225092
rect 143672 224952 143724 225004
rect 144515 224956 144567 225008
rect 403672 224980 403724 225032
rect 404515 224984 404567 225036
rect 144744 224896 144796 224948
rect 145517 224900 145569 224952
rect 404744 224924 404796 224976
rect 405517 224928 405569 224980
rect 144868 224840 144920 224892
rect 145711 224844 145763 224896
rect 404868 224868 404920 224920
rect 405711 224872 405763 224924
rect 145940 224784 145992 224836
rect 146713 224788 146765 224840
rect 405940 224812 405992 224864
rect 406713 224816 406765 224868
rect 146064 224728 146116 224780
rect 146907 224732 146959 224784
rect 406064 224756 406116 224808
rect 406907 224760 406959 224812
rect 147136 224672 147188 224724
rect 147909 224676 147961 224728
rect 407136 224700 407188 224752
rect 407909 224704 407961 224756
rect 147260 224616 147312 224668
rect 148103 224620 148155 224672
rect 407260 224644 407312 224696
rect 408103 224648 408155 224700
rect 148332 224560 148384 224612
rect 149105 224564 149157 224616
rect 408332 224588 408384 224640
rect 409105 224592 409157 224644
rect 148456 224504 148508 224556
rect 149299 224508 149351 224560
rect 408456 224532 408508 224584
rect 409299 224536 409351 224588
rect 149528 224448 149580 224500
rect 150301 224452 150353 224504
rect 409528 224476 409580 224528
rect 410301 224480 410353 224532
rect 149652 224392 149704 224444
rect 150495 224396 150547 224448
rect 409652 224420 409704 224472
rect 410495 224424 410547 224476
rect 150724 224336 150776 224388
rect 151497 224340 151549 224392
rect 410724 224364 410776 224416
rect 411497 224368 411549 224420
rect 150848 224280 150900 224332
rect 151691 224284 151743 224336
rect 410848 224308 410900 224360
rect 411691 224312 411743 224364
rect 151920 224224 151972 224276
rect 152693 224228 152745 224280
rect 411920 224252 411972 224304
rect 412693 224256 412745 224308
rect 152044 224168 152096 224220
rect 152887 224172 152939 224224
rect 412044 224196 412096 224248
rect 412887 224200 412939 224252
rect 153116 224112 153168 224164
rect 153889 224116 153941 224168
rect 413116 224140 413168 224192
rect 413889 224144 413941 224196
rect 153240 224056 153292 224108
rect 154083 224060 154135 224112
rect 413240 224084 413292 224136
rect 414083 224088 414135 224140
rect 154312 224000 154364 224052
rect 155085 224004 155137 224056
rect 414312 224028 414364 224080
rect 415085 224032 415137 224084
rect 154436 223944 154488 223996
rect 155255 223948 155307 224000
rect 414436 223972 414488 224024
rect 415255 223976 415307 224028
rect 155508 223888 155560 223940
rect 156281 223892 156333 223944
rect 415508 223916 415560 223968
rect 416281 223920 416333 223972
rect 155632 223832 155684 223884
rect 156475 223836 156527 223888
rect 415632 223860 415684 223912
rect 416475 223864 416527 223916
rect 156704 223776 156756 223828
rect 157477 223780 157529 223832
rect 416704 223804 416756 223856
rect 417477 223808 417529 223860
rect 156828 223720 156880 223772
rect 157647 223724 157699 223776
rect 416828 223748 416880 223800
rect 417647 223752 417699 223804
rect 157900 223664 157952 223716
rect 158673 223668 158725 223720
rect 417900 223692 417952 223744
rect 418673 223696 418725 223748
rect 158024 223608 158076 223660
rect 158867 223612 158919 223664
rect 418024 223636 418076 223688
rect 418867 223640 418919 223692
rect 147395 223397 147752 223457
rect 406226 223390 406583 223450
rect 134094 223102 134104 223272
rect 134104 223102 134138 223272
rect 134138 223102 134146 223272
rect 134848 223204 135066 223214
rect 134848 223170 135066 223204
rect 134848 223162 135066 223170
rect 135290 223102 135300 223272
rect 135300 223102 135334 223272
rect 135334 223102 135342 223272
rect 136044 223204 136262 223214
rect 136044 223170 136262 223204
rect 136044 223162 136262 223170
rect 136486 223102 136496 223272
rect 136496 223102 136530 223272
rect 136530 223102 136538 223272
rect 137240 223204 137458 223214
rect 137240 223170 137458 223204
rect 137240 223162 137458 223170
rect 137682 223102 137692 223272
rect 137692 223102 137726 223272
rect 137726 223102 137734 223272
rect 138436 223204 138654 223214
rect 138436 223170 138654 223204
rect 138436 223162 138654 223170
rect 138878 223102 138888 223272
rect 138888 223102 138922 223272
rect 138922 223102 138930 223272
rect 139632 223204 139850 223214
rect 139632 223170 139850 223204
rect 139632 223162 139850 223170
rect 140074 223102 140084 223272
rect 140084 223102 140118 223272
rect 140118 223102 140126 223272
rect 140828 223204 141046 223214
rect 140828 223170 141046 223204
rect 140828 223162 141046 223170
rect 141270 223102 141280 223272
rect 141280 223102 141314 223272
rect 141314 223102 141322 223272
rect 142024 223204 142242 223214
rect 142024 223170 142242 223204
rect 142024 223162 142242 223170
rect 142466 223102 142476 223272
rect 142476 223102 142510 223272
rect 142510 223102 142518 223272
rect 143220 223204 143438 223214
rect 143220 223170 143438 223204
rect 143220 223162 143438 223170
rect 143662 223102 143672 223272
rect 143672 223102 143706 223272
rect 143706 223102 143714 223272
rect 144416 223204 144634 223214
rect 144416 223170 144634 223204
rect 144416 223162 144634 223170
rect 144858 223102 144868 223272
rect 144868 223102 144902 223272
rect 144902 223102 144910 223272
rect 145612 223204 145830 223214
rect 145612 223170 145830 223204
rect 145612 223162 145830 223170
rect 146054 223102 146064 223272
rect 146064 223102 146098 223272
rect 146098 223102 146106 223272
rect 146808 223204 147026 223214
rect 146808 223170 147026 223204
rect 146808 223162 147026 223170
rect 147250 223102 147260 223272
rect 147260 223102 147294 223272
rect 147294 223102 147302 223272
rect 148004 223204 148222 223214
rect 148004 223170 148222 223204
rect 148004 223162 148222 223170
rect 148446 223102 148456 223272
rect 148456 223102 148490 223272
rect 148490 223102 148498 223272
rect 149200 223204 149418 223214
rect 149200 223170 149418 223204
rect 149200 223162 149418 223170
rect 149642 223102 149652 223272
rect 149652 223102 149686 223272
rect 149686 223102 149694 223272
rect 150396 223204 150614 223214
rect 150396 223170 150614 223204
rect 150396 223162 150614 223170
rect 150838 223102 150848 223272
rect 150848 223102 150882 223272
rect 150882 223102 150890 223272
rect 151592 223204 151810 223214
rect 151592 223170 151810 223204
rect 151592 223162 151810 223170
rect 152034 223102 152044 223272
rect 152044 223102 152078 223272
rect 152078 223102 152086 223272
rect 152788 223204 153006 223214
rect 152788 223170 153006 223204
rect 152788 223162 153006 223170
rect 153230 223102 153240 223272
rect 153240 223102 153274 223272
rect 153274 223102 153282 223272
rect 153984 223204 154202 223214
rect 153984 223170 154202 223204
rect 153984 223162 154202 223170
rect 154426 223102 154436 223272
rect 154436 223102 154470 223272
rect 154470 223102 154478 223272
rect 155180 223204 155398 223214
rect 155180 223170 155398 223204
rect 155180 223162 155398 223170
rect 155622 223102 155632 223272
rect 155632 223102 155666 223272
rect 155666 223102 155674 223272
rect 156376 223204 156594 223214
rect 156376 223170 156594 223204
rect 156376 223162 156594 223170
rect 156818 223102 156828 223272
rect 156828 223102 156862 223272
rect 156862 223102 156870 223272
rect 157572 223204 157790 223214
rect 157572 223170 157790 223204
rect 157572 223162 157790 223170
rect 158014 223102 158024 223272
rect 158024 223102 158058 223272
rect 158058 223102 158066 223272
rect 158768 223204 158986 223214
rect 158768 223170 158986 223204
rect 158768 223162 158986 223170
rect 394094 223102 394104 223272
rect 394104 223102 394138 223272
rect 394138 223102 394146 223272
rect 394848 223204 395066 223214
rect 394848 223170 395066 223204
rect 394848 223162 395066 223170
rect 395290 223102 395300 223272
rect 395300 223102 395334 223272
rect 395334 223102 395342 223272
rect 396044 223204 396262 223214
rect 396044 223170 396262 223204
rect 396044 223162 396262 223170
rect 396486 223102 396496 223272
rect 396496 223102 396530 223272
rect 396530 223102 396538 223272
rect 397240 223204 397458 223214
rect 397240 223170 397458 223204
rect 397240 223162 397458 223170
rect 397682 223102 397692 223272
rect 397692 223102 397726 223272
rect 397726 223102 397734 223272
rect 398436 223204 398654 223214
rect 398436 223170 398654 223204
rect 398436 223162 398654 223170
rect 398878 223102 398888 223272
rect 398888 223102 398922 223272
rect 398922 223102 398930 223272
rect 399632 223204 399850 223214
rect 399632 223170 399850 223204
rect 399632 223162 399850 223170
rect 400074 223102 400084 223272
rect 400084 223102 400118 223272
rect 400118 223102 400126 223272
rect 400828 223204 401046 223214
rect 400828 223170 401046 223204
rect 400828 223162 401046 223170
rect 401270 223102 401280 223272
rect 401280 223102 401314 223272
rect 401314 223102 401322 223272
rect 402024 223204 402242 223214
rect 402024 223170 402242 223204
rect 402024 223162 402242 223170
rect 402466 223102 402476 223272
rect 402476 223102 402510 223272
rect 402510 223102 402518 223272
rect 403220 223204 403438 223214
rect 403220 223170 403438 223204
rect 403220 223162 403438 223170
rect 403662 223102 403672 223272
rect 403672 223102 403706 223272
rect 403706 223102 403714 223272
rect 404416 223204 404634 223214
rect 404416 223170 404634 223204
rect 404416 223162 404634 223170
rect 404858 223102 404868 223272
rect 404868 223102 404902 223272
rect 404902 223102 404910 223272
rect 405612 223204 405830 223214
rect 405612 223170 405830 223204
rect 405612 223162 405830 223170
rect 406054 223102 406064 223272
rect 406064 223102 406098 223272
rect 406098 223102 406106 223272
rect 406808 223204 407026 223214
rect 406808 223170 407026 223204
rect 406808 223162 407026 223170
rect 407250 223102 407260 223272
rect 407260 223102 407294 223272
rect 407294 223102 407302 223272
rect 408004 223204 408222 223214
rect 408004 223170 408222 223204
rect 408004 223162 408222 223170
rect 408446 223102 408456 223272
rect 408456 223102 408490 223272
rect 408490 223102 408498 223272
rect 409200 223204 409418 223214
rect 409200 223170 409418 223204
rect 409200 223162 409418 223170
rect 409642 223102 409652 223272
rect 409652 223102 409686 223272
rect 409686 223102 409694 223272
rect 410396 223204 410614 223214
rect 410396 223170 410614 223204
rect 410396 223162 410614 223170
rect 410838 223102 410848 223272
rect 410848 223102 410882 223272
rect 410882 223102 410890 223272
rect 411592 223204 411810 223214
rect 411592 223170 411810 223204
rect 411592 223162 411810 223170
rect 412034 223102 412044 223272
rect 412044 223102 412078 223272
rect 412078 223102 412086 223272
rect 412788 223204 413006 223214
rect 412788 223170 413006 223204
rect 412788 223162 413006 223170
rect 413230 223102 413240 223272
rect 413240 223102 413274 223272
rect 413274 223102 413282 223272
rect 413984 223204 414202 223214
rect 413984 223170 414202 223204
rect 413984 223162 414202 223170
rect 414426 223102 414436 223272
rect 414436 223102 414470 223272
rect 414470 223102 414478 223272
rect 415180 223204 415398 223214
rect 415180 223170 415398 223204
rect 415180 223162 415398 223170
rect 415622 223102 415632 223272
rect 415632 223102 415666 223272
rect 415666 223102 415674 223272
rect 416376 223204 416594 223214
rect 416376 223170 416594 223204
rect 416376 223162 416594 223170
rect 416818 223102 416828 223272
rect 416828 223102 416862 223272
rect 416862 223102 416870 223272
rect 417572 223204 417790 223214
rect 417572 223170 417790 223204
rect 417572 223162 417790 223170
rect 418014 223102 418024 223272
rect 418024 223102 418058 223272
rect 418058 223102 418066 223272
rect 418768 223204 418986 223214
rect 418768 223170 418986 223204
rect 418768 223162 418986 223170
rect 146199 222856 146556 222916
rect 405030 222849 405387 222909
rect 135118 222592 135336 222602
rect 135118 222558 135336 222592
rect 135118 222550 135336 222558
rect 135936 222490 135946 222660
rect 135946 222490 135980 222660
rect 135980 222490 135988 222660
rect 136314 222592 136532 222602
rect 136314 222558 136532 222592
rect 136314 222550 136532 222558
rect 137132 222490 137142 222660
rect 137142 222490 137176 222660
rect 137176 222490 137184 222660
rect 137510 222592 137728 222602
rect 137510 222558 137728 222592
rect 137510 222550 137728 222558
rect 138328 222490 138338 222660
rect 138338 222490 138372 222660
rect 138372 222490 138380 222660
rect 138706 222592 138924 222602
rect 138706 222558 138924 222592
rect 138706 222550 138924 222558
rect 139524 222490 139534 222660
rect 139534 222490 139568 222660
rect 139568 222490 139576 222660
rect 139902 222592 140120 222602
rect 139902 222558 140120 222592
rect 139902 222550 140120 222558
rect 140720 222490 140730 222660
rect 140730 222490 140764 222660
rect 140764 222490 140772 222660
rect 141098 222592 141316 222602
rect 141098 222558 141316 222592
rect 141098 222550 141316 222558
rect 141916 222490 141926 222660
rect 141926 222490 141960 222660
rect 141960 222490 141968 222660
rect 142294 222592 142512 222602
rect 142294 222558 142512 222592
rect 142294 222550 142512 222558
rect 143112 222490 143122 222660
rect 143122 222490 143156 222660
rect 143156 222490 143164 222660
rect 143490 222592 143708 222602
rect 143490 222558 143708 222592
rect 143490 222550 143708 222558
rect 144308 222490 144318 222660
rect 144318 222490 144352 222660
rect 144352 222490 144360 222660
rect 144686 222592 144904 222602
rect 144686 222558 144904 222592
rect 144686 222550 144904 222558
rect 145504 222490 145514 222660
rect 145514 222490 145548 222660
rect 145548 222490 145556 222660
rect 145882 222592 146100 222602
rect 145882 222558 146100 222592
rect 145882 222550 146100 222558
rect 146700 222490 146710 222660
rect 146710 222490 146744 222660
rect 146744 222490 146752 222660
rect 147078 222592 147296 222602
rect 147078 222558 147296 222592
rect 147078 222550 147296 222558
rect 147896 222490 147906 222660
rect 147906 222490 147940 222660
rect 147940 222490 147948 222660
rect 148274 222592 148492 222602
rect 148274 222558 148492 222592
rect 148274 222550 148492 222558
rect 149092 222490 149102 222660
rect 149102 222490 149136 222660
rect 149136 222490 149144 222660
rect 149470 222592 149688 222602
rect 149470 222558 149688 222592
rect 149470 222550 149688 222558
rect 150288 222490 150298 222660
rect 150298 222490 150332 222660
rect 150332 222490 150340 222660
rect 150666 222592 150884 222602
rect 150666 222558 150884 222592
rect 150666 222550 150884 222558
rect 151484 222490 151494 222660
rect 151494 222490 151528 222660
rect 151528 222490 151536 222660
rect 151862 222592 152080 222602
rect 151862 222558 152080 222592
rect 151862 222550 152080 222558
rect 152680 222490 152690 222660
rect 152690 222490 152724 222660
rect 152724 222490 152732 222660
rect 153058 222592 153276 222602
rect 153058 222558 153276 222592
rect 153058 222550 153276 222558
rect 153876 222490 153886 222660
rect 153886 222490 153920 222660
rect 153920 222490 153928 222660
rect 154254 222592 154472 222602
rect 154254 222558 154472 222592
rect 154254 222550 154472 222558
rect 155072 222490 155082 222660
rect 155082 222490 155116 222660
rect 155116 222490 155124 222660
rect 155450 222592 155668 222602
rect 155450 222558 155668 222592
rect 155450 222550 155668 222558
rect 156268 222490 156278 222660
rect 156278 222490 156312 222660
rect 156312 222490 156320 222660
rect 156646 222592 156864 222602
rect 156646 222558 156864 222592
rect 156646 222550 156864 222558
rect 157464 222490 157474 222660
rect 157474 222490 157508 222660
rect 157508 222490 157516 222660
rect 158016 222490 158024 222660
rect 158024 222490 158058 222660
rect 158058 222490 158068 222660
rect 158668 222592 158886 222602
rect 158668 222558 158886 222592
rect 158668 222550 158886 222558
rect 395118 222592 395336 222602
rect 395118 222558 395336 222592
rect 395118 222550 395336 222558
rect 395936 222490 395946 222660
rect 395946 222490 395980 222660
rect 395980 222490 395988 222660
rect 396314 222592 396532 222602
rect 396314 222558 396532 222592
rect 396314 222550 396532 222558
rect 397132 222490 397142 222660
rect 397142 222490 397176 222660
rect 397176 222490 397184 222660
rect 397510 222592 397728 222602
rect 397510 222558 397728 222592
rect 397510 222550 397728 222558
rect 398328 222490 398338 222660
rect 398338 222490 398372 222660
rect 398372 222490 398380 222660
rect 398706 222592 398924 222602
rect 398706 222558 398924 222592
rect 398706 222550 398924 222558
rect 399524 222490 399534 222660
rect 399534 222490 399568 222660
rect 399568 222490 399576 222660
rect 399902 222592 400120 222602
rect 399902 222558 400120 222592
rect 399902 222550 400120 222558
rect 400720 222490 400730 222660
rect 400730 222490 400764 222660
rect 400764 222490 400772 222660
rect 401098 222592 401316 222602
rect 401098 222558 401316 222592
rect 401098 222550 401316 222558
rect 401916 222490 401926 222660
rect 401926 222490 401960 222660
rect 401960 222490 401968 222660
rect 402294 222592 402512 222602
rect 402294 222558 402512 222592
rect 402294 222550 402512 222558
rect 403112 222490 403122 222660
rect 403122 222490 403156 222660
rect 403156 222490 403164 222660
rect 403490 222592 403708 222602
rect 403490 222558 403708 222592
rect 403490 222550 403708 222558
rect 404308 222490 404318 222660
rect 404318 222490 404352 222660
rect 404352 222490 404360 222660
rect 404686 222592 404904 222602
rect 404686 222558 404904 222592
rect 404686 222550 404904 222558
rect 405504 222490 405514 222660
rect 405514 222490 405548 222660
rect 405548 222490 405556 222660
rect 405882 222592 406100 222602
rect 405882 222558 406100 222592
rect 405882 222550 406100 222558
rect 406700 222490 406710 222660
rect 406710 222490 406744 222660
rect 406744 222490 406752 222660
rect 407078 222592 407296 222602
rect 407078 222558 407296 222592
rect 407078 222550 407296 222558
rect 407896 222490 407906 222660
rect 407906 222490 407940 222660
rect 407940 222490 407948 222660
rect 408274 222592 408492 222602
rect 408274 222558 408492 222592
rect 408274 222550 408492 222558
rect 409092 222490 409102 222660
rect 409102 222490 409136 222660
rect 409136 222490 409144 222660
rect 409470 222592 409688 222602
rect 409470 222558 409688 222592
rect 409470 222550 409688 222558
rect 410288 222490 410298 222660
rect 410298 222490 410332 222660
rect 410332 222490 410340 222660
rect 410666 222592 410884 222602
rect 410666 222558 410884 222592
rect 410666 222550 410884 222558
rect 411484 222490 411494 222660
rect 411494 222490 411528 222660
rect 411528 222490 411536 222660
rect 411862 222592 412080 222602
rect 411862 222558 412080 222592
rect 411862 222550 412080 222558
rect 412680 222490 412690 222660
rect 412690 222490 412724 222660
rect 412724 222490 412732 222660
rect 413058 222592 413276 222602
rect 413058 222558 413276 222592
rect 413058 222550 413276 222558
rect 413876 222490 413886 222660
rect 413886 222490 413920 222660
rect 413920 222490 413928 222660
rect 414254 222592 414472 222602
rect 414254 222558 414472 222592
rect 414254 222550 414472 222558
rect 415072 222490 415082 222660
rect 415082 222490 415116 222660
rect 415116 222490 415124 222660
rect 415450 222592 415668 222602
rect 415450 222558 415668 222592
rect 415450 222550 415668 222558
rect 416268 222490 416278 222660
rect 416278 222490 416312 222660
rect 416312 222490 416320 222660
rect 416646 222592 416864 222602
rect 416646 222558 416864 222592
rect 416646 222550 416864 222558
rect 417464 222490 417474 222660
rect 417474 222490 417508 222660
rect 417508 222490 417516 222660
rect 418016 222490 418024 222660
rect 418024 222490 418058 222660
rect 418058 222490 418068 222660
rect 418668 222592 418886 222602
rect 418668 222558 418886 222592
rect 418668 222550 418886 222558
rect 147395 222315 147752 222375
rect 406226 222308 406583 222368
rect 676870 452706 677040 452714
rect 676870 452672 677040 452706
rect 676870 452662 677040 452672
rect 677540 452490 677550 452708
rect 677550 452490 677584 452708
rect 677584 452490 677592 452708
rect 676928 452220 676938 452438
rect 676938 452220 676972 452438
rect 676972 452220 676980 452438
rect 677482 452156 677652 452164
rect 677482 452122 677652 452156
rect 677482 452112 677652 452122
rect 676870 451510 677040 451518
rect 676870 451476 677040 451510
rect 676870 451466 677040 451476
rect 677540 451294 677550 451512
rect 677550 451294 677584 451512
rect 677584 451294 677592 451512
rect 676928 451024 676938 451242
rect 676938 451024 676972 451242
rect 676972 451024 676980 451242
rect 677482 450960 677652 450968
rect 677482 450926 677652 450960
rect 677482 450916 677652 450926
rect 676870 450314 677040 450322
rect 676870 450280 677040 450314
rect 676870 450270 677040 450280
rect 677540 450098 677550 450316
rect 677550 450098 677584 450316
rect 677584 450098 677592 450316
rect 676928 449828 676938 450046
rect 676938 449828 676972 450046
rect 676972 449828 676980 450046
rect 677482 449764 677652 449772
rect 677482 449730 677652 449764
rect 677482 449720 677652 449730
rect 676870 449118 677040 449126
rect 676870 449084 677040 449118
rect 676870 449074 677040 449084
rect 677540 448902 677550 449120
rect 677550 448902 677584 449120
rect 677584 448902 677592 449120
rect 676928 448632 676938 448850
rect 676938 448632 676972 448850
rect 676972 448632 676980 448850
rect 677482 448568 677652 448576
rect 677482 448534 677652 448568
rect 677482 448524 677652 448534
rect 676685 448095 676745 448452
rect 677767 448095 677827 448452
rect 676870 447922 677040 447930
rect 676870 447888 677040 447922
rect 676870 447878 677040 447888
rect 677540 447706 677550 447924
rect 677550 447706 677584 447924
rect 677584 447706 677592 447924
rect 676928 447436 676938 447654
rect 676938 447436 676972 447654
rect 676972 447436 676980 447654
rect 677482 447372 677652 447380
rect 677482 447338 677652 447372
rect 677482 447328 677652 447338
rect 677226 446899 677286 447256
rect 676870 446726 677040 446734
rect 676870 446692 677040 446726
rect 676870 446682 677040 446692
rect 677540 446510 677550 446728
rect 677550 446510 677584 446728
rect 677584 446510 677592 446728
rect 676928 446240 676938 446458
rect 676938 446240 676972 446458
rect 676972 446240 676980 446458
rect 677482 446176 677652 446184
rect 677482 446142 677652 446176
rect 677482 446132 677652 446142
rect 676870 445530 677040 445538
rect 676870 445496 677040 445530
rect 676870 445486 677040 445496
rect 677540 445314 677550 445532
rect 677550 445314 677584 445532
rect 677584 445314 677592 445532
rect 676928 445044 676938 445262
rect 676938 445044 676972 445262
rect 676972 445044 676980 445262
rect 677482 444980 677652 444988
rect 677482 444946 677652 444980
rect 677482 444936 677652 444946
rect 676870 444334 677040 444342
rect 676870 444300 677040 444334
rect 676870 444290 677040 444300
rect 677540 444118 677550 444336
rect 677550 444118 677584 444336
rect 677584 444118 677592 444336
rect 676928 443848 676938 444066
rect 676938 443848 676972 444066
rect 676972 443848 676980 444066
rect 677482 443784 677652 443792
rect 677482 443750 677652 443784
rect 677482 443740 677652 443750
rect 676870 443138 677040 443146
rect 676870 443104 677040 443138
rect 676870 443094 677040 443104
rect 677540 442922 677550 443140
rect 677550 442922 677584 443140
rect 677584 442922 677592 443140
rect 676928 442652 676938 442870
rect 676938 442652 676972 442870
rect 676972 442652 676980 442870
rect 677482 442588 677652 442596
rect 677482 442554 677652 442588
rect 677482 442544 677652 442554
rect 676870 441942 677040 441950
rect 676870 441908 677040 441942
rect 676870 441898 677040 441908
rect 677540 441726 677550 441944
rect 677550 441726 677584 441944
rect 677584 441726 677592 441944
rect 676928 441456 676938 441674
rect 676938 441456 676972 441674
rect 676972 441456 676980 441674
rect 677482 441392 677652 441400
rect 677482 441358 677652 441392
rect 677482 441348 677652 441358
rect 676870 440746 677040 440754
rect 676870 440712 677040 440746
rect 676870 440702 677040 440712
rect 677540 440530 677550 440748
rect 677550 440530 677584 440748
rect 677584 440530 677592 440748
rect 676928 440260 676938 440478
rect 676938 440260 676972 440478
rect 676972 440260 676980 440478
rect 677482 440196 677652 440204
rect 677482 440162 677652 440196
rect 677482 440152 677652 440162
rect 676870 439550 677040 439558
rect 676870 439516 677040 439550
rect 676870 439506 677040 439516
rect 677540 439334 677550 439552
rect 677550 439334 677584 439552
rect 677584 439334 677592 439552
<< metal2 >>
rect 417019 997567 417392 997584
rect 417019 997507 417027 997567
rect 417384 997507 417392 997567
rect 417019 997498 417392 997507
rect 664229 997485 664602 997502
rect 664229 997425 664237 997485
rect 664594 997425 664602 997485
rect 664229 997416 664602 997425
rect 168582 997238 168955 997255
rect 168582 997178 168590 997238
rect 168947 997178 168955 997238
rect 416856 997217 416862 997387
rect 416914 997217 416920 997387
rect 417514 997327 417732 997333
rect 417514 997269 417732 997275
rect 168582 997169 168955 997178
rect 167052 997002 167270 997008
rect 167052 996944 167270 996950
rect 167110 995183 167138 996944
rect 167864 996892 167870 997062
rect 167922 996892 167928 997062
rect 168248 997002 168466 997008
rect 168248 996944 168466 996950
rect 167218 996280 167224 996450
rect 167276 996280 167282 996450
rect 167234 995239 167262 996280
rect 167234 995233 167286 995239
rect 167110 995177 167162 995183
rect 167110 995119 167162 995125
rect 167234 995175 167286 995181
rect 167883 995179 167911 996892
rect 167978 996390 168196 996396
rect 167978 996332 168196 996338
rect 168077 995235 168105 996332
rect 168306 995295 168334 996944
rect 169060 996892 169066 997062
rect 169118 996892 169124 997062
rect 169444 997002 169662 997008
rect 169444 996944 169662 996950
rect 168414 996280 168420 996450
rect 168472 996280 168478 996450
rect 168430 995351 168458 996280
rect 168582 996156 168955 996170
rect 168582 996096 168590 996156
rect 168947 996096 168955 996156
rect 168582 996084 168955 996096
rect 168430 995345 168482 995351
rect 168306 995289 168358 995295
rect 168077 995229 168129 995235
rect 167110 995104 167138 995119
rect 167234 995104 167262 995175
rect 167883 995173 167935 995179
rect 167883 995115 167935 995121
rect 168077 995171 168129 995177
rect 168306 995231 168358 995237
rect 168430 995287 168482 995293
rect 169079 995291 169107 996892
rect 169174 996390 169392 996396
rect 169174 996332 169392 996338
rect 169273 995347 169301 996332
rect 169249 995341 169301 995347
rect 167883 995104 167911 995115
rect 168077 995104 168105 995171
rect 168306 995104 168334 995231
rect 168430 995104 168458 995287
rect 169079 995285 169131 995291
rect 169249 995283 169301 995289
rect 169079 995227 169131 995233
rect 169079 995104 169107 995227
rect 169273 995104 169301 995283
rect 169502 995407 169530 996944
rect 170256 996892 170262 997062
rect 170314 996892 170320 997062
rect 169778 996697 170151 996709
rect 169778 996637 169786 996697
rect 170143 996637 170151 996697
rect 169778 996623 170151 996637
rect 169610 996280 169616 996450
rect 169668 996280 169674 996450
rect 169626 995463 169654 996280
rect 169626 995457 169678 995463
rect 169502 995401 169554 995407
rect 169502 995343 169554 995349
rect 169626 995399 169678 995405
rect 170275 995403 170303 996892
rect 416588 996715 416806 996721
rect 416588 996657 416806 996663
rect 170370 996390 170588 996396
rect 170370 996332 170588 996338
rect 170469 995459 170497 996332
rect 170469 995453 170521 995459
rect 169502 995104 169530 995343
rect 169626 995104 169654 995399
rect 170275 995397 170327 995403
rect 170275 995339 170327 995345
rect 170469 995395 170521 995401
rect 170275 995104 170303 995339
rect 170469 995104 170497 995395
rect 416679 995277 416707 996657
rect 416655 995271 416707 995277
rect 416873 995221 416901 997217
rect 417502 996605 417508 996775
rect 417560 996605 417566 996775
rect 417019 996485 417392 996499
rect 417019 996425 417027 996485
rect 417384 996425 417392 996485
rect 417019 996413 417392 996425
rect 417522 995281 417550 996605
rect 416655 995213 416707 995219
rect 416679 995129 416707 995213
rect 416849 995215 416901 995221
rect 417498 995275 417550 995281
rect 417646 995225 417674 997269
rect 662857 997135 662863 997305
rect 662915 997135 662921 997305
rect 663515 997245 663733 997251
rect 663515 997187 663733 997193
rect 418215 997026 418588 997038
rect 418215 996966 418223 997026
rect 418580 996966 418588 997026
rect 418215 996952 418588 996966
rect 662589 996633 662807 996639
rect 662589 996575 662807 996581
rect 662680 995277 662708 996575
rect 417498 995217 417550 995223
rect 416849 995157 416901 995163
rect 416873 995129 416901 995157
rect 417522 995129 417550 995217
rect 417622 995219 417674 995225
rect 662656 995271 662708 995277
rect 662874 995221 662902 997135
rect 663503 996523 663509 996693
rect 663561 996523 663567 996693
rect 663523 995281 663551 996523
rect 662656 995213 662708 995219
rect 417622 995161 417674 995167
rect 417646 995129 417674 995161
rect 662680 994793 662708 995213
rect 662850 995215 662902 995221
rect 663499 995275 663551 995281
rect 663647 995225 663675 997187
rect 664053 997135 664059 997305
rect 664111 997135 664117 997305
rect 664711 997245 664929 997251
rect 664711 997187 664929 997193
rect 663785 996633 664003 996639
rect 663785 996575 664003 996581
rect 663499 995217 663551 995223
rect 662850 995157 662902 995163
rect 662874 994793 662902 995157
rect 663523 994793 663551 995217
rect 663623 995219 663675 995225
rect 663623 995161 663675 995167
rect 663876 995165 663904 996575
rect 663647 994793 663675 995161
rect 663852 995159 663904 995165
rect 664070 995109 664098 997135
rect 664699 996523 664705 996693
rect 664757 996523 664763 996693
rect 664229 996403 664602 996417
rect 664229 996343 664237 996403
rect 664594 996343 664602 996403
rect 664229 996331 664602 996343
rect 664719 995169 664747 996523
rect 663852 995101 663904 995107
rect 663876 994793 663904 995101
rect 664046 995103 664098 995109
rect 664695 995163 664747 995169
rect 664843 995113 664871 997187
rect 665249 997135 665255 997305
rect 665307 997135 665313 997305
rect 665907 997245 666125 997251
rect 665907 997187 666125 997193
rect 664981 996633 665199 996639
rect 664981 996575 665199 996581
rect 664695 995105 664747 995111
rect 664046 995045 664098 995051
rect 664070 994793 664098 995045
rect 664719 994793 664747 995105
rect 664819 995107 664871 995113
rect 664819 995049 664871 995055
rect 665072 995053 665100 996575
rect 664843 994793 664871 995049
rect 665048 995047 665100 995053
rect 665266 994997 665294 997135
rect 665425 996944 665798 996956
rect 665425 996884 665433 996944
rect 665790 996884 665798 996944
rect 665425 996870 665798 996884
rect 665895 996523 665901 996693
rect 665953 996523 665959 996693
rect 665915 995057 665943 996523
rect 665048 994989 665100 994995
rect 665072 994793 665100 994989
rect 665242 994991 665294 994997
rect 665891 995051 665943 995057
rect 666039 995001 666067 997187
rect 666445 997135 666451 997305
rect 666503 997135 666509 997305
rect 667103 997245 667321 997251
rect 667103 997187 667321 997193
rect 666177 996633 666395 996639
rect 666177 996575 666395 996581
rect 665891 994993 665943 994999
rect 665242 994933 665294 994939
rect 665266 994793 665294 994933
rect 665915 994793 665943 994993
rect 666015 994995 666067 995001
rect 666015 994937 666067 994943
rect 666268 994941 666296 996575
rect 666039 994793 666067 994937
rect 666244 994935 666296 994941
rect 666462 994885 666490 997135
rect 667091 996523 667097 996693
rect 667149 996523 667155 996693
rect 667111 994945 667139 996523
rect 666244 994877 666296 994883
rect 666268 994793 666296 994877
rect 666438 994879 666490 994885
rect 667087 994939 667139 994945
rect 667235 994889 667263 997187
rect 667087 994881 667139 994887
rect 666438 994821 666490 994827
rect 666462 994793 666490 994821
rect 667111 994793 667139 994881
rect 667211 994883 667263 994889
rect 667211 994825 667263 994831
rect 667235 994793 667263 994825
rect 40548 891200 40554 891418
rect 40606 891327 40612 891418
rect 42461 891327 42467 891351
rect 40606 891299 42467 891327
rect 42519 891327 42525 891351
rect 42519 891299 43035 891327
rect 40606 891200 40612 891299
rect 39882 891144 40052 891150
rect 42517 891133 42523 891157
rect 40052 891105 42523 891133
rect 42575 891133 42581 891157
rect 42575 891105 43035 891133
rect 39882 891086 40052 891092
rect 40494 890498 40664 890504
rect 39936 890274 39942 890492
rect 39994 890360 40000 890492
rect 42457 890484 42463 890508
rect 40664 890456 42463 890484
rect 42515 890484 42521 890508
rect 42515 890456 43035 890484
rect 40494 890440 40664 890446
rect 42513 890360 42519 890384
rect 39994 890332 42519 890360
rect 42571 890360 42577 890384
rect 42571 890332 43035 890360
rect 39994 890274 40000 890332
rect 40548 890004 40554 890222
rect 40606 890131 40612 890222
rect 40606 890103 42579 890131
rect 40606 890004 40612 890103
rect 42573 890079 42579 890103
rect 42631 890103 43035 890131
rect 42631 890079 42637 890103
rect 39882 889948 40052 889954
rect 42629 889937 42635 889961
rect 40052 889909 42635 889937
rect 42687 889937 42693 889961
rect 42687 889909 43035 889937
rect 39882 889890 40052 889896
rect 40229 889741 40315 889749
rect 40229 889384 40241 889741
rect 40301 889384 40315 889741
rect 40229 889376 40315 889384
rect 40494 889302 40664 889308
rect 39936 889078 39942 889296
rect 39994 889164 40000 889296
rect 42569 889288 42575 889312
rect 40664 889260 42575 889288
rect 42627 889288 42633 889312
rect 42627 889260 43035 889288
rect 40494 889244 40664 889250
rect 42625 889164 42631 889188
rect 39994 889136 42631 889164
rect 42683 889164 42689 889188
rect 42683 889136 43035 889164
rect 39994 889078 40000 889136
rect 40548 888808 40554 889026
rect 40606 888935 40612 889026
rect 42685 888935 42691 888959
rect 40606 888907 42691 888935
rect 42743 888935 42749 888959
rect 42743 888907 43035 888935
rect 40606 888808 40612 888907
rect 39882 888752 40052 888758
rect 42741 888741 42747 888765
rect 40052 888713 42747 888741
rect 42799 888741 42805 888765
rect 42799 888713 43035 888741
rect 39882 888694 40052 888700
rect 39683 888545 39769 888553
rect 39683 888188 39700 888545
rect 39760 888188 39769 888545
rect 39683 888180 39769 888188
rect 40768 888545 40854 888553
rect 40768 888188 40782 888545
rect 40842 888188 40854 888545
rect 40768 888180 40854 888188
rect 40494 888106 40664 888112
rect 39936 887882 39942 888100
rect 39994 887968 40000 888100
rect 42681 888092 42687 888116
rect 40664 888064 42687 888092
rect 42739 888092 42745 888116
rect 42739 888064 43035 888092
rect 40494 888048 40664 888054
rect 42737 887968 42743 887992
rect 39994 887940 42743 887968
rect 42795 887968 42801 887992
rect 42795 887940 43035 887968
rect 39994 887882 40000 887940
rect 40548 887612 40554 887830
rect 40606 887739 40612 887830
rect 40606 887711 42803 887739
rect 40606 887612 40612 887711
rect 42797 887687 42803 887711
rect 42855 887711 43035 887739
rect 42855 887687 42861 887711
rect 39882 887556 40052 887562
rect 42853 887545 42859 887569
rect 40052 887517 42859 887545
rect 42911 887545 42917 887569
rect 42911 887517 43035 887545
rect 39882 887498 40052 887504
rect 40494 886910 40664 886916
rect 39936 886686 39942 886904
rect 39994 886772 40000 886904
rect 42793 886896 42799 886920
rect 40664 886868 42799 886896
rect 42851 886896 42857 886920
rect 42851 886868 43035 886896
rect 40494 886852 40664 886858
rect 42849 886772 42855 886796
rect 39994 886744 42855 886772
rect 42907 886772 42913 886796
rect 42907 886744 43035 886772
rect 39994 886686 40000 886744
rect 40548 886416 40554 886634
rect 40606 886543 40612 886634
rect 42909 886543 42915 886567
rect 40606 886515 42915 886543
rect 42967 886543 42973 886567
rect 42967 886515 43035 886543
rect 40606 886416 40612 886515
rect 39882 886360 40052 886366
rect 42965 886349 42971 886373
rect 40052 886321 42971 886349
rect 43023 886349 43029 886373
rect 43023 886321 43035 886349
rect 39882 886302 40052 886308
rect 40494 885714 40664 885720
rect 39936 885490 39942 885708
rect 39994 885576 40000 885708
rect 42905 885700 42911 885724
rect 40664 885672 42911 885700
rect 42963 885700 42969 885724
rect 42963 885672 43035 885700
rect 40494 885656 40664 885662
rect 42961 885576 42967 885600
rect 39994 885548 42967 885576
rect 43019 885576 43025 885600
rect 43019 885548 43035 885576
rect 39994 885490 40000 885548
rect 676922 714367 676928 714458
rect 675018 714339 675092 714367
rect 675086 714315 675092 714339
rect 675144 714339 676928 714367
rect 675144 714315 675150 714339
rect 676922 714240 676928 714339
rect 676980 714240 676986 714458
rect 675030 714173 675036 714197
rect 675018 714145 675036 714173
rect 675088 714173 675094 714197
rect 677482 714184 677652 714190
rect 675088 714145 677482 714173
rect 677482 714126 677652 714132
rect 675090 713524 675096 713548
rect 675041 713496 675096 713524
rect 675148 713524 675154 713548
rect 676870 713538 677040 713544
rect 675148 713496 676870 713524
rect 676870 713480 677040 713486
rect 675034 713372 675040 713424
rect 675092 713400 675098 713424
rect 677534 713400 677540 713532
rect 675092 713372 677540 713400
rect 677534 713314 677540 713372
rect 677592 713314 677598 713532
rect 674974 713171 674980 713195
rect 674442 713143 674980 713171
rect 675032 713171 675038 713195
rect 676922 713171 676928 713262
rect 675032 713143 676928 713171
rect 676922 713044 676928 713143
rect 676980 713044 676986 713262
rect 674918 712977 674924 713001
rect 674442 712949 674924 712977
rect 674976 712977 674982 713001
rect 677482 712988 677652 712994
rect 674976 712949 677482 712977
rect 677482 712930 677652 712936
rect 674978 712328 674984 712352
rect 674442 712300 674984 712328
rect 675036 712328 675042 712352
rect 676870 712342 677040 712348
rect 675036 712300 676870 712328
rect 676870 712284 677040 712290
rect 674922 712204 674928 712228
rect 674442 712176 674928 712204
rect 674980 712204 674986 712228
rect 677534 712204 677540 712336
rect 674980 712176 677540 712204
rect 677534 712118 677540 712176
rect 677592 712118 677598 712336
rect 674862 711975 674868 711999
rect 674442 711947 674868 711975
rect 674920 711975 674926 711999
rect 676922 711975 676928 712066
rect 674920 711947 676928 711975
rect 676922 711848 676928 711947
rect 676980 711848 676986 712066
rect 674806 711781 674812 711805
rect 674442 711753 674812 711781
rect 674864 711781 674870 711805
rect 677482 711792 677652 711798
rect 674864 711753 677482 711781
rect 677482 711734 677652 711740
rect 676681 711653 676767 711661
rect 676681 711296 676693 711653
rect 676753 711296 676767 711653
rect 676681 711288 676767 711296
rect 677766 711653 677852 711661
rect 677766 711296 677775 711653
rect 677835 711296 677852 711653
rect 677766 711288 677852 711296
rect 674866 711132 674872 711156
rect 674442 711104 674872 711132
rect 674924 711132 674930 711156
rect 676870 711146 677040 711152
rect 674924 711104 676870 711132
rect 676870 711088 677040 711094
rect 674810 711008 674816 711032
rect 674442 710980 674816 711008
rect 674868 711008 674874 711032
rect 677534 711008 677540 711140
rect 674868 710980 677540 711008
rect 677534 710922 677540 710980
rect 677592 710922 677598 711140
rect 674750 710779 674756 710803
rect 674442 710751 674756 710779
rect 674808 710779 674814 710803
rect 676922 710779 676928 710870
rect 674808 710751 676928 710779
rect 676922 710652 676928 710751
rect 676980 710652 676986 710870
rect 674694 710585 674700 710609
rect 674442 710557 674700 710585
rect 674752 710585 674758 710609
rect 677482 710596 677652 710602
rect 674752 710557 677482 710585
rect 677482 710538 677652 710544
rect 677220 710457 677306 710465
rect 677220 710100 677234 710457
rect 677294 710100 677306 710457
rect 677220 710092 677306 710100
rect 674754 709936 674760 709960
rect 674442 709908 674760 709936
rect 674812 709936 674818 709960
rect 676870 709950 677040 709956
rect 674812 709908 676870 709936
rect 676870 709892 677040 709898
rect 674698 709812 674704 709836
rect 674442 709784 674704 709812
rect 674756 709812 674762 709836
rect 677534 709812 677540 709944
rect 674756 709784 677540 709812
rect 677534 709726 677540 709784
rect 677592 709726 677598 709944
rect 674638 709583 674644 709607
rect 674442 709555 674644 709583
rect 674696 709583 674702 709607
rect 676922 709583 676928 709674
rect 674696 709555 676928 709583
rect 676922 709456 676928 709555
rect 676980 709456 676986 709674
rect 674582 709389 674588 709413
rect 674442 709361 674588 709389
rect 674640 709389 674646 709413
rect 677482 709400 677652 709406
rect 674640 709361 677482 709389
rect 677482 709342 677652 709348
rect 674642 708740 674648 708764
rect 674442 708712 674648 708740
rect 674700 708740 674706 708764
rect 676870 708754 677040 708760
rect 674700 708712 676870 708740
rect 676870 708696 677040 708702
rect 674586 708616 674592 708640
rect 674442 708588 674592 708616
rect 674644 708616 674650 708640
rect 677534 708616 677540 708748
rect 674644 708588 677540 708616
rect 677534 708530 677540 708588
rect 677592 708530 677598 708748
rect 674526 708387 674532 708411
rect 674442 708359 674532 708387
rect 674584 708387 674590 708411
rect 676922 708387 676928 708478
rect 674584 708359 676928 708387
rect 676922 708260 676928 708359
rect 676980 708260 676986 708478
rect 674470 708193 674476 708217
rect 674442 708165 674476 708193
rect 674528 708193 674534 708217
rect 677482 708204 677652 708210
rect 674528 708165 677482 708193
rect 677482 708146 677652 708152
rect 674530 707544 674536 707568
rect 674442 707516 674536 707544
rect 674588 707544 674594 707568
rect 676870 707558 677040 707564
rect 674588 707516 676870 707544
rect 676870 707500 677040 707506
rect 674474 707420 674480 707444
rect 674442 707392 674480 707420
rect 674532 707420 674538 707444
rect 677534 707420 677540 707552
rect 674532 707392 677540 707420
rect 677534 707334 677540 707392
rect 677592 707334 677598 707552
rect 40573 610554 40579 610772
rect 40631 610681 40637 610772
rect 42433 610681 42439 610705
rect 40631 610653 42439 610681
rect 42491 610681 42497 610705
rect 42491 610653 43680 610681
rect 40631 610554 40637 610653
rect 39907 610498 40077 610504
rect 42489 610487 42495 610511
rect 40077 610459 42495 610487
rect 42547 610487 42553 610511
rect 42547 610459 43680 610487
rect 39907 610440 40077 610446
rect 40519 609852 40689 609858
rect 39961 609628 39967 609846
rect 40019 609714 40025 609846
rect 42429 609838 42435 609862
rect 40689 609810 42435 609838
rect 42487 609838 42493 609862
rect 42487 609810 43680 609838
rect 40519 609794 40689 609800
rect 42485 609714 42491 609738
rect 40019 609686 42491 609714
rect 42543 609714 42549 609738
rect 42543 609686 43680 609714
rect 40019 609628 40025 609686
rect 40573 609358 40579 609576
rect 40631 609485 40637 609576
rect 40631 609457 42551 609485
rect 40631 609358 40637 609457
rect 42545 609433 42551 609457
rect 42603 609457 43680 609485
rect 42603 609433 42609 609457
rect 39907 609302 40077 609308
rect 42601 609291 42607 609315
rect 40077 609263 42607 609291
rect 42659 609291 42665 609315
rect 42659 609263 43680 609291
rect 39907 609244 40077 609250
rect 40519 608656 40689 608662
rect 39961 608432 39967 608650
rect 40019 608518 40025 608650
rect 42541 608642 42547 608666
rect 40689 608614 42547 608642
rect 42599 608642 42605 608666
rect 42599 608614 43680 608642
rect 40519 608598 40689 608604
rect 42597 608518 42603 608542
rect 40019 608490 42603 608518
rect 42655 608518 42661 608542
rect 42655 608490 43680 608518
rect 40019 608432 40025 608490
rect 40573 608162 40579 608380
rect 40631 608289 40637 608380
rect 42657 608289 42663 608313
rect 40631 608261 42663 608289
rect 42715 608289 42721 608313
rect 42715 608261 43680 608289
rect 40631 608162 40637 608261
rect 39907 608106 40077 608112
rect 42713 608095 42719 608119
rect 40077 608067 42719 608095
rect 42771 608095 42777 608119
rect 42771 608067 43680 608095
rect 39907 608048 40077 608054
rect 40519 607460 40689 607466
rect 39961 607236 39967 607454
rect 40019 607322 40025 607454
rect 42653 607446 42659 607470
rect 40689 607418 42659 607446
rect 42711 607446 42717 607470
rect 42711 607418 43680 607446
rect 40519 607402 40689 607408
rect 42709 607322 42715 607346
rect 40019 607294 42715 607322
rect 42767 607322 42773 607346
rect 42767 607294 43680 607322
rect 40019 607236 40025 607294
rect 40573 606966 40579 607184
rect 40631 607093 40637 607184
rect 40631 607065 42775 607093
rect 40631 606966 40637 607065
rect 42769 607041 42775 607065
rect 42827 607065 43680 607093
rect 42827 607041 42833 607065
rect 39907 606910 40077 606916
rect 42825 606899 42831 606923
rect 40077 606871 42831 606899
rect 42883 606899 42889 606923
rect 42883 606871 43680 606899
rect 39907 606852 40077 606858
rect 40519 606264 40689 606270
rect 39961 606040 39967 606258
rect 40019 606126 40025 606258
rect 42765 606250 42771 606274
rect 40689 606222 42771 606250
rect 42823 606250 42829 606274
rect 42823 606222 43680 606250
rect 40519 606206 40689 606212
rect 42821 606126 42827 606150
rect 40019 606098 42827 606126
rect 42879 606126 42885 606150
rect 42879 606098 43680 606126
rect 40019 606040 40025 606098
rect 40573 605770 40579 605988
rect 40631 605897 40637 605988
rect 42881 605897 42887 605921
rect 40631 605869 42887 605897
rect 42939 605897 42945 605921
rect 42939 605869 43680 605897
rect 40631 605770 40637 605869
rect 39907 605714 40077 605720
rect 42937 605703 42943 605727
rect 40077 605675 42943 605703
rect 42995 605703 43001 605727
rect 42995 605675 43680 605703
rect 39907 605656 40077 605662
rect 40260 605567 40346 605575
rect 40260 605210 40272 605567
rect 40332 605210 40346 605567
rect 40260 605202 40346 605210
rect 40519 605068 40689 605074
rect 39961 604844 39967 605062
rect 40019 604930 40025 605062
rect 42877 605054 42883 605078
rect 40689 605026 42883 605054
rect 42935 605054 42941 605078
rect 42935 605026 43680 605054
rect 40519 605010 40689 605016
rect 42933 604930 42939 604954
rect 40019 604902 42939 604930
rect 42991 604930 42997 604954
rect 42991 604902 43680 604930
rect 40019 604844 40025 604902
rect 40573 604574 40579 604792
rect 40631 604701 40637 604792
rect 42993 604701 42999 604725
rect 40631 604673 42999 604701
rect 43051 604701 43057 604725
rect 43051 604673 43680 604701
rect 40631 604574 40637 604673
rect 39907 604518 40077 604524
rect 43049 604507 43055 604531
rect 40077 604479 43055 604507
rect 43107 604507 43113 604531
rect 43107 604479 43680 604507
rect 39907 604460 40077 604466
rect 39714 604371 39800 604379
rect 39714 604014 39731 604371
rect 39791 604014 39800 604371
rect 39714 604006 39800 604014
rect 40799 604371 40885 604379
rect 40799 604014 40813 604371
rect 40873 604014 40885 604371
rect 40799 604006 40885 604014
rect 40519 603872 40689 603878
rect 39961 603648 39967 603866
rect 40019 603734 40025 603866
rect 42989 603858 42995 603882
rect 40689 603830 42995 603858
rect 43047 603858 43053 603882
rect 43047 603830 43680 603858
rect 40519 603814 40689 603820
rect 43045 603734 43051 603758
rect 40019 603706 43051 603734
rect 43103 603734 43109 603758
rect 43103 603706 43680 603734
rect 40019 603648 40025 603706
rect 40573 603378 40579 603596
rect 40631 603505 40637 603596
rect 43105 603505 43111 603529
rect 40631 603477 43111 603505
rect 43163 603505 43169 603529
rect 43163 603477 43680 603505
rect 40631 603378 40637 603477
rect 39907 603322 40077 603328
rect 43161 603311 43167 603335
rect 40077 603283 43167 603311
rect 43219 603311 43225 603335
rect 43219 603283 43680 603311
rect 39907 603264 40077 603270
rect 40519 602676 40689 602682
rect 39961 602452 39967 602670
rect 40019 602538 40025 602670
rect 43101 602662 43107 602686
rect 40689 602634 43107 602662
rect 43159 602662 43165 602686
rect 43159 602634 43680 602662
rect 40519 602618 40689 602624
rect 43157 602538 43163 602562
rect 40019 602510 43163 602538
rect 43215 602538 43221 602562
rect 43215 602510 43680 602538
rect 40019 602452 40025 602510
rect 40573 602182 40579 602400
rect 40631 602309 40637 602400
rect 43217 602309 43223 602333
rect 40631 602281 43223 602309
rect 43275 602309 43281 602333
rect 43275 602281 43680 602309
rect 40631 602182 40637 602281
rect 39907 602126 40077 602132
rect 43273 602115 43279 602139
rect 40077 602087 43279 602115
rect 43331 602115 43337 602139
rect 43331 602087 43680 602115
rect 39907 602068 40077 602074
rect 40519 601480 40689 601486
rect 39961 601256 39967 601474
rect 40019 601342 40025 601474
rect 43213 601466 43219 601490
rect 40689 601438 43219 601466
rect 43271 601466 43277 601490
rect 43271 601438 43680 601466
rect 40519 601422 40689 601428
rect 43269 601342 43275 601366
rect 40019 601314 43275 601342
rect 43327 601342 43333 601366
rect 43327 601314 43680 601342
rect 40019 601256 40025 601314
rect 40573 600986 40579 601204
rect 40631 601113 40637 601204
rect 43329 601113 43335 601137
rect 40631 601085 43335 601113
rect 43387 601113 43393 601137
rect 43387 601085 43680 601113
rect 40631 600986 40637 601085
rect 39907 600930 40077 600936
rect 43385 600919 43391 600943
rect 40077 600891 43391 600919
rect 43443 600919 43449 600943
rect 43443 600891 43680 600919
rect 39907 600872 40077 600878
rect 40519 600284 40689 600290
rect 39961 600060 39967 600278
rect 40019 600146 40025 600278
rect 43325 600270 43331 600294
rect 40689 600242 43331 600270
rect 43383 600270 43389 600294
rect 43383 600242 43680 600270
rect 40519 600226 40689 600232
rect 43381 600146 43387 600170
rect 40019 600118 43387 600146
rect 43439 600146 43445 600170
rect 43439 600118 43680 600146
rect 40019 600060 40025 600118
rect 40573 599790 40579 600008
rect 40631 599917 40637 600008
rect 43441 599917 43447 599941
rect 40631 599889 43447 599917
rect 43499 599917 43505 599941
rect 43499 599889 43680 599917
rect 40631 599790 40637 599889
rect 39907 599734 40077 599740
rect 43497 599723 43503 599747
rect 40077 599695 43503 599723
rect 43555 599723 43561 599747
rect 43555 599695 43680 599723
rect 39907 599676 40077 599682
rect 40519 599088 40689 599094
rect 39961 598864 39967 599082
rect 40019 598950 40025 599082
rect 43437 599074 43443 599098
rect 40689 599046 43443 599074
rect 43495 599074 43501 599098
rect 43495 599046 43680 599074
rect 40519 599030 40689 599036
rect 43493 598950 43499 598974
rect 40019 598922 43499 598950
rect 43551 598950 43557 598974
rect 43551 598922 43680 598950
rect 40019 598864 40025 598922
rect 40573 598594 40579 598812
rect 40631 598721 40637 598812
rect 43553 598721 43559 598745
rect 40631 598693 43559 598721
rect 43611 598721 43617 598745
rect 43611 598693 43680 598721
rect 40631 598594 40637 598693
rect 39907 598538 40077 598544
rect 43609 598527 43615 598551
rect 40077 598499 43615 598527
rect 43667 598527 43673 598551
rect 43667 598499 43680 598527
rect 39907 598480 40077 598486
rect 40519 597892 40689 597898
rect 39961 597668 39967 597886
rect 40019 597754 40025 597886
rect 43549 597878 43555 597902
rect 40689 597850 43555 597878
rect 43607 597878 43613 597902
rect 43607 597850 43680 597878
rect 40519 597834 40689 597840
rect 43605 597754 43611 597778
rect 40019 597726 43611 597754
rect 43663 597754 43669 597778
rect 43663 597726 43680 597754
rect 40019 597668 40025 597726
rect 675086 453543 675092 453567
rect 673770 453515 675092 453543
rect 675144 453543 675150 453567
rect 676922 453543 676928 453634
rect 675144 453515 676928 453543
rect 676922 453416 676928 453515
rect 676980 453416 676986 453634
rect 675030 453349 675036 453373
rect 673770 453321 675036 453349
rect 675088 453349 675094 453373
rect 677482 453360 677652 453366
rect 675088 453321 677482 453349
rect 677482 453302 677652 453308
rect 675090 452700 675096 452724
rect 673770 452672 675096 452700
rect 675148 452700 675154 452724
rect 676870 452714 677040 452720
rect 675148 452672 676870 452700
rect 676870 452656 677040 452662
rect 675034 452576 675040 452600
rect 673770 452548 675040 452576
rect 675092 452576 675098 452600
rect 677534 452576 677540 452708
rect 675092 452548 677540 452576
rect 677534 452490 677540 452548
rect 677592 452490 677598 452708
rect 676922 452347 676928 452438
rect 673770 452319 674980 452347
rect 674974 452295 674980 452319
rect 675032 452319 676928 452347
rect 675032 452295 675038 452319
rect 676922 452220 676928 452319
rect 676980 452220 676986 452438
rect 674918 452153 674924 452177
rect 673770 452125 674924 452153
rect 674976 452153 674982 452177
rect 677482 452164 677652 452170
rect 674976 452125 677482 452153
rect 677482 452106 677652 452112
rect 674978 451504 674984 451528
rect 673770 451476 674984 451504
rect 675036 451504 675042 451528
rect 676870 451518 677040 451524
rect 675036 451476 676870 451504
rect 676870 451460 677040 451466
rect 674922 451380 674928 451404
rect 673770 451352 674928 451380
rect 674980 451380 674986 451404
rect 677534 451380 677540 451512
rect 674980 451352 677540 451380
rect 677534 451294 677540 451352
rect 677592 451294 677598 451512
rect 674862 451151 674868 451175
rect 673770 451123 674868 451151
rect 674920 451151 674926 451175
rect 676922 451151 676928 451242
rect 674920 451123 676928 451151
rect 676922 451024 676928 451123
rect 676980 451024 676986 451242
rect 674806 450957 674812 450981
rect 673770 450929 674812 450957
rect 674864 450957 674870 450981
rect 677482 450968 677652 450974
rect 674864 450929 677482 450957
rect 677482 450910 677652 450916
rect 674866 450308 674872 450332
rect 673770 450280 674872 450308
rect 674924 450308 674930 450332
rect 676870 450322 677040 450328
rect 674924 450280 676870 450308
rect 676870 450264 677040 450270
rect 674810 450184 674816 450208
rect 673770 450156 674816 450184
rect 674868 450184 674874 450208
rect 677534 450184 677540 450316
rect 674868 450156 677540 450184
rect 677534 450098 677540 450156
rect 677592 450098 677598 450316
rect 676922 449955 676928 450046
rect 673770 449927 674756 449955
rect 674750 449903 674756 449927
rect 674808 449927 676928 449955
rect 674808 449903 674814 449927
rect 676922 449828 676928 449927
rect 676980 449828 676986 450046
rect 674694 449761 674700 449785
rect 673770 449733 674700 449761
rect 674752 449761 674758 449785
rect 677482 449772 677652 449778
rect 674752 449733 677482 449761
rect 677482 449714 677652 449720
rect 674754 449112 674760 449136
rect 673770 449084 674760 449112
rect 674812 449112 674818 449136
rect 676870 449126 677040 449132
rect 674812 449084 676870 449112
rect 676870 449068 677040 449074
rect 674698 448988 674704 449012
rect 673770 448960 674704 448988
rect 674756 448988 674762 449012
rect 677534 448988 677540 449120
rect 674756 448960 677540 448988
rect 677534 448902 677540 448960
rect 677592 448902 677598 449120
rect 674638 448759 674644 448783
rect 673770 448731 674644 448759
rect 674696 448759 674702 448783
rect 676922 448759 676928 448850
rect 674696 448731 676928 448759
rect 676922 448632 676928 448731
rect 676980 448632 676986 448850
rect 674582 448565 674588 448589
rect 673770 448537 674588 448565
rect 674640 448565 674646 448589
rect 677482 448576 677652 448582
rect 674640 448537 677482 448565
rect 677482 448518 677652 448524
rect 676673 448452 676759 448460
rect 676673 448095 676685 448452
rect 676745 448095 676759 448452
rect 676673 448087 676759 448095
rect 677758 448452 677844 448460
rect 677758 448095 677767 448452
rect 677827 448095 677844 448452
rect 677758 448087 677844 448095
rect 674642 447916 674648 447940
rect 673770 447888 674648 447916
rect 674700 447916 674706 447940
rect 676870 447930 677040 447936
rect 674700 447888 676870 447916
rect 676870 447872 677040 447878
rect 674586 447792 674592 447816
rect 673770 447764 674592 447792
rect 674644 447792 674650 447816
rect 677534 447792 677540 447924
rect 674644 447764 677540 447792
rect 677534 447706 677540 447764
rect 677592 447706 677598 447924
rect 674526 447563 674532 447587
rect 673770 447535 674532 447563
rect 674584 447563 674590 447587
rect 676922 447563 676928 447654
rect 674584 447535 676928 447563
rect 676922 447436 676928 447535
rect 676980 447436 676986 447654
rect 674470 447369 674476 447393
rect 673770 447341 674476 447369
rect 674528 447369 674534 447393
rect 677482 447380 677652 447386
rect 674528 447341 677482 447369
rect 677482 447322 677652 447328
rect 677212 447256 677298 447264
rect 677212 446899 677226 447256
rect 677286 446899 677298 447256
rect 677212 446891 677298 446899
rect 674530 446720 674536 446744
rect 673770 446692 674536 446720
rect 674588 446720 674594 446744
rect 676870 446734 677040 446740
rect 674588 446692 676870 446720
rect 676870 446676 677040 446682
rect 674474 446596 674480 446620
rect 673770 446568 674480 446596
rect 674532 446596 674538 446620
rect 677534 446596 677540 446728
rect 674532 446568 677540 446596
rect 677534 446510 677540 446568
rect 677592 446510 677598 446728
rect 674414 446367 674420 446391
rect 673770 446339 674420 446367
rect 674472 446367 674478 446391
rect 676922 446367 676928 446458
rect 674472 446339 676928 446367
rect 676922 446240 676928 446339
rect 676980 446240 676986 446458
rect 674358 446173 674364 446197
rect 673770 446145 674364 446173
rect 674416 446173 674422 446197
rect 677482 446184 677652 446190
rect 674416 446145 677482 446173
rect 677482 446126 677652 446132
rect 674418 445524 674424 445548
rect 673770 445496 674424 445524
rect 674476 445524 674482 445548
rect 676870 445538 677040 445544
rect 674476 445496 676870 445524
rect 676870 445480 677040 445486
rect 674362 445400 674368 445424
rect 673770 445372 674368 445400
rect 674420 445400 674426 445424
rect 677534 445400 677540 445532
rect 674420 445372 677540 445400
rect 677534 445314 677540 445372
rect 677592 445314 677598 445532
rect 674302 445171 674308 445195
rect 673770 445143 674308 445171
rect 674360 445171 674366 445195
rect 676922 445171 676928 445262
rect 674360 445143 676928 445171
rect 676922 445044 676928 445143
rect 676980 445044 676986 445262
rect 674246 444977 674252 445001
rect 673770 444949 674252 444977
rect 674304 444977 674310 445001
rect 677482 444988 677652 444994
rect 674304 444949 677482 444977
rect 677482 444930 677652 444936
rect 674306 444328 674312 444352
rect 673770 444300 674312 444328
rect 674364 444328 674370 444352
rect 676870 444342 677040 444348
rect 674364 444300 676870 444328
rect 676870 444284 677040 444290
rect 674250 444204 674256 444228
rect 673770 444176 674256 444204
rect 674308 444204 674314 444228
rect 677534 444204 677540 444336
rect 674308 444176 677540 444204
rect 677534 444118 677540 444176
rect 677592 444118 677598 444336
rect 674190 443975 674196 443999
rect 673770 443947 674196 443975
rect 674248 443975 674254 443999
rect 676922 443975 676928 444066
rect 674248 443947 676928 443975
rect 676922 443848 676928 443947
rect 676980 443848 676986 444066
rect 674134 443781 674140 443805
rect 673770 443753 674140 443781
rect 674192 443781 674198 443805
rect 677482 443792 677652 443798
rect 674192 443753 677482 443781
rect 677482 443734 677652 443740
rect 674194 443132 674200 443156
rect 673770 443104 674200 443132
rect 674252 443132 674258 443156
rect 676870 443146 677040 443152
rect 674252 443104 676870 443132
rect 676870 443088 677040 443094
rect 674138 443008 674144 443032
rect 673770 442980 674144 443008
rect 674196 443008 674202 443032
rect 677534 443008 677540 443140
rect 674196 442980 677540 443008
rect 677534 442922 677540 442980
rect 677592 442922 677598 443140
rect 674078 442779 674084 442803
rect 673770 442751 674084 442779
rect 674136 442779 674142 442803
rect 676922 442779 676928 442870
rect 674136 442751 676928 442779
rect 676922 442652 676928 442751
rect 676980 442652 676986 442870
rect 674022 442585 674028 442609
rect 673770 442557 674028 442585
rect 674080 442585 674086 442609
rect 677482 442596 677652 442602
rect 674080 442557 677482 442585
rect 677482 442538 677652 442544
rect 674082 441936 674088 441960
rect 673770 441908 674088 441936
rect 674140 441936 674146 441960
rect 676870 441950 677040 441956
rect 674140 441908 676870 441936
rect 676870 441892 677040 441898
rect 674026 441812 674032 441836
rect 673770 441784 674032 441812
rect 674084 441812 674090 441836
rect 677534 441812 677540 441944
rect 674084 441784 677540 441812
rect 677534 441726 677540 441784
rect 677592 441726 677598 441944
rect 673966 441583 673972 441607
rect 673770 441555 673972 441583
rect 674024 441583 674030 441607
rect 676922 441583 676928 441674
rect 674024 441555 676928 441583
rect 676922 441456 676928 441555
rect 676980 441456 676986 441674
rect 673910 441389 673916 441413
rect 673770 441361 673916 441389
rect 673968 441389 673974 441413
rect 677482 441400 677652 441406
rect 673968 441361 677482 441389
rect 677482 441342 677652 441348
rect 673970 440740 673976 440764
rect 673770 440712 673976 440740
rect 674028 440740 674034 440764
rect 676870 440754 677040 440760
rect 674028 440712 676870 440740
rect 676870 440696 677040 440702
rect 673914 440616 673920 440640
rect 673770 440588 673920 440616
rect 673972 440616 673978 440640
rect 677534 440616 677540 440748
rect 673972 440588 677540 440616
rect 677534 440530 677540 440588
rect 677592 440530 677598 440748
rect 673854 440387 673860 440411
rect 673770 440359 673860 440387
rect 673912 440387 673918 440411
rect 676922 440387 676928 440478
rect 673912 440359 676928 440387
rect 676922 440260 676928 440359
rect 676980 440260 676986 440478
rect 673798 440193 673804 440217
rect 673770 440165 673804 440193
rect 673856 440193 673862 440217
rect 677482 440204 677652 440210
rect 673856 440165 677482 440193
rect 677482 440146 677652 440152
rect 673858 439544 673864 439568
rect 673770 439516 673864 439544
rect 673916 439544 673922 439568
rect 676870 439558 677040 439564
rect 673916 439516 676870 439544
rect 676870 439500 677040 439506
rect 673802 439420 673808 439444
rect 673770 439392 673808 439420
rect 673860 439420 673866 439444
rect 677534 439420 677540 439552
rect 673860 439392 677540 439420
rect 677534 439334 677540 439392
rect 677592 439334 677598 439552
rect 40595 352373 40601 352591
rect 40653 352500 40659 352591
rect 42405 352500 42411 352524
rect 40653 352472 42411 352500
rect 42463 352500 42469 352524
rect 42463 352472 44108 352500
rect 40653 352373 40659 352472
rect 39929 352317 40099 352323
rect 42461 352306 42467 352330
rect 40099 352278 42467 352306
rect 42519 352306 42525 352330
rect 42519 352278 44108 352306
rect 39929 352259 40099 352265
rect 40541 351671 40711 351677
rect 39983 351447 39989 351665
rect 40041 351533 40047 351665
rect 42401 351657 42407 351681
rect 40711 351629 42407 351657
rect 42459 351657 42465 351681
rect 42459 351629 44108 351657
rect 40541 351613 40711 351619
rect 42457 351533 42463 351557
rect 40041 351505 42463 351533
rect 42515 351533 42521 351557
rect 42515 351505 44108 351533
rect 40041 351447 40047 351505
rect 40595 351177 40601 351395
rect 40653 351304 40659 351395
rect 40653 351276 42523 351304
rect 40653 351177 40659 351276
rect 42517 351252 42523 351276
rect 42575 351276 44108 351304
rect 42575 351252 42581 351276
rect 39929 351121 40099 351127
rect 42573 351110 42579 351134
rect 40099 351082 42579 351110
rect 42631 351110 42637 351134
rect 42631 351082 44108 351110
rect 39929 351063 40099 351069
rect 40541 350475 40711 350481
rect 39983 350251 39989 350469
rect 40041 350337 40047 350469
rect 42513 350461 42519 350485
rect 40711 350433 42519 350461
rect 42571 350461 42577 350485
rect 42571 350433 44108 350461
rect 40541 350417 40711 350423
rect 42569 350337 42575 350361
rect 40041 350309 42575 350337
rect 42627 350337 42633 350361
rect 42627 350309 44108 350337
rect 40041 350251 40047 350309
rect 40595 349981 40601 350199
rect 40653 350108 40659 350199
rect 42629 350108 42635 350132
rect 40653 350080 42635 350108
rect 42687 350108 42693 350132
rect 42687 350080 44108 350108
rect 40653 349981 40659 350080
rect 39929 349925 40099 349931
rect 42685 349914 42691 349938
rect 40099 349886 42691 349914
rect 42743 349914 42749 349938
rect 42743 349886 44108 349914
rect 39929 349867 40099 349873
rect 40541 349279 40711 349285
rect 39983 349055 39989 349273
rect 40041 349141 40047 349273
rect 42625 349265 42631 349289
rect 40711 349237 42631 349265
rect 42683 349265 42689 349289
rect 42683 349237 44108 349265
rect 40541 349221 40711 349227
rect 42681 349141 42687 349165
rect 40041 349113 42687 349141
rect 42739 349141 42745 349165
rect 42739 349113 44108 349141
rect 40041 349055 40047 349113
rect 40595 348785 40601 349003
rect 40653 348912 40659 349003
rect 40653 348884 42747 348912
rect 40653 348785 40659 348884
rect 42741 348860 42747 348884
rect 42799 348884 44108 348912
rect 42799 348860 42805 348884
rect 39929 348729 40099 348735
rect 42797 348718 42803 348742
rect 40099 348690 42803 348718
rect 42855 348718 42861 348742
rect 42855 348690 44108 348718
rect 39929 348671 40099 348677
rect 40541 348083 40711 348089
rect 39983 347859 39989 348077
rect 40041 347945 40047 348077
rect 42737 348069 42743 348093
rect 40711 348041 42743 348069
rect 42795 348069 42801 348093
rect 42795 348041 44108 348069
rect 40541 348025 40711 348031
rect 42793 347945 42799 347969
rect 40041 347917 42799 347945
rect 42851 347945 42857 347969
rect 42851 347917 44108 347945
rect 40041 347859 40047 347917
rect 40595 347589 40601 347807
rect 40653 347716 40659 347807
rect 42853 347716 42859 347740
rect 40653 347688 42859 347716
rect 42911 347716 42917 347740
rect 42911 347688 44108 347716
rect 40653 347589 40659 347688
rect 39929 347533 40099 347539
rect 42909 347522 42915 347546
rect 40099 347494 42915 347522
rect 42967 347522 42973 347546
rect 42967 347494 44108 347522
rect 39929 347475 40099 347481
rect 40541 346887 40711 346893
rect 39983 346663 39989 346881
rect 40041 346749 40047 346881
rect 42849 346873 42855 346897
rect 40711 346845 42855 346873
rect 42907 346873 42913 346897
rect 42907 346845 44108 346873
rect 40541 346829 40711 346835
rect 42905 346749 42911 346773
rect 40041 346721 42911 346749
rect 42963 346749 42969 346773
rect 42963 346721 44108 346749
rect 40041 346663 40047 346721
rect 40595 346393 40601 346611
rect 40653 346520 40659 346611
rect 42965 346520 42971 346544
rect 40653 346492 42971 346520
rect 43023 346520 43029 346544
rect 43023 346492 44108 346520
rect 40653 346393 40659 346492
rect 39929 346337 40099 346343
rect 43021 346326 43027 346350
rect 40099 346298 43027 346326
rect 43079 346326 43085 346350
rect 43079 346298 44108 346326
rect 39929 346279 40099 346285
rect 40541 345691 40711 345697
rect 39983 345467 39989 345685
rect 40041 345553 40047 345685
rect 42961 345677 42967 345701
rect 40711 345649 42967 345677
rect 43019 345677 43025 345701
rect 43019 345649 44108 345677
rect 40541 345633 40711 345639
rect 43017 345553 43023 345577
rect 40041 345525 43023 345553
rect 43075 345553 43081 345577
rect 43075 345525 44108 345553
rect 40041 345467 40047 345525
rect 40595 345197 40601 345415
rect 40653 345324 40659 345415
rect 43077 345324 43083 345348
rect 40653 345296 43083 345324
rect 43135 345324 43141 345348
rect 43135 345296 44108 345324
rect 40653 345197 40659 345296
rect 39929 345141 40099 345147
rect 43133 345130 43139 345154
rect 40099 345102 43139 345130
rect 43191 345130 43197 345154
rect 43191 345102 44108 345130
rect 39929 345083 40099 345089
rect 40541 344495 40711 344501
rect 39983 344271 39989 344489
rect 40041 344357 40047 344489
rect 43073 344481 43079 344505
rect 40711 344453 43079 344481
rect 43131 344481 43137 344505
rect 43131 344453 44108 344481
rect 40541 344437 40711 344443
rect 43129 344357 43135 344381
rect 40041 344329 43135 344357
rect 43187 344357 43193 344381
rect 43187 344329 44108 344357
rect 40041 344271 40047 344329
rect 40595 344001 40601 344219
rect 40653 344128 40659 344219
rect 43189 344128 43195 344152
rect 40653 344100 43195 344128
rect 43247 344128 43253 344152
rect 43247 344100 44108 344128
rect 40653 344001 40659 344100
rect 39929 343945 40099 343951
rect 43245 343934 43251 343958
rect 40099 343906 43251 343934
rect 43303 343934 43309 343958
rect 43303 343906 44108 343934
rect 39929 343887 40099 343893
rect 40279 343728 40365 343736
rect 40279 343371 40291 343728
rect 40351 343371 40365 343728
rect 40279 343363 40365 343371
rect 40541 343299 40711 343305
rect 39983 343075 39989 343293
rect 40041 343161 40047 343293
rect 43185 343285 43191 343309
rect 40711 343257 43191 343285
rect 43243 343285 43249 343309
rect 43243 343257 44108 343285
rect 40541 343241 40711 343247
rect 43241 343161 43247 343185
rect 40041 343133 43247 343161
rect 43299 343161 43305 343185
rect 43299 343133 44108 343161
rect 40041 343075 40047 343133
rect 40595 342805 40601 343023
rect 40653 342932 40659 343023
rect 43301 342932 43307 342956
rect 40653 342904 43307 342932
rect 43359 342932 43365 342956
rect 43359 342904 44108 342932
rect 40653 342805 40659 342904
rect 39929 342749 40099 342755
rect 43357 342738 43363 342762
rect 40099 342710 43363 342738
rect 43415 342738 43421 342762
rect 43415 342710 44108 342738
rect 39929 342691 40099 342697
rect 39733 342532 39819 342540
rect 39733 342175 39750 342532
rect 39810 342175 39819 342532
rect 39733 342167 39819 342175
rect 40818 342532 40904 342540
rect 40818 342175 40832 342532
rect 40892 342175 40904 342532
rect 40818 342167 40904 342175
rect 40541 342103 40711 342109
rect 39983 341879 39989 342097
rect 40041 341965 40047 342097
rect 43297 342089 43303 342113
rect 40711 342061 43303 342089
rect 43355 342089 43361 342113
rect 43355 342061 44108 342089
rect 40541 342045 40711 342051
rect 43353 341965 43359 341989
rect 40041 341937 43359 341965
rect 43411 341965 43417 341989
rect 43411 341937 44108 341965
rect 40041 341879 40047 341937
rect 40595 341609 40601 341827
rect 40653 341736 40659 341827
rect 43413 341736 43419 341760
rect 40653 341708 43419 341736
rect 43471 341736 43477 341760
rect 43471 341708 44108 341736
rect 40653 341609 40659 341708
rect 39929 341553 40099 341559
rect 43469 341542 43475 341566
rect 40099 341514 43475 341542
rect 43527 341542 43533 341566
rect 43527 341514 44108 341542
rect 39929 341495 40099 341501
rect 40541 340907 40711 340913
rect 39983 340683 39989 340901
rect 40041 340769 40047 340901
rect 43409 340893 43415 340917
rect 40711 340865 43415 340893
rect 43467 340893 43473 340917
rect 43467 340865 44108 340893
rect 40541 340849 40711 340855
rect 43465 340769 43471 340793
rect 40041 340741 43471 340769
rect 43523 340769 43529 340793
rect 43523 340741 44108 340769
rect 40041 340683 40047 340741
rect 40595 340413 40601 340631
rect 40653 340540 40659 340631
rect 43525 340540 43531 340564
rect 40653 340512 43531 340540
rect 43583 340540 43589 340564
rect 43583 340512 44108 340540
rect 40653 340413 40659 340512
rect 39929 340357 40099 340363
rect 43581 340346 43587 340370
rect 40099 340318 43587 340346
rect 43639 340346 43645 340370
rect 43639 340318 44108 340346
rect 39929 340299 40099 340305
rect 40541 339711 40711 339717
rect 39983 339487 39989 339705
rect 40041 339573 40047 339705
rect 43521 339697 43527 339721
rect 40711 339669 43527 339697
rect 43579 339697 43585 339721
rect 43579 339669 44108 339697
rect 40541 339653 40711 339659
rect 43577 339573 43583 339597
rect 40041 339545 43583 339573
rect 43635 339573 43641 339597
rect 43635 339545 44108 339573
rect 40041 339487 40047 339545
rect 40595 339217 40601 339435
rect 40653 339344 40659 339435
rect 43637 339344 43643 339368
rect 40653 339316 43643 339344
rect 43695 339344 43701 339368
rect 43695 339316 44108 339344
rect 40653 339217 40659 339316
rect 39929 339161 40099 339167
rect 43693 339150 43699 339174
rect 40099 339122 43699 339150
rect 43751 339150 43757 339174
rect 43751 339122 44108 339150
rect 39929 339103 40099 339109
rect 40541 338515 40711 338521
rect 39983 338291 39989 338509
rect 40041 338377 40047 338509
rect 43633 338501 43639 338525
rect 40711 338473 43639 338501
rect 43691 338501 43697 338525
rect 43691 338473 44108 338501
rect 40541 338457 40711 338463
rect 43689 338377 43695 338401
rect 40041 338349 43695 338377
rect 43747 338377 43753 338401
rect 43747 338349 44108 338377
rect 40041 338291 40047 338349
rect 40595 338021 40601 338239
rect 40653 338148 40659 338239
rect 43749 338148 43755 338172
rect 40653 338120 43755 338148
rect 43807 338148 43813 338172
rect 43807 338120 44108 338148
rect 40653 338021 40659 338120
rect 39929 337965 40099 337971
rect 43805 337954 43811 337978
rect 40099 337926 43811 337954
rect 43863 337954 43869 337978
rect 43863 337926 44108 337954
rect 39929 337907 40099 337913
rect 40541 337319 40711 337325
rect 39983 337095 39989 337313
rect 40041 337181 40047 337313
rect 43745 337305 43751 337329
rect 40711 337277 43751 337305
rect 43803 337305 43809 337329
rect 43803 337277 44108 337305
rect 40541 337261 40711 337267
rect 43801 337181 43807 337205
rect 40041 337153 43807 337181
rect 43859 337181 43865 337205
rect 43859 337153 44108 337181
rect 40041 337095 40047 337153
rect 40595 336825 40601 337043
rect 40653 336952 40659 337043
rect 40653 336924 43867 336952
rect 40653 336825 40659 336924
rect 43861 336900 43867 336924
rect 43919 336924 44108 336952
rect 43919 336900 43925 336924
rect 39929 336769 40099 336775
rect 43917 336758 43923 336782
rect 40099 336730 43923 336758
rect 43975 336758 43981 336782
rect 43975 336730 44108 336758
rect 39929 336711 40099 336717
rect 40541 336123 40711 336129
rect 39983 335899 39989 336117
rect 40041 335985 40047 336117
rect 43857 336109 43863 336133
rect 40711 336081 43863 336109
rect 43915 336109 43921 336133
rect 43915 336081 44108 336109
rect 40541 336065 40711 336071
rect 43913 335985 43919 336009
rect 40041 335957 43919 335985
rect 43971 335985 43977 336009
rect 43971 335957 44108 335985
rect 40041 335899 40047 335957
rect 40595 335629 40601 335847
rect 40653 335756 40659 335847
rect 43973 335756 43979 335780
rect 40653 335728 43979 335756
rect 44031 335756 44037 335780
rect 44031 335728 44108 335756
rect 40653 335629 40659 335728
rect 39929 335573 40099 335579
rect 44029 335562 44035 335586
rect 40099 335534 44035 335562
rect 44087 335562 44093 335586
rect 44087 335534 44108 335562
rect 39929 335515 40099 335521
rect 40541 334927 40711 334933
rect 39983 334703 39989 334921
rect 40041 334789 40047 334921
rect 43969 334913 43975 334937
rect 40711 334885 43975 334913
rect 44027 334913 44033 334937
rect 44027 334885 44108 334913
rect 40541 334869 40711 334875
rect 44025 334789 44031 334813
rect 40041 334761 44031 334789
rect 44083 334789 44089 334813
rect 44083 334761 44108 334789
rect 40041 334703 40047 334761
rect 394104 225934 394132 225953
rect 394947 225938 394975 225953
rect 394104 225928 394156 225934
rect 134104 225906 134132 225925
rect 134947 225910 134975 225925
rect 134104 225900 134156 225906
rect 134104 225842 134156 225848
rect 134947 225904 134999 225910
rect 134947 225846 134999 225852
rect 135176 225850 135204 225925
rect 134104 223272 134132 225842
rect 134088 223102 134094 223272
rect 134146 223102 134152 223272
rect 134947 223220 134975 225846
rect 135176 225844 135228 225850
rect 135176 225786 135228 225792
rect 135300 225794 135328 225925
rect 135949 225854 135977 225925
rect 135949 225848 136001 225854
rect 135300 225788 135352 225794
rect 134848 223214 135066 223220
rect 134848 223156 135066 223162
rect 135176 222608 135204 225786
rect 135300 225730 135352 225736
rect 135949 225790 136001 225796
rect 136143 225798 136171 225925
rect 136143 225792 136195 225798
rect 135300 223272 135328 225730
rect 135284 223102 135290 223272
rect 135342 223102 135348 223272
rect 135949 222660 135977 225790
rect 136143 225734 136195 225740
rect 136372 225738 136400 225925
rect 136143 223220 136171 225734
rect 136372 225732 136424 225738
rect 136372 225674 136424 225680
rect 136496 225682 136524 225925
rect 137145 225742 137173 225925
rect 137145 225736 137197 225742
rect 136496 225676 136548 225682
rect 136044 223214 136262 223220
rect 136044 223156 136262 223162
rect 135118 222602 135336 222608
rect 135118 222544 135336 222550
rect 135930 222490 135936 222660
rect 135988 222490 135994 222660
rect 136372 222608 136400 225674
rect 136496 225618 136548 225624
rect 137145 225678 137197 225684
rect 137339 225686 137367 225925
rect 137339 225680 137391 225686
rect 136496 223272 136524 225618
rect 136480 223102 136486 223272
rect 136538 223102 136544 223272
rect 137145 222660 137173 225678
rect 137339 225622 137391 225628
rect 137568 225626 137596 225925
rect 137339 223220 137367 225622
rect 137568 225620 137620 225626
rect 137568 225562 137620 225568
rect 137692 225570 137720 225925
rect 138341 225630 138369 225925
rect 138341 225624 138393 225630
rect 137692 225564 137744 225570
rect 137240 223214 137458 223220
rect 137240 223156 137458 223162
rect 136314 222602 136532 222608
rect 136314 222544 136532 222550
rect 137126 222490 137132 222660
rect 137184 222490 137190 222660
rect 137568 222608 137596 225562
rect 137692 225506 137744 225512
rect 138341 225566 138393 225572
rect 138535 225574 138563 225925
rect 138535 225568 138587 225574
rect 137692 223272 137720 225506
rect 137676 223102 137682 223272
rect 137734 223102 137740 223272
rect 138341 222660 138369 225566
rect 138535 225510 138587 225516
rect 138764 225514 138792 225925
rect 138535 223220 138563 225510
rect 138764 225508 138816 225514
rect 138764 225450 138816 225456
rect 138888 225458 138916 225925
rect 139537 225518 139565 225925
rect 139537 225512 139589 225518
rect 138888 225452 138940 225458
rect 138436 223214 138654 223220
rect 138436 223156 138654 223162
rect 137510 222602 137728 222608
rect 137510 222544 137728 222550
rect 138322 222490 138328 222660
rect 138380 222490 138386 222660
rect 138764 222608 138792 225450
rect 138888 225394 138940 225400
rect 139537 225454 139589 225460
rect 139731 225462 139759 225925
rect 139731 225456 139783 225462
rect 138888 223272 138916 225394
rect 138872 223102 138878 223272
rect 138930 223102 138936 223272
rect 139537 222660 139565 225454
rect 139731 225398 139783 225404
rect 139960 225402 139988 225925
rect 139731 223220 139759 225398
rect 139960 225396 140012 225402
rect 139960 225338 140012 225344
rect 140084 225346 140112 225925
rect 140733 225406 140761 225925
rect 140733 225400 140785 225406
rect 140927 225350 140955 225925
rect 140084 225340 140136 225346
rect 139632 223214 139850 223220
rect 139632 223156 139850 223162
rect 138706 222602 138924 222608
rect 138706 222544 138924 222550
rect 139518 222490 139524 222660
rect 139576 222490 139582 222660
rect 139960 222608 139988 225338
rect 140084 225282 140136 225288
rect 140733 225342 140785 225348
rect 140903 225344 140955 225350
rect 140084 223272 140112 225282
rect 140068 223102 140074 223272
rect 140126 223102 140132 223272
rect 140733 222660 140761 225342
rect 140903 225286 140955 225292
rect 140927 223220 140955 225286
rect 141156 225290 141184 225925
rect 141156 225284 141208 225290
rect 141156 225226 141208 225232
rect 141280 225234 141308 225925
rect 141929 225294 141957 225925
rect 141929 225288 141981 225294
rect 141280 225228 141332 225234
rect 140828 223214 141046 223220
rect 140828 223156 141046 223162
rect 139902 222602 140120 222608
rect 139902 222544 140120 222550
rect 140714 222490 140720 222660
rect 140772 222490 140778 222660
rect 141156 222608 141184 225226
rect 141280 225170 141332 225176
rect 141929 225230 141981 225236
rect 142123 225238 142151 225925
rect 142123 225232 142175 225238
rect 141280 223272 141308 225170
rect 141264 223102 141270 223272
rect 141322 223102 141328 223272
rect 141929 222660 141957 225230
rect 142123 225174 142175 225180
rect 142352 225178 142380 225925
rect 142123 223220 142151 225174
rect 142352 225172 142404 225178
rect 142352 225114 142404 225120
rect 142476 225122 142504 225925
rect 143125 225182 143153 225925
rect 143125 225176 143177 225182
rect 143319 225126 143347 225925
rect 142476 225116 142528 225122
rect 142024 223214 142242 223220
rect 142024 223156 142242 223162
rect 141098 222602 141316 222608
rect 141098 222544 141316 222550
rect 141910 222490 141916 222660
rect 141968 222490 141974 222660
rect 142352 222608 142380 225114
rect 142476 225058 142528 225064
rect 143125 225118 143177 225124
rect 143295 225120 143347 225126
rect 142476 223272 142504 225058
rect 142460 223102 142466 223272
rect 142518 223102 142524 223272
rect 143125 222660 143153 225118
rect 143295 225062 143347 225068
rect 143319 223220 143347 225062
rect 143548 225066 143576 225925
rect 143548 225060 143600 225066
rect 143548 225002 143600 225008
rect 143672 225010 143700 225925
rect 144321 225070 144349 225925
rect 144321 225064 144373 225070
rect 143672 225004 143724 225010
rect 143220 223214 143438 223220
rect 143220 223156 143438 223162
rect 142294 222602 142512 222608
rect 142294 222544 142512 222550
rect 143106 222490 143112 222660
rect 143164 222490 143170 222660
rect 143548 222608 143576 225002
rect 143672 224946 143724 224952
rect 144321 225006 144373 225012
rect 144515 225014 144543 225925
rect 144515 225008 144567 225014
rect 143672 223272 143700 224946
rect 143656 223102 143662 223272
rect 143714 223102 143720 223272
rect 144321 222660 144349 225006
rect 144515 224950 144567 224956
rect 144744 224954 144772 225925
rect 144515 223220 144543 224950
rect 144744 224948 144796 224954
rect 144744 224890 144796 224896
rect 144868 224898 144896 225925
rect 145517 224958 145545 225925
rect 145517 224952 145569 224958
rect 144868 224892 144920 224898
rect 144416 223214 144634 223220
rect 144416 223156 144634 223162
rect 143490 222602 143708 222608
rect 143490 222544 143708 222550
rect 144302 222490 144308 222660
rect 144360 222490 144366 222660
rect 144744 222608 144772 224890
rect 144868 224834 144920 224840
rect 145517 224894 145569 224900
rect 145711 224902 145739 225925
rect 145711 224896 145763 224902
rect 144868 223272 144896 224834
rect 144852 223102 144858 223272
rect 144910 223102 144916 223272
rect 145517 222660 145545 224894
rect 145711 224838 145763 224844
rect 145940 224842 145968 225925
rect 145711 223220 145739 224838
rect 145940 224836 145992 224842
rect 145940 224778 145992 224784
rect 146064 224786 146092 225925
rect 146713 224846 146741 225925
rect 146713 224840 146765 224846
rect 146064 224780 146116 224786
rect 145612 223214 145830 223220
rect 145612 223156 145830 223162
rect 144686 222602 144904 222608
rect 144686 222544 144904 222550
rect 145498 222490 145504 222660
rect 145556 222490 145562 222660
rect 145940 222608 145968 224778
rect 146064 224722 146116 224728
rect 146713 224782 146765 224788
rect 146907 224790 146935 225925
rect 146907 224784 146959 224790
rect 146064 223272 146092 224722
rect 146048 223102 146054 223272
rect 146106 223102 146112 223272
rect 146191 222916 146564 222930
rect 146191 222856 146199 222916
rect 146556 222856 146564 222916
rect 146191 222844 146564 222856
rect 146713 222660 146741 224782
rect 146907 224726 146959 224732
rect 147136 224730 147164 225925
rect 146907 223220 146935 224726
rect 147136 224724 147188 224730
rect 147136 224666 147188 224672
rect 147260 224674 147288 225925
rect 147909 224734 147937 225925
rect 147909 224728 147961 224734
rect 147260 224668 147312 224674
rect 146808 223214 147026 223220
rect 146808 223156 147026 223162
rect 145882 222602 146100 222608
rect 145882 222544 146100 222550
rect 146694 222490 146700 222660
rect 146752 222490 146758 222660
rect 147136 222608 147164 224666
rect 147260 224610 147312 224616
rect 147909 224670 147961 224676
rect 148103 224678 148131 225925
rect 148103 224672 148155 224678
rect 147260 223272 147288 224610
rect 147387 223457 147760 223469
rect 147387 223397 147395 223457
rect 147752 223397 147760 223457
rect 147387 223383 147760 223397
rect 147244 223102 147250 223272
rect 147302 223102 147308 223272
rect 147909 222660 147937 224670
rect 148103 224614 148155 224620
rect 148332 224618 148360 225925
rect 148103 223220 148131 224614
rect 148332 224612 148384 224618
rect 148332 224554 148384 224560
rect 148456 224562 148484 225925
rect 149105 224622 149133 225925
rect 149105 224616 149157 224622
rect 148456 224556 148508 224562
rect 148004 223214 148222 223220
rect 148004 223156 148222 223162
rect 147078 222602 147296 222608
rect 147078 222544 147296 222550
rect 147890 222490 147896 222660
rect 147948 222490 147954 222660
rect 148332 222608 148360 224554
rect 148456 224498 148508 224504
rect 149105 224558 149157 224564
rect 149299 224566 149327 225925
rect 149299 224560 149351 224566
rect 148456 223272 148484 224498
rect 148440 223102 148446 223272
rect 148498 223102 148504 223272
rect 149105 222660 149133 224558
rect 149299 224502 149351 224508
rect 149528 224506 149556 225925
rect 149299 223220 149327 224502
rect 149528 224500 149580 224506
rect 149528 224442 149580 224448
rect 149652 224450 149680 225925
rect 150301 224510 150329 225925
rect 150301 224504 150353 224510
rect 149652 224444 149704 224450
rect 149200 223214 149418 223220
rect 149200 223156 149418 223162
rect 148274 222602 148492 222608
rect 148274 222544 148492 222550
rect 149086 222490 149092 222660
rect 149144 222490 149150 222660
rect 149528 222608 149556 224442
rect 149652 224386 149704 224392
rect 150301 224446 150353 224452
rect 150495 224454 150523 225925
rect 150495 224448 150547 224454
rect 149652 223272 149680 224386
rect 149636 223102 149642 223272
rect 149694 223102 149700 223272
rect 150301 222660 150329 224446
rect 150495 224390 150547 224396
rect 150724 224394 150752 225925
rect 150495 223220 150523 224390
rect 150724 224388 150776 224394
rect 150724 224330 150776 224336
rect 150848 224338 150876 225925
rect 151497 224398 151525 225925
rect 151497 224392 151549 224398
rect 150848 224332 150900 224338
rect 150396 223214 150614 223220
rect 150396 223156 150614 223162
rect 149470 222602 149688 222608
rect 149470 222544 149688 222550
rect 150282 222490 150288 222660
rect 150340 222490 150346 222660
rect 150724 222608 150752 224330
rect 150848 224274 150900 224280
rect 151497 224334 151549 224340
rect 151691 224342 151719 225925
rect 151691 224336 151743 224342
rect 150848 223272 150876 224274
rect 150832 223102 150838 223272
rect 150890 223102 150896 223272
rect 151497 222660 151525 224334
rect 151691 224278 151743 224284
rect 151920 224282 151948 225925
rect 151691 223220 151719 224278
rect 151920 224276 151972 224282
rect 151920 224218 151972 224224
rect 152044 224226 152072 225925
rect 152693 224286 152721 225925
rect 152693 224280 152745 224286
rect 152044 224220 152096 224226
rect 151592 223214 151810 223220
rect 151592 223156 151810 223162
rect 150666 222602 150884 222608
rect 150666 222544 150884 222550
rect 151478 222490 151484 222660
rect 151536 222490 151542 222660
rect 151920 222608 151948 224218
rect 152044 224162 152096 224168
rect 152693 224222 152745 224228
rect 152887 224230 152915 225925
rect 152887 224224 152939 224230
rect 152044 223272 152072 224162
rect 152028 223102 152034 223272
rect 152086 223102 152092 223272
rect 152693 222660 152721 224222
rect 152887 224166 152939 224172
rect 153116 224170 153144 225925
rect 152887 223220 152915 224166
rect 153116 224164 153168 224170
rect 153116 224106 153168 224112
rect 153240 224114 153268 225925
rect 153889 224174 153917 225925
rect 153889 224168 153941 224174
rect 153240 224108 153292 224114
rect 152788 223214 153006 223220
rect 152788 223156 153006 223162
rect 151862 222602 152080 222608
rect 151862 222544 152080 222550
rect 152674 222490 152680 222660
rect 152732 222490 152738 222660
rect 153116 222608 153144 224106
rect 153240 224050 153292 224056
rect 153889 224110 153941 224116
rect 154083 224118 154111 225925
rect 154083 224112 154135 224118
rect 153240 223272 153268 224050
rect 153224 223102 153230 223272
rect 153282 223102 153288 223272
rect 153889 222660 153917 224110
rect 154083 224054 154135 224060
rect 154312 224058 154340 225925
rect 154083 223220 154111 224054
rect 154312 224052 154364 224058
rect 154312 223994 154364 224000
rect 154436 224002 154464 225925
rect 155085 224062 155113 225925
rect 155085 224056 155137 224062
rect 155279 224006 155307 225925
rect 154436 223996 154488 224002
rect 153984 223214 154202 223220
rect 153984 223156 154202 223162
rect 153058 222602 153276 222608
rect 153058 222544 153276 222550
rect 153870 222490 153876 222660
rect 153928 222490 153934 222660
rect 154312 222608 154340 223994
rect 154436 223938 154488 223944
rect 155085 223998 155137 224004
rect 155255 224000 155307 224006
rect 154436 223272 154464 223938
rect 154420 223102 154426 223272
rect 154478 223102 154484 223272
rect 155085 222660 155113 223998
rect 155255 223942 155307 223948
rect 155279 223220 155307 223942
rect 155508 223946 155536 225925
rect 155508 223940 155560 223946
rect 155508 223882 155560 223888
rect 155632 223890 155660 225925
rect 156281 223950 156309 225925
rect 156281 223944 156333 223950
rect 155632 223884 155684 223890
rect 155180 223214 155398 223220
rect 155180 223156 155398 223162
rect 154254 222602 154472 222608
rect 154254 222544 154472 222550
rect 155066 222490 155072 222660
rect 155124 222490 155130 222660
rect 155508 222608 155536 223882
rect 155632 223826 155684 223832
rect 156281 223886 156333 223892
rect 156475 223894 156503 225925
rect 156475 223888 156527 223894
rect 155632 223272 155660 223826
rect 155616 223102 155622 223272
rect 155674 223102 155680 223272
rect 156281 222660 156309 223886
rect 156475 223830 156527 223836
rect 156704 223834 156732 225925
rect 156475 223220 156503 223830
rect 156704 223828 156756 223834
rect 156704 223770 156756 223776
rect 156828 223778 156856 225925
rect 157477 223838 157505 225925
rect 157477 223832 157529 223838
rect 157671 223782 157699 225925
rect 156828 223772 156880 223778
rect 156376 223214 156594 223220
rect 156376 223156 156594 223162
rect 155450 222602 155668 222608
rect 155450 222544 155668 222550
rect 156262 222490 156268 222660
rect 156320 222490 156326 222660
rect 156704 222608 156732 223770
rect 156828 223714 156880 223720
rect 157477 223774 157529 223780
rect 157647 223776 157699 223782
rect 156828 223272 156856 223714
rect 156812 223102 156818 223272
rect 156870 223102 156876 223272
rect 157477 222660 157505 223774
rect 157647 223718 157699 223724
rect 157671 223220 157699 223718
rect 157900 223722 157928 225925
rect 157900 223716 157952 223722
rect 157900 223658 157952 223664
rect 158024 223666 158052 225925
rect 158673 223726 158701 225925
rect 158673 223720 158725 223726
rect 158024 223660 158076 223666
rect 157572 223214 157790 223220
rect 157572 223156 157790 223162
rect 157900 222848 157928 223658
rect 158024 223602 158076 223608
rect 158673 223662 158725 223668
rect 158867 223670 158895 225925
rect 394104 225870 394156 225876
rect 394947 225932 394999 225938
rect 394947 225874 394999 225880
rect 395176 225878 395204 225953
rect 158867 223664 158919 223670
rect 158024 223272 158052 223602
rect 158008 223102 158014 223272
rect 158066 223102 158072 223272
rect 158673 222848 158701 223662
rect 158867 223606 158919 223612
rect 158867 223220 158895 223606
rect 394104 223272 394132 225870
rect 158768 223214 158986 223220
rect 158768 223156 158986 223162
rect 394088 223102 394094 223272
rect 394146 223102 394152 223272
rect 394947 223220 394975 225874
rect 395176 225872 395228 225878
rect 395176 225814 395228 225820
rect 395300 225822 395328 225953
rect 395949 225882 395977 225953
rect 395949 225876 396001 225882
rect 395300 225816 395352 225822
rect 394848 223214 395066 223220
rect 394848 223156 395066 223162
rect 157900 222820 158055 222848
rect 158673 222820 158828 222848
rect 158027 222660 158055 222820
rect 156646 222602 156864 222608
rect 156646 222544 156864 222550
rect 157458 222490 157464 222660
rect 157516 222490 157522 222660
rect 158010 222490 158016 222660
rect 158068 222490 158074 222660
rect 158800 222608 158828 222820
rect 395176 222608 395204 225814
rect 395300 225758 395352 225764
rect 395949 225818 396001 225824
rect 396143 225826 396171 225953
rect 396143 225820 396195 225826
rect 395300 223272 395328 225758
rect 395284 223102 395290 223272
rect 395342 223102 395348 223272
rect 395949 222660 395977 225818
rect 396143 225762 396195 225768
rect 396372 225766 396400 225953
rect 396143 223220 396171 225762
rect 396372 225760 396424 225766
rect 396372 225702 396424 225708
rect 396496 225710 396524 225953
rect 397145 225770 397173 225953
rect 397145 225764 397197 225770
rect 396496 225704 396548 225710
rect 396044 223214 396262 223220
rect 396044 223156 396262 223162
rect 158668 222602 158886 222608
rect 158668 222544 158886 222550
rect 395118 222602 395336 222608
rect 395118 222544 395336 222550
rect 395930 222490 395936 222660
rect 395988 222490 395994 222660
rect 396372 222608 396400 225702
rect 396496 225646 396548 225652
rect 397145 225706 397197 225712
rect 397339 225714 397367 225953
rect 397339 225708 397391 225714
rect 396496 223272 396524 225646
rect 396480 223102 396486 223272
rect 396538 223102 396544 223272
rect 397145 222660 397173 225706
rect 397339 225650 397391 225656
rect 397568 225654 397596 225953
rect 397339 223220 397367 225650
rect 397568 225648 397620 225654
rect 397568 225590 397620 225596
rect 397692 225598 397720 225953
rect 398341 225658 398369 225953
rect 398341 225652 398393 225658
rect 397692 225592 397744 225598
rect 397240 223214 397458 223220
rect 397240 223156 397458 223162
rect 396314 222602 396532 222608
rect 396314 222544 396532 222550
rect 397126 222490 397132 222660
rect 397184 222490 397190 222660
rect 397568 222608 397596 225590
rect 397692 225534 397744 225540
rect 398341 225594 398393 225600
rect 398535 225602 398563 225953
rect 398535 225596 398587 225602
rect 397692 223272 397720 225534
rect 397676 223102 397682 223272
rect 397734 223102 397740 223272
rect 398341 222660 398369 225594
rect 398535 225538 398587 225544
rect 398764 225542 398792 225953
rect 398535 223220 398563 225538
rect 398764 225536 398816 225542
rect 398764 225478 398816 225484
rect 398888 225486 398916 225953
rect 399537 225546 399565 225953
rect 399537 225540 399589 225546
rect 398888 225480 398940 225486
rect 398436 223214 398654 223220
rect 398436 223156 398654 223162
rect 397510 222602 397728 222608
rect 397510 222544 397728 222550
rect 398322 222490 398328 222660
rect 398380 222490 398386 222660
rect 398764 222608 398792 225478
rect 398888 225422 398940 225428
rect 399537 225482 399589 225488
rect 399731 225490 399759 225953
rect 399731 225484 399783 225490
rect 398888 223272 398916 225422
rect 398872 223102 398878 223272
rect 398930 223102 398936 223272
rect 399537 222660 399565 225482
rect 399731 225426 399783 225432
rect 399960 225430 399988 225953
rect 399731 223220 399759 225426
rect 399960 225424 400012 225430
rect 399960 225366 400012 225372
rect 400084 225374 400112 225953
rect 400733 225434 400761 225953
rect 400733 225428 400785 225434
rect 400927 225378 400955 225953
rect 400084 225368 400136 225374
rect 399632 223214 399850 223220
rect 399632 223156 399850 223162
rect 398706 222602 398924 222608
rect 398706 222544 398924 222550
rect 399518 222490 399524 222660
rect 399576 222490 399582 222660
rect 399960 222608 399988 225366
rect 400084 225310 400136 225316
rect 400733 225370 400785 225376
rect 400903 225372 400955 225378
rect 400084 223272 400112 225310
rect 400068 223102 400074 223272
rect 400126 223102 400132 223272
rect 400733 222660 400761 225370
rect 400903 225314 400955 225320
rect 400927 223220 400955 225314
rect 401156 225318 401184 225953
rect 401156 225312 401208 225318
rect 401156 225254 401208 225260
rect 401280 225262 401308 225953
rect 401929 225322 401957 225953
rect 401929 225316 401981 225322
rect 401280 225256 401332 225262
rect 400828 223214 401046 223220
rect 400828 223156 401046 223162
rect 399902 222602 400120 222608
rect 399902 222544 400120 222550
rect 400714 222490 400720 222660
rect 400772 222490 400778 222660
rect 401156 222608 401184 225254
rect 401280 225198 401332 225204
rect 401929 225258 401981 225264
rect 402123 225266 402151 225953
rect 402123 225260 402175 225266
rect 401280 223272 401308 225198
rect 401264 223102 401270 223272
rect 401322 223102 401328 223272
rect 401929 222660 401957 225258
rect 402123 225202 402175 225208
rect 402352 225206 402380 225953
rect 402123 223220 402151 225202
rect 402352 225200 402404 225206
rect 402352 225142 402404 225148
rect 402476 225150 402504 225953
rect 403125 225210 403153 225953
rect 403125 225204 403177 225210
rect 403319 225154 403347 225953
rect 402476 225144 402528 225150
rect 402024 223214 402242 223220
rect 402024 223156 402242 223162
rect 401098 222602 401316 222608
rect 401098 222544 401316 222550
rect 401910 222490 401916 222660
rect 401968 222490 401974 222660
rect 402352 222608 402380 225142
rect 402476 225086 402528 225092
rect 403125 225146 403177 225152
rect 403295 225148 403347 225154
rect 402476 223272 402504 225086
rect 402460 223102 402466 223272
rect 402518 223102 402524 223272
rect 403125 222660 403153 225146
rect 403295 225090 403347 225096
rect 403319 223220 403347 225090
rect 403548 225094 403576 225953
rect 403548 225088 403600 225094
rect 403548 225030 403600 225036
rect 403672 225038 403700 225953
rect 404321 225098 404349 225953
rect 404321 225092 404373 225098
rect 403672 225032 403724 225038
rect 403220 223214 403438 223220
rect 403220 223156 403438 223162
rect 402294 222602 402512 222608
rect 402294 222544 402512 222550
rect 403106 222490 403112 222660
rect 403164 222490 403170 222660
rect 403548 222608 403576 225030
rect 403672 224974 403724 224980
rect 404321 225034 404373 225040
rect 404515 225042 404543 225953
rect 404515 225036 404567 225042
rect 403672 223272 403700 224974
rect 403656 223102 403662 223272
rect 403714 223102 403720 223272
rect 404321 222660 404349 225034
rect 404515 224978 404567 224984
rect 404744 224982 404772 225953
rect 404515 223220 404543 224978
rect 404744 224976 404796 224982
rect 404744 224918 404796 224924
rect 404868 224926 404896 225953
rect 405517 224986 405545 225953
rect 405517 224980 405569 224986
rect 404868 224920 404920 224926
rect 404416 223214 404634 223220
rect 404416 223156 404634 223162
rect 403490 222602 403708 222608
rect 403490 222544 403708 222550
rect 404302 222490 404308 222660
rect 404360 222490 404366 222660
rect 404744 222608 404772 224918
rect 404868 224862 404920 224868
rect 405517 224922 405569 224928
rect 405711 224930 405739 225953
rect 405711 224924 405763 224930
rect 404868 223272 404896 224862
rect 404852 223102 404858 223272
rect 404910 223102 404916 223272
rect 405022 222909 405395 222923
rect 405022 222849 405030 222909
rect 405387 222849 405395 222909
rect 405022 222837 405395 222849
rect 405517 222660 405545 224922
rect 405711 224866 405763 224872
rect 405940 224870 405968 225953
rect 405711 223220 405739 224866
rect 405940 224864 405992 224870
rect 405940 224806 405992 224812
rect 406064 224814 406092 225953
rect 406713 224874 406741 225953
rect 406713 224868 406765 224874
rect 406064 224808 406116 224814
rect 405612 223214 405830 223220
rect 405612 223156 405830 223162
rect 404686 222602 404904 222608
rect 404686 222544 404904 222550
rect 405498 222490 405504 222660
rect 405556 222490 405562 222660
rect 405940 222608 405968 224806
rect 406064 224750 406116 224756
rect 406713 224810 406765 224816
rect 406907 224818 406935 225953
rect 406907 224812 406959 224818
rect 406064 223272 406092 224750
rect 406218 223450 406591 223462
rect 406218 223390 406226 223450
rect 406583 223390 406591 223450
rect 406218 223376 406591 223390
rect 406048 223102 406054 223272
rect 406106 223102 406112 223272
rect 406713 222660 406741 224810
rect 406907 224754 406959 224760
rect 407136 224758 407164 225953
rect 406907 223220 406935 224754
rect 407136 224752 407188 224758
rect 407136 224694 407188 224700
rect 407260 224702 407288 225953
rect 407909 224762 407937 225953
rect 407909 224756 407961 224762
rect 407260 224696 407312 224702
rect 406808 223214 407026 223220
rect 406808 223156 407026 223162
rect 405882 222602 406100 222608
rect 405882 222544 406100 222550
rect 406694 222490 406700 222660
rect 406752 222490 406758 222660
rect 407136 222608 407164 224694
rect 407260 224638 407312 224644
rect 407909 224698 407961 224704
rect 408103 224706 408131 225953
rect 408103 224700 408155 224706
rect 407260 223272 407288 224638
rect 407244 223102 407250 223272
rect 407302 223102 407308 223272
rect 407909 222660 407937 224698
rect 408103 224642 408155 224648
rect 408332 224646 408360 225953
rect 408103 223220 408131 224642
rect 408332 224640 408384 224646
rect 408332 224582 408384 224588
rect 408456 224590 408484 225953
rect 409105 224650 409133 225953
rect 409105 224644 409157 224650
rect 408456 224584 408508 224590
rect 408004 223214 408222 223220
rect 408004 223156 408222 223162
rect 407078 222602 407296 222608
rect 407078 222544 407296 222550
rect 407890 222490 407896 222660
rect 407948 222490 407954 222660
rect 408332 222608 408360 224582
rect 408456 224526 408508 224532
rect 409105 224586 409157 224592
rect 409299 224594 409327 225953
rect 409299 224588 409351 224594
rect 408456 223272 408484 224526
rect 408440 223102 408446 223272
rect 408498 223102 408504 223272
rect 409105 222660 409133 224586
rect 409299 224530 409351 224536
rect 409528 224534 409556 225953
rect 409299 223220 409327 224530
rect 409528 224528 409580 224534
rect 409528 224470 409580 224476
rect 409652 224478 409680 225953
rect 410301 224538 410329 225953
rect 410301 224532 410353 224538
rect 409652 224472 409704 224478
rect 409200 223214 409418 223220
rect 409200 223156 409418 223162
rect 408274 222602 408492 222608
rect 408274 222544 408492 222550
rect 409086 222490 409092 222660
rect 409144 222490 409150 222660
rect 409528 222608 409556 224470
rect 409652 224414 409704 224420
rect 410301 224474 410353 224480
rect 410495 224482 410523 225953
rect 410495 224476 410547 224482
rect 409652 223272 409680 224414
rect 409636 223102 409642 223272
rect 409694 223102 409700 223272
rect 410301 222660 410329 224474
rect 410495 224418 410547 224424
rect 410724 224422 410752 225953
rect 410495 223220 410523 224418
rect 410724 224416 410776 224422
rect 410724 224358 410776 224364
rect 410848 224366 410876 225953
rect 411497 224426 411525 225953
rect 411497 224420 411549 224426
rect 410848 224360 410900 224366
rect 410396 223214 410614 223220
rect 410396 223156 410614 223162
rect 409470 222602 409688 222608
rect 409470 222544 409688 222550
rect 410282 222490 410288 222660
rect 410340 222490 410346 222660
rect 410724 222608 410752 224358
rect 410848 224302 410900 224308
rect 411497 224362 411549 224368
rect 411691 224370 411719 225953
rect 411691 224364 411743 224370
rect 410848 223272 410876 224302
rect 410832 223102 410838 223272
rect 410890 223102 410896 223272
rect 411497 222660 411525 224362
rect 411691 224306 411743 224312
rect 411920 224310 411948 225953
rect 411691 223220 411719 224306
rect 411920 224304 411972 224310
rect 411920 224246 411972 224252
rect 412044 224254 412072 225953
rect 412693 224314 412721 225953
rect 412693 224308 412745 224314
rect 412044 224248 412096 224254
rect 411592 223214 411810 223220
rect 411592 223156 411810 223162
rect 410666 222602 410884 222608
rect 410666 222544 410884 222550
rect 411478 222490 411484 222660
rect 411536 222490 411542 222660
rect 411920 222608 411948 224246
rect 412044 224190 412096 224196
rect 412693 224250 412745 224256
rect 412887 224258 412915 225953
rect 412887 224252 412939 224258
rect 412044 223272 412072 224190
rect 412028 223102 412034 223272
rect 412086 223102 412092 223272
rect 412693 222660 412721 224250
rect 412887 224194 412939 224200
rect 413116 224198 413144 225953
rect 412887 223220 412915 224194
rect 413116 224192 413168 224198
rect 413116 224134 413168 224140
rect 413240 224142 413268 225953
rect 413889 224202 413917 225953
rect 413889 224196 413941 224202
rect 413240 224136 413292 224142
rect 412788 223214 413006 223220
rect 412788 223156 413006 223162
rect 411862 222602 412080 222608
rect 411862 222544 412080 222550
rect 412674 222490 412680 222660
rect 412732 222490 412738 222660
rect 413116 222608 413144 224134
rect 413240 224078 413292 224084
rect 413889 224138 413941 224144
rect 414083 224146 414111 225953
rect 414083 224140 414135 224146
rect 413240 223272 413268 224078
rect 413224 223102 413230 223272
rect 413282 223102 413288 223272
rect 413889 222660 413917 224138
rect 414083 224082 414135 224088
rect 414312 224086 414340 225953
rect 414083 223220 414111 224082
rect 414312 224080 414364 224086
rect 414312 224022 414364 224028
rect 414436 224030 414464 225953
rect 415085 224090 415113 225953
rect 415085 224084 415137 224090
rect 415279 224034 415307 225953
rect 414436 224024 414488 224030
rect 413984 223214 414202 223220
rect 413984 223156 414202 223162
rect 413058 222602 413276 222608
rect 413058 222544 413276 222550
rect 413870 222490 413876 222660
rect 413928 222490 413934 222660
rect 414312 222608 414340 224022
rect 414436 223966 414488 223972
rect 415085 224026 415137 224032
rect 415255 224028 415307 224034
rect 414436 223272 414464 223966
rect 414420 223102 414426 223272
rect 414478 223102 414484 223272
rect 415085 222660 415113 224026
rect 415255 223970 415307 223976
rect 415279 223220 415307 223970
rect 415508 223974 415536 225953
rect 415508 223968 415560 223974
rect 415508 223910 415560 223916
rect 415632 223918 415660 225953
rect 416281 223978 416309 225953
rect 416281 223972 416333 223978
rect 415632 223912 415684 223918
rect 415180 223214 415398 223220
rect 415180 223156 415398 223162
rect 414254 222602 414472 222608
rect 414254 222544 414472 222550
rect 415066 222490 415072 222660
rect 415124 222490 415130 222660
rect 415508 222608 415536 223910
rect 415632 223854 415684 223860
rect 416281 223914 416333 223920
rect 416475 223922 416503 225953
rect 416475 223916 416527 223922
rect 415632 223272 415660 223854
rect 415616 223102 415622 223272
rect 415674 223102 415680 223272
rect 416281 222660 416309 223914
rect 416475 223858 416527 223864
rect 416704 223862 416732 225953
rect 416475 223220 416503 223858
rect 416704 223856 416756 223862
rect 416704 223798 416756 223804
rect 416828 223806 416856 225953
rect 417477 223866 417505 225953
rect 417477 223860 417529 223866
rect 417671 223810 417699 225953
rect 416828 223800 416880 223806
rect 416376 223214 416594 223220
rect 416376 223156 416594 223162
rect 415450 222602 415668 222608
rect 415450 222544 415668 222550
rect 416262 222490 416268 222660
rect 416320 222490 416326 222660
rect 416704 222608 416732 223798
rect 416828 223742 416880 223748
rect 417477 223802 417529 223808
rect 417647 223804 417699 223810
rect 416828 223272 416856 223742
rect 416812 223102 416818 223272
rect 416870 223102 416876 223272
rect 417477 222660 417505 223802
rect 417647 223746 417699 223752
rect 417671 223220 417699 223746
rect 417900 223750 417928 225953
rect 417900 223744 417952 223750
rect 417900 223686 417952 223692
rect 418024 223694 418052 225953
rect 418673 223754 418701 225953
rect 418673 223748 418725 223754
rect 418024 223688 418076 223694
rect 417572 223214 417790 223220
rect 417572 223156 417790 223162
rect 417900 222834 417928 223686
rect 418024 223630 418076 223636
rect 418673 223690 418725 223696
rect 418867 223698 418895 225953
rect 418867 223692 418919 223698
rect 418024 223272 418052 223630
rect 418008 223102 418014 223272
rect 418066 223102 418072 223272
rect 418673 222834 418701 223690
rect 418867 223634 418919 223640
rect 418867 223220 418895 223634
rect 418768 223214 418986 223220
rect 418768 223156 418986 223162
rect 417900 222806 418055 222834
rect 418673 222806 418828 222834
rect 418027 222660 418055 222806
rect 416646 222602 416864 222608
rect 416646 222544 416864 222550
rect 417458 222490 417464 222660
rect 417516 222490 417522 222660
rect 418010 222490 418016 222660
rect 418068 222490 418074 222660
rect 418800 222608 418828 222806
rect 418668 222602 418886 222608
rect 418668 222544 418886 222550
rect 147387 222375 147760 222384
rect 147387 222315 147395 222375
rect 147752 222315 147760 222375
rect 147387 222298 147760 222315
rect 406218 222368 406591 222377
rect 406218 222308 406226 222368
rect 406583 222308 406591 222368
rect 406218 222291 406591 222308
<< via2 >>
rect 417027 997507 417384 997567
rect 664237 997425 664594 997485
rect 168590 997178 168947 997238
rect 168590 996096 168947 996156
rect 169786 996637 170143 996697
rect 417027 996425 417384 996485
rect 418223 996966 418580 997026
rect 664237 996343 664594 996403
rect 665433 996884 665790 996944
rect 40241 889384 40301 889741
rect 39700 888188 39760 888545
rect 40782 888188 40842 888545
rect 676693 711296 676753 711653
rect 677775 711296 677835 711653
rect 677234 710100 677294 710457
rect 40272 605210 40332 605567
rect 39731 604014 39791 604371
rect 40813 604014 40873 604371
rect 676685 448095 676745 448452
rect 677767 448095 677827 448452
rect 677226 446899 677286 447256
rect 40291 343371 40351 343728
rect 39750 342175 39810 342532
rect 40832 342175 40892 342532
rect 146199 222856 146556 222916
rect 147395 223397 147752 223457
rect 405030 222849 405387 222909
rect 406226 223390 406583 223450
rect 147395 222315 147752 222375
rect 406226 222308 406583 222368
<< metal3 >>
rect 168581 997238 168954 997586
rect 168581 997178 168590 997238
rect 168947 997178 168954 997238
rect 168581 996156 168954 997178
rect 169779 996697 170149 997586
rect 169779 996637 169786 996697
rect 170143 996637 170149 996697
rect 169779 996623 170149 996637
rect 417018 997567 417391 997915
rect 417018 997507 417027 997567
rect 417384 997507 417391 997567
rect 417018 996485 417391 997507
rect 418216 997026 418586 997915
rect 418216 996966 418223 997026
rect 418580 996966 418586 997026
rect 418216 996952 418586 996966
rect 664228 997485 664601 997833
rect 664228 997425 664237 997485
rect 664594 997425 664601 997485
rect 417018 996425 417027 996485
rect 417384 996425 417391 996485
rect 417018 996410 417391 996425
rect 664228 996403 664601 997425
rect 665426 996944 665796 997833
rect 665426 996884 665433 996944
rect 665790 996884 665796 996944
rect 665426 996870 665796 996884
rect 664228 996343 664237 996403
rect 664594 996343 664601 996403
rect 664228 996328 664601 996343
rect 168581 996096 168590 996156
rect 168947 996096 168954 996156
rect 168581 996081 168954 996096
rect 39352 889741 40315 889747
rect 39352 889384 40241 889741
rect 40301 889384 40315 889741
rect 39352 889377 40315 889384
rect 39352 888545 40857 888552
rect 39352 888188 39700 888545
rect 39760 888188 40782 888545
rect 40842 888188 40857 888545
rect 39352 888179 40857 888188
rect 676678 711653 678183 711662
rect 676678 711296 676693 711653
rect 676753 711296 677775 711653
rect 677835 711296 678183 711653
rect 676678 711289 678183 711296
rect 677220 710457 678183 710464
rect 677220 710100 677234 710457
rect 677294 710100 678183 710457
rect 677220 710094 678183 710100
rect 39383 605567 40346 605573
rect 39383 605210 40272 605567
rect 40332 605210 40346 605567
rect 39383 605203 40346 605210
rect 39383 604371 40888 604378
rect 39383 604014 39731 604371
rect 39791 604014 40813 604371
rect 40873 604014 40888 604371
rect 39383 604005 40888 604014
rect 676670 448452 678175 448461
rect 676670 448095 676685 448452
rect 676745 448095 677767 448452
rect 677827 448095 678175 448452
rect 676670 448088 678175 448095
rect 677212 447256 678175 447263
rect 677212 446899 677226 447256
rect 677286 446899 678175 447256
rect 677212 446893 678175 446899
rect 39402 343728 40365 343734
rect 39402 343371 40291 343728
rect 40351 343371 40365 343728
rect 39402 343364 40365 343371
rect 39402 342532 40907 342539
rect 39402 342175 39750 342532
rect 39810 342175 40832 342532
rect 40892 342175 40907 342532
rect 39402 342166 40907 342175
rect 147388 223457 147761 223472
rect 147388 223397 147395 223457
rect 147752 223397 147761 223457
rect 146193 222916 146563 222930
rect 146193 222856 146199 222916
rect 146556 222856 146563 222916
rect 146193 221967 146563 222856
rect 147388 222375 147761 223397
rect 406219 223450 406592 223465
rect 406219 223390 406226 223450
rect 406583 223390 406592 223450
rect 147388 222315 147395 222375
rect 147752 222315 147761 222375
rect 147388 221967 147761 222315
rect 405024 222909 405394 222923
rect 405024 222849 405030 222909
rect 405387 222849 405394 222909
rect 405024 221960 405394 222849
rect 406219 222368 406592 223390
rect 406219 222308 406226 222368
rect 406583 222308 406592 222368
rect 406219 221960 406592 222308
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 134996 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_2
timestamp 1663859327
transform 1 0 153028 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_3
timestamp 1663859327
transform -1 0 154132 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_4
timestamp 1663859327
transform 1 0 155420 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_5
timestamp 1663859327
transform -1 0 156524 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_6
timestamp 1663859327
transform 1 0 156616 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_7
timestamp 1663859327
transform -1 0 157720 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_8
timestamp 1663859327
transform -1 0 158916 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_9
timestamp 1663859327
transform -1 0 158916 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_10
timestamp 1663859327
transform -1 0 417762 0 -1 997540
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_11
timestamp 1663859327
transform 1 0 416658 0 1 996452
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_12
timestamp 1663859327
transform 0 -1 677805 1 0 439304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_13
timestamp 1663859327
transform 0 1 676717 -1 0 440408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_14
timestamp 1663859327
transform 0 1 676717 -1 0 448780
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_15
timestamp 1663859327
transform 0 -1 677805 1 0 447676
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_16
timestamp 1663859327
transform 0 1 676717 -1 0 452368
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_17
timestamp 1663859327
transform 0 -1 677805 1 0 451264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_18
timestamp 1663859327
transform 0 1 676717 -1 0 449976
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_19
timestamp 1663859327
transform 0 -1 677805 1 0 448872
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_20
timestamp 1663859327
transform 0 1 676717 -1 0 451172
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_21
timestamp 1663859327
transform 0 -1 677805 1 0 450068
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_22
timestamp 1663859327
transform 0 1 676717 -1 0 453564
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_23
timestamp 1663859327
transform 0 -1 677805 1 0 452460
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_24
timestamp 1663859327
transform 0 -1 677805 1 0 707304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_25
timestamp 1663859327
transform 0 1 676717 -1 0 708408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_26
timestamp 1663859327
transform 0 1 676717 -1 0 709604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_27
timestamp 1663859327
transform 0 -1 677805 1 0 708500
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_28
timestamp 1663859327
transform 0 1 676717 -1 0 710800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_29
timestamp 1663859327
transform 0 -1 677805 1 0 709696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_30
timestamp 1663859327
transform 0 1 676717 -1 0 711996
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_31
timestamp 1663859327
transform 0 -1 677805 1 0 710892
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_32
timestamp 1663859327
transform 0 1 676717 -1 0 714388
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_33
timestamp 1663859327
transform 0 -1 677805 1 0 713284
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_34
timestamp 1663859327
transform 0 1 676717 -1 0 446388
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_35
timestamp 1663859327
transform 0 -1 677805 1 0 445284
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_36
timestamp 1663859327
transform 0 1 676717 -1 0 447584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_37
timestamp 1663859327
transform 0 -1 677805 1 0 446480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_38
timestamp 1663859327
transform -1 0 169322 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_39
timestamp 1663859327
transform -1 0 168126 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_40
timestamp 1663859327
transform 0 -1 677805 1 0 712088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_41
timestamp 1663859327
transform 0 1 676717 -1 0 713192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_42
timestamp 1663859327
transform -1 0 170518 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_43
timestamp 1663859327
transform 1 0 169414 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_44
timestamp 1663859327
transform 1 0 168218 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_45
timestamp 1663859327
transform 1 0 167022 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_46
timestamp 1663859327
transform 0 1 676717 -1 0 441604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_47
timestamp 1663859327
transform 0 -1 677805 1 0 440500
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_48
timestamp 1663859327
transform 0 -1 677805 1 0 441696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_49
timestamp 1663859327
transform 0 1 676717 -1 0 442800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_50
timestamp 1663859327
transform 0 -1 677805 1 0 442892
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_51
timestamp 1663859327
transform 0 1 676717 -1 0 443996
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_52
timestamp 1663859327
transform 0 -1 677805 1 0 444088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_53
timestamp 1663859327
transform 0 1 676717 -1 0 445192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_54
timestamp 1663859327
transform 1 0 151832 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_55
timestamp 1663859327
transform -1 0 152936 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_56
timestamp 1663859327
transform 1 0 150636 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_57
timestamp 1663859327
transform -1 0 151740 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_58
timestamp 1663859327
transform 1 0 149440 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_59
timestamp 1663859327
transform -1 0 150544 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_60
timestamp 1663859327
transform 1 0 148244 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_61
timestamp 1663859327
transform -1 0 149348 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_62
timestamp 1663859327
transform 1 0 147048 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_63
timestamp 1663859327
transform -1 0 148152 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_64
timestamp 1663859327
transform 1 0 145852 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_65
timestamp 1663859327
transform -1 0 146956 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_66
timestamp 1663859327
transform -1 0 145760 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_67
timestamp 1663859327
transform 1 0 144656 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_68
timestamp 1663859327
transform 1 0 143460 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_69
timestamp 1663859327
transform -1 0 144564 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_70
timestamp 1663859327
transform 1 0 142264 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_71
timestamp 1663859327
transform -1 0 143368 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_72
timestamp 1663859327
transform 1 0 141068 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_73
timestamp 1663859327
transform -1 0 142172 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_74
timestamp 1663859327
transform 1 0 139872 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_75
timestamp 1663859327
transform -1 0 140976 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_76
timestamp 1663859327
transform 1 0 138676 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_77
timestamp 1663859327
transform -1 0 139780 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_78
timestamp 1663859327
transform -1 0 138584 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_79
timestamp 1663859327
transform 1 0 137480 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_80
timestamp 1663859327
transform 1 0 136284 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_81
timestamp 1663859327
transform -1 0 137388 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_82
timestamp 1663859327
transform 1 0 135088 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_83
timestamp 1663859327
transform -1 0 136192 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_84
timestamp 1663859327
transform -1 0 155328 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_85
timestamp 1663859327
transform 1 0 154224 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_86
timestamp 1663859327
transform -1 0 394996 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_88
timestamp 1663859327
transform -1 0 396192 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_89
timestamp 1663859327
transform 1 0 395088 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_90
timestamp 1663859327
transform 1 0 396284 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_91
timestamp 1663859327
transform -1 0 397388 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_92
timestamp 1663859327
transform -1 0 398584 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_93
timestamp 1663859327
transform 1 0 397480 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_94
timestamp 1663859327
transform -1 0 399780 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_95
timestamp 1663859327
transform 1 0 398676 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_96
timestamp 1663859327
transform 1 0 399872 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_97
timestamp 1663859327
transform 1 0 401068 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_98
timestamp 1663859327
transform -1 0 400976 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_99
timestamp 1663859327
transform -1 0 402172 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_100
timestamp 1663859327
transform 1 0 402264 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_101
timestamp 1663859327
transform 1 0 403460 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_102
timestamp 1663859327
transform 1 0 404656 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_103
timestamp 1663859327
transform -1 0 403368 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_104
timestamp 1663859327
transform -1 0 404564 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_105
timestamp 1663859327
transform -1 0 405760 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_106
timestamp 1663859327
transform -1 0 406956 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_107
timestamp 1663859327
transform 1 0 405852 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_108
timestamp 1663859327
transform -1 0 408152 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_109
timestamp 1663859327
transform 1 0 407048 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_110
timestamp 1663859327
transform 1 0 408244 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_111
timestamp 1663859327
transform -1 0 409348 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_112
timestamp 1663859327
transform 1 0 409440 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_113
timestamp 1663859327
transform -1 0 410544 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_114
timestamp 1663859327
transform 1 0 410636 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_115
timestamp 1663859327
transform -1 0 411740 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_116
timestamp 1663859327
transform 1 0 411832 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_117
timestamp 1663859327
transform -1 0 412936 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_118
timestamp 1663859327
transform -1 0 414132 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_119
timestamp 1663859327
transform 1 0 413028 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_120
timestamp 1663859327
transform -1 0 415328 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_121
timestamp 1663859327
transform 1 0 414224 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_122
timestamp 1663859327
transform 1 0 415420 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_123
timestamp 1663859327
transform -1 0 416524 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_124
timestamp 1663859327
transform 1 0 416616 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_125
timestamp 1663859327
transform -1 0 418916 0 1 222337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_126
timestamp 1663859327
transform -1 0 417720 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_127
timestamp 1663859327
transform -1 0 418916 0 -1 223425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_128
timestamp 1663859327
transform 0 -1 40864 -1 0 335777
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_129
timestamp 1663859327
transform 0 1 39776 1 0 334673
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_130
timestamp 1663859327
transform 0 -1 40864 -1 0 336973
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_131
timestamp 1663859327
transform 0 1 39776 1 0 335869
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_132
timestamp 1663859327
transform 0 -1 40864 -1 0 338169
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_133
timestamp 1663859327
transform 0 1 39776 1 0 337065
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_134
timestamp 1663859327
transform 0 -1 40864 -1 0 341757
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_135
timestamp 1663859327
transform 0 1 39776 1 0 340653
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_136
timestamp 1663859327
transform 0 -1 40864 -1 0 340561
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_137
timestamp 1663859327
transform 0 1 39776 1 0 339457
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_138
timestamp 1663859327
transform 0 1 39776 1 0 338261
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_139
timestamp 1663859327
transform 0 -1 40864 -1 0 339365
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_140
timestamp 1663859327
transform 0 1 39776 1 0 343045
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_141
timestamp 1663859327
transform 0 -1 40864 -1 0 344149
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_142
timestamp 1663859327
transform 0 1 39776 1 0 341849
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_143
timestamp 1663859327
transform 0 -1 40864 -1 0 342953
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_144
timestamp 1663859327
transform 0 -1 40864 -1 0 347737
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_145
timestamp 1663859327
transform 0 1 39776 1 0 346633
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_146
timestamp 1663859327
transform 0 1 39776 1 0 345437
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_147
timestamp 1663859327
transform 0 -1 40864 -1 0 346541
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_148
timestamp 1663859327
transform 0 1 39776 1 0 344241
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_149
timestamp 1663859327
transform 0 -1 40864 -1 0 345345
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_150
timestamp 1663859327
transform 0 -1 40864 -1 0 351325
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_151
timestamp 1663859327
transform 0 1 39776 1 0 350221
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_152
timestamp 1663859327
transform 0 -1 40864 -1 0 350129
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_153
timestamp 1663859327
transform 0 1 39776 1 0 349025
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_154
timestamp 1663859327
transform 0 1 39776 1 0 347829
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_155
timestamp 1663859327
transform 0 -1 40864 -1 0 348933
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_156
timestamp 1663859327
transform 0 -1 40864 -1 0 352521
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_157
timestamp 1663859327
transform 0 1 39776 1 0 351417
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_158
timestamp 1663859327
transform 0 1 39754 1 0 609598
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_159
timestamp 1663859327
transform 0 -1 40842 -1 0 610702
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_160
timestamp 1663859327
transform 0 1 39754 1 0 608402
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_161
timestamp 1663859327
transform 0 -1 40842 -1 0 609506
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_162
timestamp 1663859327
transform 0 1 39754 1 0 607206
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_163
timestamp 1663859327
transform 0 -1 40842 -1 0 608310
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_164
timestamp 1663859327
transform 0 1 39754 1 0 606010
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_165
timestamp 1663859327
transform 0 -1 40842 -1 0 607114
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_166
timestamp 1663859327
transform 0 1 39754 1 0 604814
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_167
timestamp 1663859327
transform 0 -1 40842 -1 0 605918
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_168
timestamp 1663859327
transform 0 1 39754 1 0 603618
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_169
timestamp 1663859327
transform 0 -1 40842 -1 0 604722
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_170
timestamp 1663859327
transform 0 1 39754 1 0 602422
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_171
timestamp 1663859327
transform 0 -1 40842 -1 0 603526
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_172
timestamp 1663859327
transform 0 -1 40842 -1 0 602330
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_173
timestamp 1663859327
transform 0 1 39754 1 0 601226
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_174
timestamp 1663859327
transform 0 1 39754 1 0 600030
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_175
timestamp 1663859327
transform 0 -1 40842 -1 0 601134
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_176
timestamp 1663859327
transform 0 1 39754 1 0 598834
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_177
timestamp 1663859327
transform 0 -1 40842 -1 0 599938
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_178
timestamp 1663859327
transform 0 1 39754 1 0 597638
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_179
timestamp 1663859327
transform 0 -1 40842 -1 0 598742
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_180
timestamp 1663859327
transform 1 0 662659 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_181
timestamp 1663859327
transform 0 -1 40817 -1 0 890152
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_182
timestamp 1663859327
transform 0 1 39729 1 0 889048
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_183
timestamp 1663859327
transform 0 -1 40817 -1 0 891348
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_184
timestamp 1663859327
transform 0 1 39729 1 0 890244
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_185
timestamp 1663859327
transform 0 1 39729 1 0 885460
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_186
timestamp 1663859327
transform 0 -1 40817 -1 0 886564
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_187
timestamp 1663859327
transform 0 1 39729 1 0 886656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_188
timestamp 1663859327
transform 0 -1 40817 -1 0 887760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_189
timestamp 1663859327
transform 0 -1 40817 -1 0 888956
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_190
timestamp 1663859327
transform 0 1 39729 1 0 887852
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_191
timestamp 1663859327
transform 1 0 663855 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_192
timestamp 1663859327
transform 1 0 665051 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_193
timestamp 1663859327
transform 1 0 666247 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_194
timestamp 1663859327
transform -1 0 663763 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_195
timestamp 1663859327
transform -1 0 664959 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_196
timestamp 1663859327
transform -1 0 666155 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_197
timestamp 1663859327
transform -1 0 667351 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 0 -1 677805 -1 0 707304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1663859327
transform 0 -1 677805 -1 0 708500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1663859327
transform -1 0 133892 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1663859327
transform -1 0 155420 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1663859327
transform -1 0 155420 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1663859327
transform -1 0 153028 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1663859327
transform -1 0 153028 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1663859327
transform -1 0 156616 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1663859327
transform -1 0 156616 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1663859327
transform -1 0 157812 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1663859327
transform -1 0 157812 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1663859327
transform -1 0 159008 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1663859327
transform -1 0 159008 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1663859327
transform 1 0 417762 0 1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1663859327
transform 1 0 417762 0 -1 997540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1663859327
transform 0 1 676717 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1663859327
transform 0 -1 677805 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1663859327
transform 0 1 676717 -1 0 451264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1663859327
transform 0 -1 677805 -1 0 451264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1663859327
transform 0 1 676717 -1 0 448872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1663859327
transform 0 -1 677805 -1 0 448872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1663859327
transform 0 1 676717 -1 0 450068
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1663859327
transform 0 -1 677805 -1 0 450068
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1663859327
transform 0 1 676717 -1 0 452460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1663859327
transform 0 -1 677805 -1 0 452460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1663859327
transform 0 -1 677805 -1 0 453656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1663859327
transform 0 1 676717 -1 0 453656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1663859327
transform 0 1 676717 -1 0 707304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1663859327
transform 0 1 676717 -1 0 708500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1663859327
transform 0 1 676717 -1 0 709696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1663859327
transform 0 -1 677805 -1 0 709696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1663859327
transform 0 1 676717 -1 0 710892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1663859327
transform 0 -1 677805 -1 0 710892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1663859327
transform 0 1 676717 -1 0 712088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1663859327
transform 0 -1 677805 -1 0 712088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1663859327
transform 0 1 676717 -1 0 714480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1663859327
transform 0 -1 677805 -1 0 714480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1663859327
transform 0 1 676717 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1663859327
transform 0 -1 677805 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1663859327
transform 1 0 416566 0 1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1663859327
transform 1 0 416566 0 -1 997540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1663859327
transform -1 0 169414 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1663859327
transform -1 0 169414 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1663859327
transform 0 -1 677805 -1 0 713284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1663859327
transform 0 1 676717 -1 0 713284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1663859327
transform -1 0 170610 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1663859327
transform -1 0 170610 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1663859327
transform -1 0 168218 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1663859327
transform -1 0 168218 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1663859327
transform -1 0 167022 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1663859327
transform -1 0 167022 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1663859327
transform 0 -1 677805 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1663859327
transform 0 1 676717 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1663859327
transform 0 -1 677805 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1663859327
transform 0 1 676717 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1663859327
transform 0 -1 677805 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1663859327
transform 0 1 676717 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1663859327
transform 0 -1 677805 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1663859327
transform 0 1 676717 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1663859327
transform 0 -1 677805 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1663859327
transform 0 1 676717 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1663859327
transform 0 -1 677805 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1663859327
transform 0 1 676717 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1663859327
transform -1 0 151832 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1663859327
transform -1 0 151832 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1663859327
transform -1 0 150636 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1663859327
transform -1 0 150636 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1663859327
transform -1 0 149440 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1663859327
transform -1 0 149440 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1663859327
transform -1 0 148244 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1663859327
transform -1 0 148244 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1663859327
transform -1 0 147048 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1663859327
transform -1 0 147048 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1663859327
transform -1 0 145852 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1663859327
transform -1 0 145852 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1663859327
transform -1 0 144656 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1663859327
transform -1 0 144656 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1663859327
transform -1 0 143460 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1663859327
transform -1 0 143460 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1663859327
transform -1 0 142264 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1663859327
transform -1 0 142264 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1663859327
transform -1 0 141068 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1663859327
transform -1 0 141068 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1663859327
transform -1 0 139872 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1663859327
transform -1 0 139872 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1663859327
transform -1 0 138676 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1663859327
transform -1 0 138676 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1663859327
transform -1 0 137480 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1663859327
transform -1 0 137480 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1663859327
transform -1 0 136284 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1663859327
transform -1 0 136284 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1663859327
transform -1 0 135088 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1663859327
transform -1 0 135088 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1663859327
transform -1 0 154224 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1663859327
transform -1 0 154224 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1663859327
transform -1 0 393892 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1663859327
transform -1 0 395088 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1663859327
transform -1 0 395088 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1663859327
transform -1 0 396284 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1663859327
transform -1 0 396284 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1663859327
transform -1 0 398676 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1663859327
transform -1 0 398676 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1663859327
transform -1 0 397480 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1663859327
transform -1 0 397480 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1663859327
transform -1 0 399872 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1663859327
transform -1 0 401068 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1663859327
transform -1 0 402264 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1663859327
transform -1 0 399872 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1663859327
transform -1 0 401068 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1663859327
transform -1 0 402264 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1663859327
transform -1 0 403460 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1663859327
transform -1 0 404656 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1663859327
transform -1 0 403460 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1663859327
transform -1 0 404656 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1663859327
transform -1 0 405852 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1663859327
transform -1 0 405852 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1663859327
transform -1 0 407048 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1663859327
transform -1 0 407048 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1663859327
transform -1 0 408244 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1663859327
transform -1 0 408244 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1663859327
transform -1 0 409440 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1663859327
transform -1 0 409440 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1663859327
transform -1 0 410636 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1663859327
transform -1 0 410636 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1663859327
transform -1 0 411832 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1663859327
transform -1 0 411832 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1663859327
transform -1 0 413028 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1663859327
transform -1 0 413028 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1663859327
transform -1 0 414224 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1663859327
transform -1 0 414224 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1663859327
transform -1 0 415420 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1663859327
transform -1 0 415420 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1663859327
transform -1 0 416616 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1663859327
transform -1 0 417812 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1663859327
transform -1 0 419008 0 1 222337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1663859327
transform -1 0 416616 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1663859327
transform -1 0 417812 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1663859327
transform -1 0 419008 0 -1 223425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1663859327
transform 0 -1 40864 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1663859327
transform 0 1 39776 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1663859327
transform 0 -1 40864 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1663859327
transform 0 1 39776 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1663859327
transform 0 -1 40864 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1663859327
transform 0 1 39776 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1663859327
transform 0 1 39776 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1663859327
transform 0 -1 40864 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1663859327
transform 0 1 39776 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1663859327
transform 0 -1 40864 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1663859327
transform 0 1 39776 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1663859327
transform 0 -1 40864 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1663859327
transform 0 -1 40864 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1663859327
transform 0 1 39776 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1663859327
transform 0 -1 40864 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1663859327
transform 0 1 39776 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1663859327
transform 0 -1 40864 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1663859327
transform 0 1 39776 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1663859327
transform 0 -1 40864 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1663859327
transform 0 1 39776 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1663859327
transform 0 -1 40864 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1663859327
transform 0 1 39776 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1663859327
transform 0 -1 40864 -1 0 350221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1663859327
transform 0 1 39776 -1 0 350221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1663859327
transform 0 -1 40864 -1 0 349025
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1663859327
transform 0 1 39776 -1 0 349025
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1663859327
transform 0 1 39776 -1 0 347829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1663859327
transform 0 -1 40864 -1 0 347829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1663859327
transform 0 1 39776 -1 0 352613
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1663859327
transform 0 -1 40864 -1 0 352613
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1663859327
transform 0 -1 40864 -1 0 351417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1663859327
transform 0 1 39776 -1 0 351417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1663859327
transform 0 1 39754 -1 0 610794
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1663859327
transform 0 -1 40842 -1 0 610794
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1663859327
transform 0 1 39754 -1 0 609598
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1663859327
transform 0 -1 40842 -1 0 609598
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1663859327
transform 0 1 39754 -1 0 608402
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1663859327
transform 0 -1 40842 -1 0 608402
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1663859327
transform 0 1 39754 -1 0 607206
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1663859327
transform 0 -1 40842 -1 0 607206
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1663859327
transform 0 1 39754 -1 0 606010
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1663859327
transform 0 -1 40842 -1 0 606010
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1663859327
transform 0 1 39754 -1 0 604814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1663859327
transform 0 -1 40842 -1 0 604814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1663859327
transform 0 1 39754 -1 0 603618
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1663859327
transform 0 -1 40842 -1 0 603618
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1663859327
transform 0 -1 40842 -1 0 602422
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1663859327
transform 0 1 39754 -1 0 602422
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1663859327
transform 0 1 39754 -1 0 601226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1663859327
transform 0 -1 40842 -1 0 601226
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1663859327
transform 0 1 39754 -1 0 598834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1663859327
transform 0 1 39754 -1 0 600030
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1663859327
transform 0 -1 40842 -1 0 598834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1663859327
transform 0 -1 40842 -1 0 600030
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1663859327
transform 0 1 39754 -1 0 597638
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1663859327
transform 0 -1 40842 -1 0 597638
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1663859327
transform 0 1 39729 -1 0 890244
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1663859327
transform 0 -1 40817 -1 0 890244
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1663859327
transform 0 -1 40817 -1 0 891440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1663859327
transform 0 1 39729 -1 0 891440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1663859327
transform 0 -1 40817 -1 0 885460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1663859327
transform 0 1 39729 -1 0 885460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1663859327
transform 0 -1 40817 -1 0 886656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1663859327
transform 0 1 39729 -1 0 886656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1663859327
transform 0 1 39729 -1 0 887852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1663859327
transform 0 -1 40817 -1 0 887852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1663859327
transform 0 1 39729 -1 0 889048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1663859327
transform 0 -1 40817 -1 0 889048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1663859327
transform 1 0 662567 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1663859327
transform 1 0 663763 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1663859327
transform 1 0 664959 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1663859327
transform 1 0 666155 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1663859327
transform 1 0 662567 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1663859327
transform 1 0 663763 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1663859327
transform 1 0 664959 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1663859327
transform 1 0 666155 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1663859327
transform 1 0 667351 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1663859327
transform 1 0 667351 0 -1 997458
box -38 -48 130 592
<< labels >>
flabel metal1 416107 995163 416416 995191 0 FreeSans 288 0 0 0 mgmt_io_out_buf[18]
port 1 nsew signal output
flabel metal1 661923 994827 662232 994855 0 FreeSans 288 0 0 0 mgmt_io_out_buf[15]
port 7 nsew signal output
flabel metal1 674476 714634 674504 714921 0 FreeSans 288 90 0 0 mgmt_io_out_buf[13]
port 12 nsew signal output
flabel metal1 673804 453768 673832 454055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[7]
port 19 nsew signal output
flabel metal1 133123 223608 133374 223636 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[37]
port 93 nsew signal output
flabel metal1 170830 995121 171110 995149 0 FreeSans 288 0 0 0 mgmt_io_out_buf[21]
port 54 nsew signal output
flabel metal1 42995 891682 43023 891917 0 FreeSans 288 90 0 0 mgmt_io_out_buf[23]
port 59 nsew signal output
flabel metal1 43639 611095 43667 611356 0 FreeSans 288 90 0 0 mgmt_io_out_buf[29]
port 67 nsew signal output
flabel metal3 664263 997712 664569 997806 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 665458 997701 665764 997795 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 418245 997803 418551 997897 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 417057 997799 417363 997893 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 169809 997465 170115 997559 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 168616 997465 168922 997559 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 146226 221997 146532 222091 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 147432 221997 147738 222091 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 405051 221984 405357 222078 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 406244 221978 406550 222072 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 39436 343400 39526 343697 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 39434 342201 39524 342498 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 39413 605236 39503 605533 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 39413 604045 39503 604342 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 39382 889409 39472 889706 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 39385 888211 39475 888508 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 678061 710130 678151 710427 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 678070 711327 678160 711624 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 678062 446931 678152 447228 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 678064 448130 678154 448427 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal1 673832 215050 673860 215337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[7]
port 25 nsew signal input
flabel metal1 673720 215050 673748 215333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[33]
port 105 nsew signal input
flabel metal1 673888 214850 673916 215137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[7]
port 48 nsew signal output
flabel metal1 673944 214650 673972 214937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[8]
port 26 nsew signal input
flabel metal1 674000 214450 674028 214737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[8]
port 47 nsew signal output
flabel metal1 674056 214250 674084 214537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[9]
port 27 nsew signal input
flabel metal1 674112 214050 674140 214337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[9]
port 46 nsew signal output
flabel metal1 674168 213850 674196 214137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[10]
port 28 nsew signal input
flabel metal1 674224 213650 674252 213937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[10]
port 45 nsew signal output
flabel metal1 674280 213450 674308 213737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[11]
port 29 nsew signal input
flabel metal1 674336 213250 674364 213537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[11]
port 44 nsew signal output
flabel metal1 674392 213050 674420 213337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[12]
port 30 nsew signal input
flabel metal1 674448 212850 674476 213137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[12]
port 43 nsew signal output
flabel metal1 674504 212650 674532 212937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[13]
port 31 nsew signal input
flabel metal1 674560 212450 674588 212737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[13]
port 42 nsew signal output
flabel metal1 674616 212250 674644 212537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[14]
port 32 nsew signal input
flabel metal1 674672 212050 674700 212337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[14]
port 41 nsew signal output
flabel metal1 674728 211850 674756 212137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[15]
port 33 nsew signal input
flabel metal1 674784 211650 674812 211937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[15]
port 40 nsew signal output
flabel metal1 674840 211450 674868 211737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[16]
port 34 nsew signal input
flabel metal1 674896 211250 674924 211537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[16]
port 39 nsew signal output
flabel metal1 674952 211050 674980 211337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[17]
port 35 nsew signal input
flabel metal1 675008 210850 675036 211137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[17]
port 38 nsew signal output
flabel metal1 675064 210650 675092 210937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[18]
port 36 nsew signal input
flabel metal1 675120 210450 675148 210737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[18]
port 37 nsew signal output
flabel metal1 673664 215250 673692 215533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[33]
port 134 nsew signal output
flabel metal1 673608 215450 673636 215733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[32]
port 106 nsew signal input
flabel metal1 673552 215650 673580 215933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[32]
port 133 nsew signal output
flabel metal1 673496 215850 673524 216133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[31]
port 107 nsew signal input
flabel metal1 673440 216050 673468 216333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[31]
port 132 nsew signal output
flabel metal1 673384 216250 673412 216533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[30]
port 108 nsew signal input
flabel metal1 673328 216450 673356 216733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[30]
port 131 nsew signal output
flabel metal1 673272 216650 673300 216933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[29]
port 109 nsew signal input
flabel metal1 673216 216850 673244 217133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[29]
port 130 nsew signal output
flabel metal1 673160 217050 673188 217333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[28]
port 110 nsew signal input
flabel metal1 673104 217250 673132 217533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[28]
port 129 nsew signal output
flabel metal1 673048 217450 673076 217733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[27]
port 111 nsew signal input
flabel metal1 672992 217650 673020 217933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[27]
port 128 nsew signal output
flabel metal1 672936 217850 672964 218133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[26]
port 112 nsew signal input
flabel metal1 672880 218050 672908 218333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[26]
port 127 nsew signal output
flabel metal1 672824 218250 672852 218533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[25]
port 113 nsew signal input
flabel metal1 672768 218450 672796 218733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[25]
port 126 nsew signal output
flabel metal1 672712 218650 672740 218933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[24]
port 114 nsew signal input
flabel metal1 672656 218850 672684 219133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[24]
port 125 nsew signal output
flabel metal1 672600 219050 672628 219333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[23]
port 115 nsew signal input
flabel metal1 672544 219250 672572 219533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[23]
port 124 nsew signal output
flabel metal1 672488 219450 672516 219733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[22]
port 116 nsew signal input
flabel metal1 672432 219650 672460 219933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[22]
port 123 nsew signal output
flabel metal1 672376 219850 672404 220133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[21]
port 117 nsew signal input
flabel metal1 672320 220050 672348 220333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[21]
port 122 nsew signal output
flabel metal1 672264 220250 672292 220533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[20]
port 118 nsew signal input
flabel metal1 672208 220450 672236 220733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[20]
port 121 nsew signal output
flabel metal1 672152 220650 672180 220933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[19]
port 119 nsew signal input
flabel metal1 671480 223050 671508 223287 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[37]
port 94 nsew signal input
flabel metal1 672096 220850 672124 221133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[19]
port 120 nsew signal output
flabel metal1 672040 221050 672068 221287 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[34]
port 101 nsew signal input
flabel metal1 671984 221250 672012 221487 0 FreeSans 288 90 0 0 mgmt_io_in_buf[34]
port 100 nsew signal output
flabel metal1 671928 221450 671956 221687 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[35]
port 102 nsew signal input
flabel metal1 671872 221650 671900 221887 0 FreeSans 288 90 0 0 mgmt_io_in_buf[35]
port 99 nsew signal output
flabel metal1 671816 221850 671844 222087 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[36]
port 103 nsew signal input
flabel metal1 671760 222050 671788 222287 0 FreeSans 288 90 0 0 mgmt_io_in_buf[36]
port 98 nsew signal output
flabel metal1 671704 222250 671732 222487 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[37]
port 104 nsew signal input
flabel metal1 671648 222450 671676 222687 0 FreeSans 288 90 0 0 mgmt_io_in_buf[37]
port 97 nsew signal output
flabel metal1 671592 222650 671620 222887 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[35]
port 96 nsew signal input
flabel metal1 671536 222850 671564 223087 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[36]
port 95 nsew signal input
flabel metal1 132923 223664 133174 223692 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[36]
port 92 nsew signal output
flabel metal1 132723 223720 132974 223748 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[35]
port 91 nsew signal output
flabel metal1 132523 223776 132774 223804 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[37]
port 87 nsew signal input
flabel metal1 132323 223832 132574 223860 0 FreeSans 288 0 0 0 mgmt_io_out_buf[37]
port 86 nsew signal output
flabel metal1 132123 223888 132374 223916 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[36]
port 88 nsew signal input
flabel metal1 131923 223944 132174 223972 0 FreeSans 288 0 0 0 mgmt_io_out_buf[36]
port 85 nsew signal output
flabel metal1 131723 224000 131974 224028 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[35]
port 89 nsew signal input
flabel metal1 131523 224056 131774 224084 0 FreeSans 288 0 0 0 mgmt_io_out_buf[35]
port 84 nsew signal output
flabel metal1 131323 224112 131574 224140 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[34]
port 90 nsew signal input
flabel metal1 131123 224168 131374 224196 0 FreeSans 288 0 0 0 mgmt_io_out_buf[34]
port 83 nsew signal output
flabel metal1 44003 353236 44031 353530 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[33]
port 78 nsew signal input
flabel metal1 43947 353436 43975 353730 0 FreeSans 288 90 0 0 mgmt_io_out_buf[32]
port 76 nsew signal output
flabel metal1 43891 353636 43919 353930 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[32]
port 79 nsew signal input
flabel metal1 43835 353836 43863 354130 0 FreeSans 288 90 0 0 mgmt_io_out_buf[31]
port 75 nsew signal output
flabel metal1 43779 354036 43807 354330 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[31]
port 80 nsew signal input
flabel metal1 43723 354236 43751 354530 0 FreeSans 288 90 0 0 mgmt_io_out_buf[30]
port 74 nsew signal output
flabel metal1 43667 354436 43695 354730 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[30]
port 81 nsew signal input
flabel metal1 43583 611295 43611 611556 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[29]
port 68 nsew signal input
flabel metal1 43527 611495 43555 611756 0 FreeSans 288 90 0 0 mgmt_io_out_buf[28]
port 66 nsew signal output
flabel metal1 43471 611695 43499 611956 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[28]
port 69 nsew signal input
flabel metal1 43415 611895 43443 612156 0 FreeSans 288 90 0 0 mgmt_io_out_buf[27]
port 65 nsew signal output
flabel metal1 43359 612095 43387 612356 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[27]
port 70 nsew signal input
flabel metal1 43303 612295 43331 612556 0 FreeSans 288 90 0 0 mgmt_io_out_buf[26]
port 64 nsew signal output
flabel metal1 43247 612495 43275 612756 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[26]
port 71 nsew signal input
flabel metal1 43191 612695 43219 612956 0 FreeSans 288 90 0 0 mgmt_io_out_buf[25]
port 63 nsew signal output
flabel metal1 43135 612895 43163 613156 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[25]
port 72 nsew signal input
flabel metal1 43079 613095 43107 613356 0 FreeSans 288 90 0 0 mgmt_io_out_buf[24]
port 62 nsew signal output
flabel metal1 43023 613295 43051 613556 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[24]
port 73 nsew signal input
flabel metal1 42939 891882 42967 892117 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[23]
port 60 nsew signal input
flabel metal1 42883 892082 42911 892317 0 FreeSans 288 90 0 0 mgmt_io_out_buf[22]
port 58 nsew signal output
flabel metal1 42827 892282 42855 892517 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[22]
port 61 nsew signal input
flabel metal1 171030 995177 171310 995205 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[21]
port 53 nsew signal input
flabel metal1 171231 995233 171511 995261 0 FreeSans 288 0 0 0 mgmt_io_out_buf[20]
port 55 nsew signal output
flabel metal1 171431 995289 171711 995317 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[20]
port 52 nsew signal input
flabel metal1 171629 995345 171909 995373 0 FreeSans 288 0 0 0 mgmt_io_out_buf[19]
port 56 nsew signal output
flabel metal1 171829 995401 172109 995429 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[19]
port 50 nsew signal input
flabel metal1 415907 995219 416216 995247 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[18]
port 0 nsew signal input
flabel metal1 661723 994883 662032 994911 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[15]
port 6 nsew signal input
flabel metal1 661523 994939 661832 994967 0 FreeSans 288 0 0 0 mgmt_io_out_buf[16]
port 3 nsew signal output
flabel metal1 661323 994995 661632 995023 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[16]
port 5 nsew signal input
flabel metal1 661123 995051 661432 995079 0 FreeSans 288 0 0 0 mgmt_io_out_buf[17]
port 2 nsew signal output
flabel metal1 660923 995107 661232 995135 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[17]
port 4 nsew signal input
flabel metal1 674532 714834 674560 715121 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[13]
port 10 nsew signal input
flabel metal1 674588 715034 674616 715321 0 FreeSans 288 90 0 0 mgmt_io_out_buf[14]
port 11 nsew signal output
flabel metal1 674644 715234 674672 715521 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[14]
port 9 nsew signal input
flabel metal1 673860 453968 673888 454255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[7]
port 18 nsew signal input
flabel metal1 673916 454168 673944 454455 0 FreeSans 288 90 0 0 mgmt_io_out_buf[8]
port 20 nsew signal output
flabel metal1 673972 454368 674000 454655 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[8]
port 17 nsew signal input
flabel metal1 674028 454568 674056 454855 0 FreeSans 288 90 0 0 mgmt_io_out_buf[9]
port 21 nsew signal output
flabel metal1 674084 454768 674112 455055 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[9]
port 16 nsew signal input
flabel metal1 674140 454968 674168 455255 0 FreeSans 288 90 0 0 mgmt_io_out_buf[10]
port 22 nsew signal output
flabel metal1 674196 455168 674224 455455 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[10]
port 15 nsew signal input
flabel metal1 674252 455368 674280 455655 0 FreeSans 288 90 0 0 mgmt_io_out_buf[11]
port 23 nsew signal output
flabel metal1 674308 455568 674336 455855 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[11]
port 14 nsew signal input
flabel metal1 674364 455768 674392 456055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[12]
port 24 nsew signal output
flabel metal1 674420 455968 674448 456255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[12]
port 13 nsew signal input
flabel metal1 44059 353036 44087 353330 0 FreeSans 288 90 0 0 mgmt_io_out_buf[33]
port 77 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
