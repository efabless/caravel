magic
tech sky130A
magscale 1 2
timestamp 1675171987
<< viali >>
rect 2421 2397 2455 2431
<< metal1 >>
rect 92 3834 4232 3856
rect 92 3782 858 3834
rect 910 3782 922 3834
rect 974 3782 986 3834
rect 1038 3782 1050 3834
rect 1102 3782 1114 3834
rect 1166 3782 2378 3834
rect 2430 3782 2442 3834
rect 2494 3782 2506 3834
rect 2558 3782 2570 3834
rect 2622 3782 2634 3834
rect 2686 3782 3898 3834
rect 3950 3782 3962 3834
rect 4014 3782 4026 3834
rect 4078 3782 4090 3834
rect 4142 3782 4154 3834
rect 4206 3782 4232 3834
rect 92 3760 4232 3782
rect 92 3290 4232 3312
rect 92 3238 138 3290
rect 190 3238 202 3290
rect 254 3238 266 3290
rect 318 3238 330 3290
rect 382 3238 394 3290
rect 446 3238 1658 3290
rect 1710 3238 1722 3290
rect 1774 3238 1786 3290
rect 1838 3238 1850 3290
rect 1902 3238 1914 3290
rect 1966 3238 3178 3290
rect 3230 3238 3242 3290
rect 3294 3238 3306 3290
rect 3358 3238 3370 3290
rect 3422 3238 3434 3290
rect 3486 3238 4232 3290
rect 92 3216 4232 3238
rect 92 2746 4232 2768
rect 92 2694 858 2746
rect 910 2694 922 2746
rect 974 2694 986 2746
rect 1038 2694 1050 2746
rect 1102 2694 1114 2746
rect 1166 2694 2378 2746
rect 2430 2694 2442 2746
rect 2494 2694 2506 2746
rect 2558 2694 2570 2746
rect 2622 2694 2634 2746
rect 2686 2694 3898 2746
rect 3950 2694 3962 2746
rect 4014 2694 4026 2746
rect 4078 2694 4090 2746
rect 4142 2694 4154 2746
rect 4206 2694 4232 2746
rect 92 2672 4232 2694
rect 2130 2388 2136 2440
rect 2188 2428 2194 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2188 2400 2421 2428
rect 2188 2388 2194 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 92 2202 4232 2224
rect 92 2150 138 2202
rect 190 2150 202 2202
rect 254 2150 266 2202
rect 318 2150 330 2202
rect 382 2150 394 2202
rect 446 2150 1658 2202
rect 1710 2150 1722 2202
rect 1774 2150 1786 2202
rect 1838 2150 1850 2202
rect 1902 2150 1914 2202
rect 1966 2150 3178 2202
rect 3230 2150 3242 2202
rect 3294 2150 3306 2202
rect 3358 2150 3370 2202
rect 3422 2150 3434 2202
rect 3486 2150 4232 2202
rect 92 2128 4232 2150
rect 92 1658 4232 1680
rect 92 1606 858 1658
rect 910 1606 922 1658
rect 974 1606 986 1658
rect 1038 1606 1050 1658
rect 1102 1606 1114 1658
rect 1166 1606 2378 1658
rect 2430 1606 2442 1658
rect 2494 1606 2506 1658
rect 2558 1606 2570 1658
rect 2622 1606 2634 1658
rect 2686 1606 3898 1658
rect 3950 1606 3962 1658
rect 4014 1606 4026 1658
rect 4078 1606 4090 1658
rect 4142 1606 4154 1658
rect 4206 1606 4232 1658
rect 92 1584 4232 1606
rect 92 1114 4232 1136
rect 92 1062 138 1114
rect 190 1062 202 1114
rect 254 1062 266 1114
rect 318 1062 330 1114
rect 382 1062 394 1114
rect 446 1062 1658 1114
rect 1710 1062 1722 1114
rect 1774 1062 1786 1114
rect 1838 1062 1850 1114
rect 1902 1062 1914 1114
rect 1966 1062 3178 1114
rect 3230 1062 3242 1114
rect 3294 1062 3306 1114
rect 3358 1062 3370 1114
rect 3422 1062 3434 1114
rect 3486 1062 4232 1114
rect 92 1040 4232 1062
rect 92 570 4232 592
rect 92 518 858 570
rect 910 518 922 570
rect 974 518 986 570
rect 1038 518 1050 570
rect 1102 518 1114 570
rect 1166 518 2378 570
rect 2430 518 2442 570
rect 2494 518 2506 570
rect 2558 518 2570 570
rect 2622 518 2634 570
rect 2686 518 3898 570
rect 3950 518 3962 570
rect 4014 518 4026 570
rect 4078 518 4090 570
rect 4142 518 4154 570
rect 4206 518 4232 570
rect 92 496 4232 518
<< via1 >>
rect 858 3782 910 3834
rect 922 3782 974 3834
rect 986 3782 1038 3834
rect 1050 3782 1102 3834
rect 1114 3782 1166 3834
rect 2378 3782 2430 3834
rect 2442 3782 2494 3834
rect 2506 3782 2558 3834
rect 2570 3782 2622 3834
rect 2634 3782 2686 3834
rect 3898 3782 3950 3834
rect 3962 3782 4014 3834
rect 4026 3782 4078 3834
rect 4090 3782 4142 3834
rect 4154 3782 4206 3834
rect 138 3238 190 3290
rect 202 3238 254 3290
rect 266 3238 318 3290
rect 330 3238 382 3290
rect 394 3238 446 3290
rect 1658 3238 1710 3290
rect 1722 3238 1774 3290
rect 1786 3238 1838 3290
rect 1850 3238 1902 3290
rect 1914 3238 1966 3290
rect 3178 3238 3230 3290
rect 3242 3238 3294 3290
rect 3306 3238 3358 3290
rect 3370 3238 3422 3290
rect 3434 3238 3486 3290
rect 858 2694 910 2746
rect 922 2694 974 2746
rect 986 2694 1038 2746
rect 1050 2694 1102 2746
rect 1114 2694 1166 2746
rect 2378 2694 2430 2746
rect 2442 2694 2494 2746
rect 2506 2694 2558 2746
rect 2570 2694 2622 2746
rect 2634 2694 2686 2746
rect 3898 2694 3950 2746
rect 3962 2694 4014 2746
rect 4026 2694 4078 2746
rect 4090 2694 4142 2746
rect 4154 2694 4206 2746
rect 2136 2388 2188 2440
rect 138 2150 190 2202
rect 202 2150 254 2202
rect 266 2150 318 2202
rect 330 2150 382 2202
rect 394 2150 446 2202
rect 1658 2150 1710 2202
rect 1722 2150 1774 2202
rect 1786 2150 1838 2202
rect 1850 2150 1902 2202
rect 1914 2150 1966 2202
rect 3178 2150 3230 2202
rect 3242 2150 3294 2202
rect 3306 2150 3358 2202
rect 3370 2150 3422 2202
rect 3434 2150 3486 2202
rect 858 1606 910 1658
rect 922 1606 974 1658
rect 986 1606 1038 1658
rect 1050 1606 1102 1658
rect 1114 1606 1166 1658
rect 2378 1606 2430 1658
rect 2442 1606 2494 1658
rect 2506 1606 2558 1658
rect 2570 1606 2622 1658
rect 2634 1606 2686 1658
rect 3898 1606 3950 1658
rect 3962 1606 4014 1658
rect 4026 1606 4078 1658
rect 4090 1606 4142 1658
rect 4154 1606 4206 1658
rect 138 1062 190 1114
rect 202 1062 254 1114
rect 266 1062 318 1114
rect 330 1062 382 1114
rect 394 1062 446 1114
rect 1658 1062 1710 1114
rect 1722 1062 1774 1114
rect 1786 1062 1838 1114
rect 1850 1062 1902 1114
rect 1914 1062 1966 1114
rect 3178 1062 3230 1114
rect 3242 1062 3294 1114
rect 3306 1062 3358 1114
rect 3370 1062 3422 1114
rect 3434 1062 3486 1114
rect 858 518 910 570
rect 922 518 974 570
rect 986 518 1038 570
rect 1050 518 1102 570
rect 1114 518 1166 570
rect 2378 518 2430 570
rect 2442 518 2494 570
rect 2506 518 2558 570
rect 2570 518 2622 570
rect 2634 518 2686 570
rect 3898 518 3950 570
rect 3962 518 4014 570
rect 4026 518 4078 570
rect 4090 518 4142 570
rect 4154 518 4206 570
<< metal2 >>
rect 132 3932 452 3944
rect 132 3876 144 3932
rect 200 3876 224 3932
rect 280 3876 304 3932
rect 360 3876 384 3932
rect 440 3876 452 3932
rect 132 3852 452 3876
rect 1652 3932 1972 3944
rect 1652 3876 1664 3932
rect 1720 3876 1744 3932
rect 1800 3876 1824 3932
rect 1880 3876 1904 3932
rect 1960 3876 1972 3932
rect 132 3796 144 3852
rect 200 3796 224 3852
rect 280 3796 304 3852
rect 360 3796 384 3852
rect 440 3796 452 3852
rect 132 3772 452 3796
rect 132 3716 144 3772
rect 200 3716 224 3772
rect 280 3716 304 3772
rect 360 3716 384 3772
rect 440 3716 452 3772
rect 132 3692 452 3716
rect 132 3636 144 3692
rect 200 3636 224 3692
rect 280 3636 304 3692
rect 360 3636 384 3692
rect 440 3636 452 3692
rect 132 3290 452 3636
rect 132 3238 138 3290
rect 190 3238 202 3290
rect 254 3238 266 3290
rect 318 3238 330 3290
rect 382 3238 394 3290
rect 446 3238 452 3290
rect 132 2412 452 3238
rect 132 2356 144 2412
rect 200 2356 224 2412
rect 280 2356 304 2412
rect 360 2356 384 2412
rect 440 2356 452 2412
rect 132 2332 452 2356
rect 132 2276 144 2332
rect 200 2276 224 2332
rect 280 2276 304 2332
rect 360 2276 384 2332
rect 440 2276 452 2332
rect 132 2252 452 2276
rect 132 2202 144 2252
rect 200 2202 224 2252
rect 280 2202 304 2252
rect 360 2202 384 2252
rect 440 2202 452 2252
rect 132 2150 138 2202
rect 200 2196 202 2202
rect 382 2196 384 2202
rect 190 2172 202 2196
rect 254 2172 266 2196
rect 318 2172 330 2196
rect 382 2172 394 2196
rect 200 2150 202 2172
rect 382 2150 384 2172
rect 446 2150 452 2202
rect 132 2116 144 2150
rect 200 2116 224 2150
rect 280 2116 304 2150
rect 360 2116 384 2150
rect 440 2116 452 2150
rect 132 1114 452 2116
rect 132 1062 138 1114
rect 190 1062 202 1114
rect 254 1062 266 1114
rect 318 1062 330 1114
rect 382 1062 394 1114
rect 446 1062 452 1114
rect 132 892 452 1062
rect 132 836 144 892
rect 200 836 224 892
rect 280 836 304 892
rect 360 836 384 892
rect 440 836 452 892
rect 132 812 452 836
rect 132 756 144 812
rect 200 756 224 812
rect 280 756 304 812
rect 360 756 384 812
rect 440 756 452 812
rect 132 732 452 756
rect 132 676 144 732
rect 200 676 224 732
rect 280 676 304 732
rect 360 676 384 732
rect 440 676 452 732
rect 132 652 452 676
rect 132 596 144 652
rect 200 596 224 652
rect 280 596 304 652
rect 360 596 384 652
rect 440 596 452 652
rect 132 496 452 596
rect 852 3834 1172 3856
rect 852 3782 858 3834
rect 910 3782 922 3834
rect 974 3782 986 3834
rect 1038 3782 1050 3834
rect 1102 3782 1114 3834
rect 1166 3782 1172 3834
rect 852 3132 1172 3782
rect 852 3076 864 3132
rect 920 3076 944 3132
rect 1000 3076 1024 3132
rect 1080 3076 1104 3132
rect 1160 3076 1172 3132
rect 852 3052 1172 3076
rect 852 2996 864 3052
rect 920 2996 944 3052
rect 1000 2996 1024 3052
rect 1080 2996 1104 3052
rect 1160 2996 1172 3052
rect 852 2972 1172 2996
rect 852 2916 864 2972
rect 920 2916 944 2972
rect 1000 2916 1024 2972
rect 1080 2916 1104 2972
rect 1160 2916 1172 2972
rect 852 2892 1172 2916
rect 852 2836 864 2892
rect 920 2836 944 2892
rect 1000 2836 1024 2892
rect 1080 2836 1104 2892
rect 1160 2836 1172 2892
rect 852 2746 1172 2836
rect 852 2694 858 2746
rect 910 2694 922 2746
rect 974 2694 986 2746
rect 1038 2694 1050 2746
rect 1102 2694 1114 2746
rect 1166 2694 1172 2746
rect 852 1658 1172 2694
rect 852 1606 858 1658
rect 910 1612 922 1658
rect 974 1612 986 1658
rect 1038 1612 1050 1658
rect 1102 1612 1114 1658
rect 920 1606 922 1612
rect 1102 1606 1104 1612
rect 1166 1606 1172 1658
rect 852 1556 864 1606
rect 920 1556 944 1606
rect 1000 1556 1024 1606
rect 1080 1556 1104 1606
rect 1160 1556 1172 1606
rect 852 1532 1172 1556
rect 852 1476 864 1532
rect 920 1476 944 1532
rect 1000 1476 1024 1532
rect 1080 1476 1104 1532
rect 1160 1476 1172 1532
rect 852 1452 1172 1476
rect 852 1396 864 1452
rect 920 1396 944 1452
rect 1000 1396 1024 1452
rect 1080 1396 1104 1452
rect 1160 1396 1172 1452
rect 852 1372 1172 1396
rect 852 1316 864 1372
rect 920 1316 944 1372
rect 1000 1316 1024 1372
rect 1080 1316 1104 1372
rect 1160 1316 1172 1372
rect 852 570 1172 1316
rect 852 518 858 570
rect 910 518 922 570
rect 974 518 986 570
rect 1038 518 1050 570
rect 1102 518 1114 570
rect 1166 518 1172 570
rect 852 496 1172 518
rect 1652 3852 1972 3876
rect 3172 3932 3492 3944
rect 3172 3876 3184 3932
rect 3240 3876 3264 3932
rect 3320 3876 3344 3932
rect 3400 3876 3424 3932
rect 3480 3876 3492 3932
rect 1652 3796 1664 3852
rect 1720 3796 1744 3852
rect 1800 3796 1824 3852
rect 1880 3796 1904 3852
rect 1960 3796 1972 3852
rect 1652 3772 1972 3796
rect 1652 3716 1664 3772
rect 1720 3716 1744 3772
rect 1800 3716 1824 3772
rect 1880 3716 1904 3772
rect 1960 3716 1972 3772
rect 1652 3692 1972 3716
rect 1652 3636 1664 3692
rect 1720 3636 1744 3692
rect 1800 3636 1824 3692
rect 1880 3636 1904 3692
rect 1960 3636 1972 3692
rect 1652 3290 1972 3636
rect 1652 3238 1658 3290
rect 1710 3238 1722 3290
rect 1774 3238 1786 3290
rect 1838 3238 1850 3290
rect 1902 3238 1914 3290
rect 1966 3238 1972 3290
rect 1652 2412 1972 3238
rect 2372 3834 2692 3856
rect 2372 3782 2378 3834
rect 2430 3782 2442 3834
rect 2494 3782 2506 3834
rect 2558 3782 2570 3834
rect 2622 3782 2634 3834
rect 2686 3782 2692 3834
rect 2372 3132 2692 3782
rect 2372 3076 2384 3132
rect 2440 3076 2464 3132
rect 2520 3076 2544 3132
rect 2600 3076 2624 3132
rect 2680 3076 2692 3132
rect 2372 3052 2692 3076
rect 2372 2996 2384 3052
rect 2440 2996 2464 3052
rect 2520 2996 2544 3052
rect 2600 2996 2624 3052
rect 2680 2996 2692 3052
rect 2372 2972 2692 2996
rect 2372 2916 2384 2972
rect 2440 2916 2464 2972
rect 2520 2916 2544 2972
rect 2600 2916 2624 2972
rect 2680 2916 2692 2972
rect 2372 2892 2692 2916
rect 2372 2836 2384 2892
rect 2440 2836 2464 2892
rect 2520 2836 2544 2892
rect 2600 2836 2624 2892
rect 2680 2836 2692 2892
rect 2372 2746 2692 2836
rect 2372 2694 2378 2746
rect 2430 2694 2442 2746
rect 2494 2694 2506 2746
rect 2558 2694 2570 2746
rect 2622 2694 2634 2746
rect 2686 2694 2692 2746
rect 1652 2356 1664 2412
rect 1720 2356 1744 2412
rect 1800 2356 1824 2412
rect 1880 2356 1904 2412
rect 1960 2356 1972 2412
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 1652 2332 1972 2356
rect 1652 2276 1664 2332
rect 1720 2276 1744 2332
rect 1800 2276 1824 2332
rect 1880 2276 1904 2332
rect 1960 2276 1972 2332
rect 1652 2252 1972 2276
rect 1652 2202 1664 2252
rect 1720 2202 1744 2252
rect 1800 2202 1824 2252
rect 1880 2202 1904 2252
rect 1960 2202 1972 2252
rect 1652 2150 1658 2202
rect 1720 2196 1722 2202
rect 1902 2196 1904 2202
rect 1710 2172 1722 2196
rect 1774 2172 1786 2196
rect 1838 2172 1850 2196
rect 1902 2172 1914 2196
rect 1720 2150 1722 2172
rect 1902 2150 1904 2172
rect 1966 2150 1972 2202
rect 1652 2116 1664 2150
rect 1720 2116 1744 2150
rect 1800 2116 1824 2150
rect 1880 2116 1904 2150
rect 1960 2116 1972 2150
rect 1652 1114 1972 2116
rect 1652 1062 1658 1114
rect 1710 1062 1722 1114
rect 1774 1062 1786 1114
rect 1838 1062 1850 1114
rect 1902 1062 1914 1114
rect 1966 1062 1972 1114
rect 1652 892 1972 1062
rect 1652 836 1664 892
rect 1720 836 1744 892
rect 1800 836 1824 892
rect 1880 836 1904 892
rect 1960 836 1972 892
rect 1652 812 1972 836
rect 1652 756 1664 812
rect 1720 756 1744 812
rect 1800 756 1824 812
rect 1880 756 1904 812
rect 1960 756 1972 812
rect 1652 732 1972 756
rect 1652 676 1664 732
rect 1720 676 1744 732
rect 1800 676 1824 732
rect 1880 676 1904 732
rect 1960 676 1972 732
rect 1652 652 1972 676
rect 1652 596 1664 652
rect 1720 596 1744 652
rect 1800 596 1824 652
rect 1880 596 1904 652
rect 1960 596 1972 652
rect 1652 496 1972 596
rect 2148 400 2176 2382
rect 2372 1658 2692 2694
rect 2372 1606 2378 1658
rect 2430 1612 2442 1658
rect 2494 1612 2506 1658
rect 2558 1612 2570 1658
rect 2622 1612 2634 1658
rect 2440 1606 2442 1612
rect 2622 1606 2624 1612
rect 2686 1606 2692 1658
rect 2372 1556 2384 1606
rect 2440 1556 2464 1606
rect 2520 1556 2544 1606
rect 2600 1556 2624 1606
rect 2680 1556 2692 1606
rect 2372 1532 2692 1556
rect 2372 1476 2384 1532
rect 2440 1476 2464 1532
rect 2520 1476 2544 1532
rect 2600 1476 2624 1532
rect 2680 1476 2692 1532
rect 2372 1452 2692 1476
rect 2372 1396 2384 1452
rect 2440 1396 2464 1452
rect 2520 1396 2544 1452
rect 2600 1396 2624 1452
rect 2680 1396 2692 1452
rect 2372 1372 2692 1396
rect 2372 1316 2384 1372
rect 2440 1316 2464 1372
rect 2520 1316 2544 1372
rect 2600 1316 2624 1372
rect 2680 1316 2692 1372
rect 2372 570 2692 1316
rect 2372 518 2378 570
rect 2430 518 2442 570
rect 2494 518 2506 570
rect 2558 518 2570 570
rect 2622 518 2634 570
rect 2686 518 2692 570
rect 2372 496 2692 518
rect 3172 3852 3492 3876
rect 3172 3796 3184 3852
rect 3240 3796 3264 3852
rect 3320 3796 3344 3852
rect 3400 3796 3424 3852
rect 3480 3796 3492 3852
rect 3172 3772 3492 3796
rect 3172 3716 3184 3772
rect 3240 3716 3264 3772
rect 3320 3716 3344 3772
rect 3400 3716 3424 3772
rect 3480 3716 3492 3772
rect 3172 3692 3492 3716
rect 3172 3636 3184 3692
rect 3240 3636 3264 3692
rect 3320 3636 3344 3692
rect 3400 3636 3424 3692
rect 3480 3636 3492 3692
rect 3172 3290 3492 3636
rect 3172 3238 3178 3290
rect 3230 3238 3242 3290
rect 3294 3238 3306 3290
rect 3358 3238 3370 3290
rect 3422 3238 3434 3290
rect 3486 3238 3492 3290
rect 3172 2412 3492 3238
rect 3172 2356 3184 2412
rect 3240 2356 3264 2412
rect 3320 2356 3344 2412
rect 3400 2356 3424 2412
rect 3480 2356 3492 2412
rect 3172 2332 3492 2356
rect 3172 2276 3184 2332
rect 3240 2276 3264 2332
rect 3320 2276 3344 2332
rect 3400 2276 3424 2332
rect 3480 2276 3492 2332
rect 3172 2252 3492 2276
rect 3172 2202 3184 2252
rect 3240 2202 3264 2252
rect 3320 2202 3344 2252
rect 3400 2202 3424 2252
rect 3480 2202 3492 2252
rect 3172 2150 3178 2202
rect 3240 2196 3242 2202
rect 3422 2196 3424 2202
rect 3230 2172 3242 2196
rect 3294 2172 3306 2196
rect 3358 2172 3370 2196
rect 3422 2172 3434 2196
rect 3240 2150 3242 2172
rect 3422 2150 3424 2172
rect 3486 2150 3492 2202
rect 3172 2116 3184 2150
rect 3240 2116 3264 2150
rect 3320 2116 3344 2150
rect 3400 2116 3424 2150
rect 3480 2116 3492 2150
rect 3172 1114 3492 2116
rect 3172 1062 3178 1114
rect 3230 1062 3242 1114
rect 3294 1062 3306 1114
rect 3358 1062 3370 1114
rect 3422 1062 3434 1114
rect 3486 1062 3492 1114
rect 3172 892 3492 1062
rect 3172 836 3184 892
rect 3240 836 3264 892
rect 3320 836 3344 892
rect 3400 836 3424 892
rect 3480 836 3492 892
rect 3172 812 3492 836
rect 3172 756 3184 812
rect 3240 756 3264 812
rect 3320 756 3344 812
rect 3400 756 3424 812
rect 3480 756 3492 812
rect 3172 732 3492 756
rect 3172 676 3184 732
rect 3240 676 3264 732
rect 3320 676 3344 732
rect 3400 676 3424 732
rect 3480 676 3492 732
rect 3172 652 3492 676
rect 3172 596 3184 652
rect 3240 596 3264 652
rect 3320 596 3344 652
rect 3400 596 3424 652
rect 3480 596 3492 652
rect 3172 496 3492 596
rect 3892 3834 4212 3856
rect 3892 3782 3898 3834
rect 3950 3782 3962 3834
rect 4014 3782 4026 3834
rect 4078 3782 4090 3834
rect 4142 3782 4154 3834
rect 4206 3782 4212 3834
rect 3892 3132 4212 3782
rect 3892 3076 3904 3132
rect 3960 3076 3984 3132
rect 4040 3076 4064 3132
rect 4120 3076 4144 3132
rect 4200 3076 4212 3132
rect 3892 3052 4212 3076
rect 3892 2996 3904 3052
rect 3960 2996 3984 3052
rect 4040 2996 4064 3052
rect 4120 2996 4144 3052
rect 4200 2996 4212 3052
rect 3892 2972 4212 2996
rect 3892 2916 3904 2972
rect 3960 2916 3984 2972
rect 4040 2916 4064 2972
rect 4120 2916 4144 2972
rect 4200 2916 4212 2972
rect 3892 2892 4212 2916
rect 3892 2836 3904 2892
rect 3960 2836 3984 2892
rect 4040 2836 4064 2892
rect 4120 2836 4144 2892
rect 4200 2836 4212 2892
rect 3892 2746 4212 2836
rect 3892 2694 3898 2746
rect 3950 2694 3962 2746
rect 4014 2694 4026 2746
rect 4078 2694 4090 2746
rect 4142 2694 4154 2746
rect 4206 2694 4212 2746
rect 3892 1658 4212 2694
rect 3892 1606 3898 1658
rect 3950 1612 3962 1658
rect 4014 1612 4026 1658
rect 4078 1612 4090 1658
rect 4142 1612 4154 1658
rect 3960 1606 3962 1612
rect 4142 1606 4144 1612
rect 4206 1606 4212 1658
rect 3892 1556 3904 1606
rect 3960 1556 3984 1606
rect 4040 1556 4064 1606
rect 4120 1556 4144 1606
rect 4200 1556 4212 1606
rect 3892 1532 4212 1556
rect 3892 1476 3904 1532
rect 3960 1476 3984 1532
rect 4040 1476 4064 1532
rect 4120 1476 4144 1532
rect 4200 1476 4212 1532
rect 3892 1452 4212 1476
rect 3892 1396 3904 1452
rect 3960 1396 3984 1452
rect 4040 1396 4064 1452
rect 4120 1396 4144 1452
rect 4200 1396 4212 1452
rect 3892 1372 4212 1396
rect 3892 1316 3904 1372
rect 3960 1316 3984 1372
rect 4040 1316 4064 1372
rect 4120 1316 4144 1372
rect 4200 1316 4212 1372
rect 3892 570 4212 1316
rect 3892 518 3898 570
rect 3950 518 3962 570
rect 4014 518 4026 570
rect 4078 518 4090 570
rect 4142 518 4154 570
rect 4206 518 4212 570
rect 3892 496 4212 518
rect 2134 0 2190 400
<< via2 >>
rect 144 3876 200 3932
rect 224 3876 280 3932
rect 304 3876 360 3932
rect 384 3876 440 3932
rect 1664 3876 1720 3932
rect 1744 3876 1800 3932
rect 1824 3876 1880 3932
rect 1904 3876 1960 3932
rect 144 3796 200 3852
rect 224 3796 280 3852
rect 304 3796 360 3852
rect 384 3796 440 3852
rect 144 3716 200 3772
rect 224 3716 280 3772
rect 304 3716 360 3772
rect 384 3716 440 3772
rect 144 3636 200 3692
rect 224 3636 280 3692
rect 304 3636 360 3692
rect 384 3636 440 3692
rect 144 2356 200 2412
rect 224 2356 280 2412
rect 304 2356 360 2412
rect 384 2356 440 2412
rect 144 2276 200 2332
rect 224 2276 280 2332
rect 304 2276 360 2332
rect 384 2276 440 2332
rect 144 2202 200 2252
rect 224 2202 280 2252
rect 304 2202 360 2252
rect 384 2202 440 2252
rect 144 2196 190 2202
rect 190 2196 200 2202
rect 224 2196 254 2202
rect 254 2196 266 2202
rect 266 2196 280 2202
rect 304 2196 318 2202
rect 318 2196 330 2202
rect 330 2196 360 2202
rect 384 2196 394 2202
rect 394 2196 440 2202
rect 144 2150 190 2172
rect 190 2150 200 2172
rect 224 2150 254 2172
rect 254 2150 266 2172
rect 266 2150 280 2172
rect 304 2150 318 2172
rect 318 2150 330 2172
rect 330 2150 360 2172
rect 384 2150 394 2172
rect 394 2150 440 2172
rect 144 2116 200 2150
rect 224 2116 280 2150
rect 304 2116 360 2150
rect 384 2116 440 2150
rect 144 836 200 892
rect 224 836 280 892
rect 304 836 360 892
rect 384 836 440 892
rect 144 756 200 812
rect 224 756 280 812
rect 304 756 360 812
rect 384 756 440 812
rect 144 676 200 732
rect 224 676 280 732
rect 304 676 360 732
rect 384 676 440 732
rect 144 596 200 652
rect 224 596 280 652
rect 304 596 360 652
rect 384 596 440 652
rect 864 3076 920 3132
rect 944 3076 1000 3132
rect 1024 3076 1080 3132
rect 1104 3076 1160 3132
rect 864 2996 920 3052
rect 944 2996 1000 3052
rect 1024 2996 1080 3052
rect 1104 2996 1160 3052
rect 864 2916 920 2972
rect 944 2916 1000 2972
rect 1024 2916 1080 2972
rect 1104 2916 1160 2972
rect 864 2836 920 2892
rect 944 2836 1000 2892
rect 1024 2836 1080 2892
rect 1104 2836 1160 2892
rect 864 1606 910 1612
rect 910 1606 920 1612
rect 944 1606 974 1612
rect 974 1606 986 1612
rect 986 1606 1000 1612
rect 1024 1606 1038 1612
rect 1038 1606 1050 1612
rect 1050 1606 1080 1612
rect 1104 1606 1114 1612
rect 1114 1606 1160 1612
rect 864 1556 920 1606
rect 944 1556 1000 1606
rect 1024 1556 1080 1606
rect 1104 1556 1160 1606
rect 864 1476 920 1532
rect 944 1476 1000 1532
rect 1024 1476 1080 1532
rect 1104 1476 1160 1532
rect 864 1396 920 1452
rect 944 1396 1000 1452
rect 1024 1396 1080 1452
rect 1104 1396 1160 1452
rect 864 1316 920 1372
rect 944 1316 1000 1372
rect 1024 1316 1080 1372
rect 1104 1316 1160 1372
rect 3184 3876 3240 3932
rect 3264 3876 3320 3932
rect 3344 3876 3400 3932
rect 3424 3876 3480 3932
rect 1664 3796 1720 3852
rect 1744 3796 1800 3852
rect 1824 3796 1880 3852
rect 1904 3796 1960 3852
rect 1664 3716 1720 3772
rect 1744 3716 1800 3772
rect 1824 3716 1880 3772
rect 1904 3716 1960 3772
rect 1664 3636 1720 3692
rect 1744 3636 1800 3692
rect 1824 3636 1880 3692
rect 1904 3636 1960 3692
rect 2384 3076 2440 3132
rect 2464 3076 2520 3132
rect 2544 3076 2600 3132
rect 2624 3076 2680 3132
rect 2384 2996 2440 3052
rect 2464 2996 2520 3052
rect 2544 2996 2600 3052
rect 2624 2996 2680 3052
rect 2384 2916 2440 2972
rect 2464 2916 2520 2972
rect 2544 2916 2600 2972
rect 2624 2916 2680 2972
rect 2384 2836 2440 2892
rect 2464 2836 2520 2892
rect 2544 2836 2600 2892
rect 2624 2836 2680 2892
rect 1664 2356 1720 2412
rect 1744 2356 1800 2412
rect 1824 2356 1880 2412
rect 1904 2356 1960 2412
rect 1664 2276 1720 2332
rect 1744 2276 1800 2332
rect 1824 2276 1880 2332
rect 1904 2276 1960 2332
rect 1664 2202 1720 2252
rect 1744 2202 1800 2252
rect 1824 2202 1880 2252
rect 1904 2202 1960 2252
rect 1664 2196 1710 2202
rect 1710 2196 1720 2202
rect 1744 2196 1774 2202
rect 1774 2196 1786 2202
rect 1786 2196 1800 2202
rect 1824 2196 1838 2202
rect 1838 2196 1850 2202
rect 1850 2196 1880 2202
rect 1904 2196 1914 2202
rect 1914 2196 1960 2202
rect 1664 2150 1710 2172
rect 1710 2150 1720 2172
rect 1744 2150 1774 2172
rect 1774 2150 1786 2172
rect 1786 2150 1800 2172
rect 1824 2150 1838 2172
rect 1838 2150 1850 2172
rect 1850 2150 1880 2172
rect 1904 2150 1914 2172
rect 1914 2150 1960 2172
rect 1664 2116 1720 2150
rect 1744 2116 1800 2150
rect 1824 2116 1880 2150
rect 1904 2116 1960 2150
rect 1664 836 1720 892
rect 1744 836 1800 892
rect 1824 836 1880 892
rect 1904 836 1960 892
rect 1664 756 1720 812
rect 1744 756 1800 812
rect 1824 756 1880 812
rect 1904 756 1960 812
rect 1664 676 1720 732
rect 1744 676 1800 732
rect 1824 676 1880 732
rect 1904 676 1960 732
rect 1664 596 1720 652
rect 1744 596 1800 652
rect 1824 596 1880 652
rect 1904 596 1960 652
rect 2384 1606 2430 1612
rect 2430 1606 2440 1612
rect 2464 1606 2494 1612
rect 2494 1606 2506 1612
rect 2506 1606 2520 1612
rect 2544 1606 2558 1612
rect 2558 1606 2570 1612
rect 2570 1606 2600 1612
rect 2624 1606 2634 1612
rect 2634 1606 2680 1612
rect 2384 1556 2440 1606
rect 2464 1556 2520 1606
rect 2544 1556 2600 1606
rect 2624 1556 2680 1606
rect 2384 1476 2440 1532
rect 2464 1476 2520 1532
rect 2544 1476 2600 1532
rect 2624 1476 2680 1532
rect 2384 1396 2440 1452
rect 2464 1396 2520 1452
rect 2544 1396 2600 1452
rect 2624 1396 2680 1452
rect 2384 1316 2440 1372
rect 2464 1316 2520 1372
rect 2544 1316 2600 1372
rect 2624 1316 2680 1372
rect 3184 3796 3240 3852
rect 3264 3796 3320 3852
rect 3344 3796 3400 3852
rect 3424 3796 3480 3852
rect 3184 3716 3240 3772
rect 3264 3716 3320 3772
rect 3344 3716 3400 3772
rect 3424 3716 3480 3772
rect 3184 3636 3240 3692
rect 3264 3636 3320 3692
rect 3344 3636 3400 3692
rect 3424 3636 3480 3692
rect 3184 2356 3240 2412
rect 3264 2356 3320 2412
rect 3344 2356 3400 2412
rect 3424 2356 3480 2412
rect 3184 2276 3240 2332
rect 3264 2276 3320 2332
rect 3344 2276 3400 2332
rect 3424 2276 3480 2332
rect 3184 2202 3240 2252
rect 3264 2202 3320 2252
rect 3344 2202 3400 2252
rect 3424 2202 3480 2252
rect 3184 2196 3230 2202
rect 3230 2196 3240 2202
rect 3264 2196 3294 2202
rect 3294 2196 3306 2202
rect 3306 2196 3320 2202
rect 3344 2196 3358 2202
rect 3358 2196 3370 2202
rect 3370 2196 3400 2202
rect 3424 2196 3434 2202
rect 3434 2196 3480 2202
rect 3184 2150 3230 2172
rect 3230 2150 3240 2172
rect 3264 2150 3294 2172
rect 3294 2150 3306 2172
rect 3306 2150 3320 2172
rect 3344 2150 3358 2172
rect 3358 2150 3370 2172
rect 3370 2150 3400 2172
rect 3424 2150 3434 2172
rect 3434 2150 3480 2172
rect 3184 2116 3240 2150
rect 3264 2116 3320 2150
rect 3344 2116 3400 2150
rect 3424 2116 3480 2150
rect 3184 836 3240 892
rect 3264 836 3320 892
rect 3344 836 3400 892
rect 3424 836 3480 892
rect 3184 756 3240 812
rect 3264 756 3320 812
rect 3344 756 3400 812
rect 3424 756 3480 812
rect 3184 676 3240 732
rect 3264 676 3320 732
rect 3344 676 3400 732
rect 3424 676 3480 732
rect 3184 596 3240 652
rect 3264 596 3320 652
rect 3344 596 3400 652
rect 3424 596 3480 652
rect 3904 3076 3960 3132
rect 3984 3076 4040 3132
rect 4064 3076 4120 3132
rect 4144 3076 4200 3132
rect 3904 2996 3960 3052
rect 3984 2996 4040 3052
rect 4064 2996 4120 3052
rect 4144 2996 4200 3052
rect 3904 2916 3960 2972
rect 3984 2916 4040 2972
rect 4064 2916 4120 2972
rect 4144 2916 4200 2972
rect 3904 2836 3960 2892
rect 3984 2836 4040 2892
rect 4064 2836 4120 2892
rect 4144 2836 4200 2892
rect 3904 1606 3950 1612
rect 3950 1606 3960 1612
rect 3984 1606 4014 1612
rect 4014 1606 4026 1612
rect 4026 1606 4040 1612
rect 4064 1606 4078 1612
rect 4078 1606 4090 1612
rect 4090 1606 4120 1612
rect 4144 1606 4154 1612
rect 4154 1606 4200 1612
rect 3904 1556 3960 1606
rect 3984 1556 4040 1606
rect 4064 1556 4120 1606
rect 4144 1556 4200 1606
rect 3904 1476 3960 1532
rect 3984 1476 4040 1532
rect 4064 1476 4120 1532
rect 4144 1476 4200 1532
rect 3904 1396 3960 1452
rect 3984 1396 4040 1452
rect 4064 1396 4120 1452
rect 4144 1396 4200 1452
rect 3904 1316 3960 1372
rect 3984 1316 4040 1372
rect 4064 1316 4120 1372
rect 4144 1316 4200 1372
<< metal3 >>
rect 44 3932 4280 3944
rect 44 3876 144 3932
rect 200 3876 224 3932
rect 280 3876 304 3932
rect 360 3876 384 3932
rect 440 3876 1664 3932
rect 1720 3876 1744 3932
rect 1800 3876 1824 3932
rect 1880 3876 1904 3932
rect 1960 3876 3184 3932
rect 3240 3876 3264 3932
rect 3320 3876 3344 3932
rect 3400 3876 3424 3932
rect 3480 3876 4280 3932
rect 44 3852 4280 3876
rect 44 3796 144 3852
rect 200 3796 224 3852
rect 280 3796 304 3852
rect 360 3796 384 3852
rect 440 3796 1664 3852
rect 1720 3796 1744 3852
rect 1800 3796 1824 3852
rect 1880 3796 1904 3852
rect 1960 3796 3184 3852
rect 3240 3796 3264 3852
rect 3320 3796 3344 3852
rect 3400 3796 3424 3852
rect 3480 3796 4280 3852
rect 44 3772 4280 3796
rect 44 3716 144 3772
rect 200 3716 224 3772
rect 280 3716 304 3772
rect 360 3716 384 3772
rect 440 3716 1664 3772
rect 1720 3716 1744 3772
rect 1800 3716 1824 3772
rect 1880 3716 1904 3772
rect 1960 3716 3184 3772
rect 3240 3716 3264 3772
rect 3320 3716 3344 3772
rect 3400 3716 3424 3772
rect 3480 3716 4280 3772
rect 44 3692 4280 3716
rect 44 3636 144 3692
rect 200 3636 224 3692
rect 280 3636 304 3692
rect 360 3636 384 3692
rect 440 3636 1664 3692
rect 1720 3636 1744 3692
rect 1800 3636 1824 3692
rect 1880 3636 1904 3692
rect 1960 3636 3184 3692
rect 3240 3636 3264 3692
rect 3320 3636 3344 3692
rect 3400 3636 3424 3692
rect 3480 3636 4280 3692
rect 44 3624 4280 3636
rect 44 3132 4280 3144
rect 44 3076 864 3132
rect 920 3076 944 3132
rect 1000 3076 1024 3132
rect 1080 3076 1104 3132
rect 1160 3076 2384 3132
rect 2440 3076 2464 3132
rect 2520 3076 2544 3132
rect 2600 3076 2624 3132
rect 2680 3076 3904 3132
rect 3960 3076 3984 3132
rect 4040 3076 4064 3132
rect 4120 3076 4144 3132
rect 4200 3076 4280 3132
rect 44 3052 4280 3076
rect 44 2996 864 3052
rect 920 2996 944 3052
rect 1000 2996 1024 3052
rect 1080 2996 1104 3052
rect 1160 2996 2384 3052
rect 2440 2996 2464 3052
rect 2520 2996 2544 3052
rect 2600 2996 2624 3052
rect 2680 2996 3904 3052
rect 3960 2996 3984 3052
rect 4040 2996 4064 3052
rect 4120 2996 4144 3052
rect 4200 2996 4280 3052
rect 44 2972 4280 2996
rect 44 2916 864 2972
rect 920 2916 944 2972
rect 1000 2916 1024 2972
rect 1080 2916 1104 2972
rect 1160 2916 2384 2972
rect 2440 2916 2464 2972
rect 2520 2916 2544 2972
rect 2600 2916 2624 2972
rect 2680 2916 3904 2972
rect 3960 2916 3984 2972
rect 4040 2916 4064 2972
rect 4120 2916 4144 2972
rect 4200 2916 4280 2972
rect 44 2892 4280 2916
rect 44 2836 864 2892
rect 920 2836 944 2892
rect 1000 2836 1024 2892
rect 1080 2836 1104 2892
rect 1160 2836 2384 2892
rect 2440 2836 2464 2892
rect 2520 2836 2544 2892
rect 2600 2836 2624 2892
rect 2680 2836 3904 2892
rect 3960 2836 3984 2892
rect 4040 2836 4064 2892
rect 4120 2836 4144 2892
rect 4200 2836 4280 2892
rect 44 2824 4280 2836
rect 44 2412 4280 2424
rect 44 2356 144 2412
rect 200 2356 224 2412
rect 280 2356 304 2412
rect 360 2356 384 2412
rect 440 2356 1664 2412
rect 1720 2356 1744 2412
rect 1800 2356 1824 2412
rect 1880 2356 1904 2412
rect 1960 2356 3184 2412
rect 3240 2356 3264 2412
rect 3320 2356 3344 2412
rect 3400 2356 3424 2412
rect 3480 2356 4280 2412
rect 44 2332 4280 2356
rect 44 2276 144 2332
rect 200 2276 224 2332
rect 280 2276 304 2332
rect 360 2276 384 2332
rect 440 2276 1664 2332
rect 1720 2276 1744 2332
rect 1800 2276 1824 2332
rect 1880 2276 1904 2332
rect 1960 2276 3184 2332
rect 3240 2276 3264 2332
rect 3320 2276 3344 2332
rect 3400 2276 3424 2332
rect 3480 2276 4280 2332
rect 44 2252 4280 2276
rect 44 2196 144 2252
rect 200 2196 224 2252
rect 280 2196 304 2252
rect 360 2196 384 2252
rect 440 2196 1664 2252
rect 1720 2196 1744 2252
rect 1800 2196 1824 2252
rect 1880 2196 1904 2252
rect 1960 2196 3184 2252
rect 3240 2196 3264 2252
rect 3320 2196 3344 2252
rect 3400 2196 3424 2252
rect 3480 2196 4280 2252
rect 44 2172 4280 2196
rect 44 2116 144 2172
rect 200 2116 224 2172
rect 280 2116 304 2172
rect 360 2116 384 2172
rect 440 2116 1664 2172
rect 1720 2116 1744 2172
rect 1800 2116 1824 2172
rect 1880 2116 1904 2172
rect 1960 2116 3184 2172
rect 3240 2116 3264 2172
rect 3320 2116 3344 2172
rect 3400 2116 3424 2172
rect 3480 2116 4280 2172
rect 44 2104 4280 2116
rect 44 1612 4280 1624
rect 44 1556 864 1612
rect 920 1556 944 1612
rect 1000 1556 1024 1612
rect 1080 1556 1104 1612
rect 1160 1556 2384 1612
rect 2440 1556 2464 1612
rect 2520 1556 2544 1612
rect 2600 1556 2624 1612
rect 2680 1556 3904 1612
rect 3960 1556 3984 1612
rect 4040 1556 4064 1612
rect 4120 1556 4144 1612
rect 4200 1556 4280 1612
rect 44 1532 4280 1556
rect 44 1476 864 1532
rect 920 1476 944 1532
rect 1000 1476 1024 1532
rect 1080 1476 1104 1532
rect 1160 1476 2384 1532
rect 2440 1476 2464 1532
rect 2520 1476 2544 1532
rect 2600 1476 2624 1532
rect 2680 1476 3904 1532
rect 3960 1476 3984 1532
rect 4040 1476 4064 1532
rect 4120 1476 4144 1532
rect 4200 1476 4280 1532
rect 44 1452 4280 1476
rect 44 1396 864 1452
rect 920 1396 944 1452
rect 1000 1396 1024 1452
rect 1080 1396 1104 1452
rect 1160 1396 2384 1452
rect 2440 1396 2464 1452
rect 2520 1396 2544 1452
rect 2600 1396 2624 1452
rect 2680 1396 3904 1452
rect 3960 1396 3984 1452
rect 4040 1396 4064 1452
rect 4120 1396 4144 1452
rect 4200 1396 4280 1452
rect 44 1372 4280 1396
rect 44 1316 864 1372
rect 920 1316 944 1372
rect 1000 1316 1024 1372
rect 1080 1316 1104 1372
rect 1160 1316 2384 1372
rect 2440 1316 2464 1372
rect 2520 1316 2544 1372
rect 2600 1316 2624 1372
rect 2680 1316 3904 1372
rect 3960 1316 3984 1372
rect 4040 1316 4064 1372
rect 4120 1316 4144 1372
rect 4200 1316 4280 1372
rect 44 1304 4280 1316
rect 44 892 4280 904
rect 44 836 144 892
rect 200 836 224 892
rect 280 836 304 892
rect 360 836 384 892
rect 440 836 1664 892
rect 1720 836 1744 892
rect 1800 836 1824 892
rect 1880 836 1904 892
rect 1960 836 3184 892
rect 3240 836 3264 892
rect 3320 836 3344 892
rect 3400 836 3424 892
rect 3480 836 4280 892
rect 44 812 4280 836
rect 44 756 144 812
rect 200 756 224 812
rect 280 756 304 812
rect 360 756 384 812
rect 440 756 1664 812
rect 1720 756 1744 812
rect 1800 756 1824 812
rect 1880 756 1904 812
rect 1960 756 3184 812
rect 3240 756 3264 812
rect 3320 756 3344 812
rect 3400 756 3424 812
rect 3480 756 4280 812
rect 44 732 4280 756
rect 44 676 144 732
rect 200 676 224 732
rect 280 676 304 732
rect 360 676 384 732
rect 440 676 1664 732
rect 1720 676 1744 732
rect 1800 676 1824 732
rect 1880 676 1904 732
rect 1960 676 3184 732
rect 3240 676 3264 732
rect 3320 676 3344 732
rect 3400 676 3424 732
rect 3480 676 4280 732
rect 44 652 4280 676
rect 44 596 144 652
rect 200 596 224 652
rect 280 596 304 652
rect 360 596 384 652
rect 440 596 1664 652
rect 1720 596 1744 652
rect 1800 596 1824 652
rect 1880 596 1904 652
rect 1960 596 3184 652
rect 3240 596 3264 652
rect 3320 596 3344 652
rect 3400 596 3424 652
rect 3480 596 4280 652
rect 44 584 4280 596
use sky130_fd_sc_hd__decap_4  FILLER_0_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 368 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 920 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15
timestamp 1673029049
transform 1 0 1472 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17
timestamp 1673029049
transform 1 0 1656 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp 1673029049
transform 1 0 2208 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25
timestamp 1673029049
transform 1 0 2392 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31
timestamp 1673029049
transform 1 0 2944 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33
timestamp 1673029049
transform 1 0 3128 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39
timestamp 1673029049
transform 1 0 3680 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1673029049
transform 1 0 3864 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 368 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1472 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1673029049
transform 1 0 1748 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1673029049
transform 1 0 2852 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_35
timestamp 1673029049
transform 1 0 3312 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_41
timestamp 1673029049
transform 1 0 3864 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1673029049
transform 1 0 368 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1673029049
transform 1 0 736 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1673029049
transform 1 0 920 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_21
timestamp 1673029049
transform 1 0 2024 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_26
timestamp 1673029049
transform 1 0 2484 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1673029049
transform 1 0 3588 0 1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1673029049
transform 1 0 368 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1673029049
transform 1 0 1472 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_18
timestamp 1673029049
transform 1 0 1748 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_24
timestamp 1673029049
transform 1 0 2300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_28
timestamp 1673029049
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35
timestamp 1673029049
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1673029049
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1673029049
transform 1 0 368 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1673029049
transform 1 0 736 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1673029049
transform 1 0 920 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_21
timestamp 1673029049
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_26
timestamp 1673029049
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1673029049
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1673029049
transform 1 0 368 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1673029049
transform 1 0 736 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_9
timestamp 1673029049
transform 1 0 920 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1673029049
transform 1 0 1472 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_17
timestamp 1673029049
transform 1 0 1656 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1673029049
transform 1 0 2208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_25
timestamp 1673029049
transform 1 0 2392 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1673029049
transform 1 0 2944 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_33
timestamp 1673029049
transform 1 0 3128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp 1673029049
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_41
timestamp 1673029049
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 92 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 4232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 92 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 4232 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 92 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 4232 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 92 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 92 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 92 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 4232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1673029049
transform 1 0 1564 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1673029049
transform 1 0 2300 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1673029049
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1673029049
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1673029049
transform 1 0 1656 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1673029049
transform 1 0 3220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1673029049
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1673029049
transform 1 0 2392 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1673029049
transform 1 0 1656 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1673029049
transform 1 0 3220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1673029049
transform 1 0 828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1673029049
transform 1 0 2392 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1673029049
transform 1 0 828 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1673029049
transform 1 0 1564 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1673029049
transform 1 0 2300 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1673029049
transform 1 0 3036 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1673029049
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2392 0 -1 2720
box -38 -48 314 592
<< labels >>
flabel metal2 s 2134 0 2190 400 0 FreeSans 224 90 0 0 gpio_logic1
port 0 nsew signal tristate
flabel metal2 s 132 496 452 3944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 1652 496 1972 3944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 3172 496 3492 3944 0 FreeSans 1792 90 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 44 584 4280 904 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 44 2104 4280 2424 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal3 s 44 3624 4280 3944 0 FreeSans 1920 0 0 0 vccd1
port 1 nsew power bidirectional
flabel metal2 s 852 496 1172 3856 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 2372 496 2692 3856 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal2 s 3892 496 4212 3856 0 FreeSans 1792 90 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 44 1304 4280 1624 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
flabel metal3 s 44 2824 4280 3144 0 FreeSans 1920 0 0 0 vssd1
port 2 nsew ground bidirectional
rlabel metal1 2162 3264 2162 3264 0 vccd1
rlabel metal1 2162 3808 2162 3808 0 vssd1
rlabel metal2 2162 1384 2162 1384 0 gpio_logic1
<< properties >>
string FIXED_BBOX 0 0 4400 4400
<< end >>
