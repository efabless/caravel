magic
tech sky130A
magscale 1 2
timestamp 1699123252
<< viali >>
rect 7205 13481 7239 13515
rect 10701 13481 10735 13515
rect 11161 13481 11195 13515
rect 16405 13481 16439 13515
rect 2973 13413 3007 13447
rect 1501 13345 1535 13379
rect 4445 13345 4479 13379
rect 7573 13345 7607 13379
rect 8493 13345 8527 13379
rect 9505 13345 9539 13379
rect 15117 13345 15151 13379
rect 17693 13345 17727 13379
rect 3249 13277 3283 13311
rect 4997 13277 5031 13311
rect 6469 13277 6503 13311
rect 7941 13277 7975 13311
rect 9770 13255 9804 13289
rect 9965 13277 9999 13311
rect 10425 13277 10459 13311
rect 11253 13277 11287 13311
rect 11621 13277 11655 13311
rect 12633 13277 12667 13311
rect 12817 13277 12851 13311
rect 13737 13277 13771 13311
rect 14381 13277 14415 13311
rect 14565 13277 14599 13311
rect 14933 13277 14967 13311
rect 15577 13277 15611 13311
rect 16773 13277 16807 13311
rect 17141 13277 17175 13311
rect 18061 13277 18095 13311
rect 3893 13209 3927 13243
rect 3985 13209 4019 13243
rect 5457 13209 5491 13243
rect 5549 13209 5583 13243
rect 5825 13209 5859 13243
rect 8401 13209 8435 13243
rect 9321 13209 9355 13243
rect 9873 13209 9907 13243
rect 12081 13209 12115 13243
rect 12173 13209 12207 13243
rect 13185 13209 13219 13243
rect 15853 13209 15887 13243
rect 17601 13209 17635 13243
rect 1869 13141 1903 13175
rect 2513 13141 2547 13175
rect 3433 13141 3467 13175
rect 6009 13141 6043 13175
rect 6653 13141 6687 13175
rect 7665 13141 7699 13175
rect 12633 13141 12667 13175
rect 13093 13141 13127 13175
rect 13553 13141 13587 13175
rect 14381 13141 14415 13175
rect 15393 13141 15427 13175
rect 15945 13141 15979 13175
rect 17969 13141 18003 13175
rect 3065 12869 3099 12903
rect 4169 12869 4203 12903
rect 6101 12869 6135 12903
rect 8953 12869 8987 12903
rect 12725 12869 12759 12903
rect 13829 12869 13863 12903
rect 13921 12869 13955 12903
rect 15209 12869 15243 12903
rect 16221 12869 16255 12903
rect 17417 12869 17451 12903
rect 18245 12869 18279 12903
rect 2513 12801 2547 12835
rect 2789 12801 2823 12835
rect 3709 12801 3743 12835
rect 4537 12801 4571 12835
rect 6009 12801 6043 12835
rect 6469 12801 6503 12835
rect 6929 12801 6963 12835
rect 7389 12801 7423 12835
rect 8861 12801 8895 12835
rect 9413 12801 9447 12835
rect 9695 12801 9729 12835
rect 10609 12801 10643 12835
rect 11989 12801 12023 12835
rect 12909 12801 12943 12835
rect 13645 12801 13679 12835
rect 14473 12801 14507 12835
rect 15393 12801 15427 12835
rect 16773 12801 16807 12835
rect 17693 12801 17727 12835
rect 18061 12801 18095 12835
rect 11253 12733 11287 12767
rect 15669 12733 15703 12767
rect 16129 12733 16163 12767
rect 2421 12665 2455 12699
rect 11713 12665 11747 12699
rect 1685 12597 1719 12631
rect 2053 12597 2087 12631
rect 4077 12597 4111 12631
rect 6561 12597 6595 12631
rect 7021 12597 7055 12631
rect 9229 12597 9263 12631
rect 13369 12597 13403 12631
rect 5089 12393 5123 12427
rect 9229 12393 9263 12427
rect 13185 12393 13219 12427
rect 17693 12325 17727 12359
rect 4537 12257 4571 12291
rect 4721 12257 4755 12291
rect 7297 12257 7331 12291
rect 9965 12257 9999 12291
rect 12173 12257 12207 12291
rect 12725 12257 12759 12291
rect 15209 12257 15243 12291
rect 17325 12257 17359 12291
rect 1685 12189 1719 12223
rect 1869 12189 1903 12223
rect 2973 12189 3007 12223
rect 3341 12189 3375 12223
rect 5549 12189 5583 12223
rect 6469 12189 6503 12223
rect 6745 12189 6779 12223
rect 7665 12189 7699 12223
rect 8309 12189 8343 12223
rect 9143 12189 9177 12223
rect 9321 12189 9355 12223
rect 10793 12189 10827 12223
rect 11253 12189 11287 12223
rect 11437 12189 11471 12223
rect 12633 12189 12667 12223
rect 13082 12167 13116 12201
rect 13461 12189 13495 12223
rect 13553 12189 13587 12223
rect 14197 12189 14231 12223
rect 14289 12189 14323 12223
rect 14657 12189 14691 12223
rect 15117 12189 15151 12223
rect 15761 12189 15795 12223
rect 16681 12189 16715 12223
rect 18153 12189 18187 12223
rect 3985 12121 4019 12155
rect 4169 12121 4203 12155
rect 4629 12121 4663 12155
rect 5825 12121 5859 12155
rect 6837 12121 6871 12155
rect 8585 12121 8619 12155
rect 10149 12121 10183 12155
rect 11713 12121 11747 12155
rect 11805 12121 11839 12155
rect 17601 12121 17635 12155
rect 1685 12053 1719 12087
rect 2421 12053 2455 12087
rect 2881 12053 2915 12087
rect 3433 12053 3467 12087
rect 10057 12053 10091 12087
rect 10517 12053 10551 12087
rect 10977 12053 11011 12087
rect 4261 11849 4295 11883
rect 6009 11849 6043 11883
rect 8861 11849 8895 11883
rect 9413 11849 9447 11883
rect 11621 11849 11655 11883
rect 13093 11849 13127 11883
rect 14013 11849 14047 11883
rect 15853 11849 15887 11883
rect 2053 11781 2087 11815
rect 8309 11781 8343 11815
rect 8401 11781 8435 11815
rect 10333 11781 10367 11815
rect 11161 11781 11195 11815
rect 18429 11781 18463 11815
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 2421 11713 2455 11747
rect 3893 11713 3927 11747
rect 4445 11713 4479 11747
rect 5457 11713 5491 11747
rect 5917 11713 5951 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 7381 11719 7415 11753
rect 7573 11713 7607 11747
rect 8861 11713 8895 11747
rect 9045 11713 9079 11747
rect 9321 11713 9355 11747
rect 9965 11713 9999 11747
rect 10793 11713 10827 11747
rect 11253 11713 11287 11747
rect 11989 11713 12023 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 14013 11713 14047 11747
rect 14197 11703 14231 11737
rect 14473 11713 14507 11747
rect 15485 11713 15519 11747
rect 16129 11713 16163 11747
rect 16865 11713 16899 11747
rect 17785 11713 17819 11747
rect 4997 11645 5031 11679
rect 5549 11645 5583 11679
rect 6653 11645 6687 11679
rect 7481 11645 7515 11679
rect 7849 11645 7883 11679
rect 9781 11645 9815 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 15209 11645 15243 11679
rect 15393 11645 15427 11679
rect 3709 11577 3743 11611
rect 10241 11577 10275 11611
rect 16221 11577 16255 11611
rect 7113 11509 7147 11543
rect 10701 11509 10735 11543
rect 12725 11509 12759 11543
rect 13645 11509 13679 11543
rect 14565 11509 14599 11543
rect 3985 11305 4019 11339
rect 6285 11305 6319 11339
rect 6653 11305 6687 11339
rect 8585 11305 8619 11339
rect 9413 11305 9447 11339
rect 10701 11305 10735 11339
rect 11529 11305 11563 11339
rect 15209 11305 15243 11339
rect 5825 11237 5859 11271
rect 14197 11237 14231 11271
rect 16129 11237 16163 11271
rect 16957 11237 16991 11271
rect 2329 11169 2363 11203
rect 2881 11169 2915 11203
rect 11161 11169 11195 11203
rect 13369 11169 13403 11203
rect 13461 11169 13495 11203
rect 17049 11169 17083 11203
rect 17877 11169 17911 11203
rect 1685 11101 1719 11135
rect 1869 11101 1903 11135
rect 4353 11101 4387 11135
rect 5549 11101 5583 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 7113 11101 7147 11135
rect 7297 11101 7331 11135
rect 8033 11101 8067 11135
rect 8493 11101 8527 11135
rect 8677 11101 8711 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9965 11101 9999 11135
rect 10149 11101 10183 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 12081 11101 12115 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 14322 11101 14356 11135
rect 14749 11101 14783 11135
rect 14841 11101 14875 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 15669 11101 15703 11135
rect 16037 11101 16071 11135
rect 16497 11101 16531 11135
rect 17325 11101 17359 11135
rect 18337 11101 18371 11135
rect 1777 11033 1811 11067
rect 2789 11033 2823 11067
rect 3341 11033 3375 11067
rect 7389 11033 7423 11067
rect 10057 11033 10091 11067
rect 12449 11033 12483 11067
rect 17785 11033 17819 11067
rect 3525 10965 3559 10999
rect 4077 10965 4111 10999
rect 7941 10965 7975 10999
rect 14381 10965 14415 10999
rect 18245 10965 18279 10999
rect 7573 10761 7607 10795
rect 9965 10761 9999 10795
rect 11161 10761 11195 10795
rect 12541 10761 12575 10795
rect 13001 10761 13035 10795
rect 14657 10761 14691 10795
rect 15025 10761 15059 10795
rect 16313 10761 16347 10795
rect 3341 10693 3375 10727
rect 4353 10693 4387 10727
rect 5181 10693 5215 10727
rect 6561 10693 6595 10727
rect 9321 10693 9355 10727
rect 12265 10693 12299 10727
rect 18337 10693 18371 10727
rect 1501 10625 1535 10659
rect 2053 10625 2087 10659
rect 2329 10625 2363 10659
rect 3985 10625 4019 10659
rect 4261 10625 4295 10659
rect 4721 10625 4755 10659
rect 5365 10625 5399 10659
rect 6101 10625 6135 10659
rect 7757 10625 7791 10659
rect 7849 10625 7883 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 11069 10625 11103 10659
rect 11253 10625 11287 10659
rect 11897 10625 11931 10659
rect 12909 10625 12943 10659
rect 13645 10625 13679 10659
rect 13737 10625 13771 10659
rect 14381 10625 14415 10659
rect 15393 10625 15427 10659
rect 15577 10625 15611 10659
rect 16037 10625 16071 10659
rect 16770 10625 16804 10659
rect 18245 10625 18279 10659
rect 2789 10557 2823 10591
rect 6469 10557 6503 10591
rect 7021 10557 7055 10591
rect 7573 10557 7607 10591
rect 11713 10557 11747 10591
rect 13185 10557 13219 10591
rect 14657 10557 14691 10591
rect 15485 10557 15519 10591
rect 2237 10489 2271 10523
rect 3249 10489 3283 10523
rect 4905 10489 4939 10523
rect 8125 10489 8159 10523
rect 8861 10489 8895 10523
rect 11897 10489 11931 10523
rect 1593 10421 1627 10455
rect 3709 10421 3743 10455
rect 14013 10421 14047 10455
rect 14473 10421 14507 10455
rect 15945 10421 15979 10455
rect 5549 10217 5583 10251
rect 8125 10217 8159 10251
rect 8585 10217 8619 10251
rect 9321 10217 9355 10251
rect 9873 10217 9907 10251
rect 13277 10217 13311 10251
rect 14381 10217 14415 10251
rect 18429 10217 18463 10251
rect 11345 10149 11379 10183
rect 1593 10081 1627 10115
rect 3525 10081 3559 10115
rect 6745 10081 6779 10115
rect 7481 10081 7515 10115
rect 10241 10081 10275 10115
rect 11713 10081 11747 10115
rect 14197 10081 14231 10115
rect 15761 10081 15795 10115
rect 1961 10013 1995 10047
rect 3433 10013 3467 10047
rect 4077 10013 4111 10047
rect 4813 10013 4847 10047
rect 5457 10013 5491 10047
rect 7389 10013 7423 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 8677 10013 8711 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 9781 10013 9815 10047
rect 10793 10013 10827 10047
rect 10970 10013 11004 10047
rect 11253 10013 11287 10047
rect 11897 10013 11931 10047
rect 12081 10013 12115 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13185 10013 13219 10047
rect 13645 10013 13679 10047
rect 14473 10013 14507 10047
rect 15301 10013 15335 10047
rect 15669 10013 15703 10047
rect 16037 10013 16071 10047
rect 16313 10013 16347 10047
rect 16957 10013 16991 10047
rect 17969 10013 18003 10047
rect 3893 9945 3927 9979
rect 6193 9945 6227 9979
rect 6285 9945 6319 9979
rect 7113 9945 7147 9979
rect 9965 9945 9999 9979
rect 10885 9945 10919 9979
rect 17233 9945 17267 9979
rect 12541 9877 12575 9911
rect 13737 9877 13771 9911
rect 14197 9877 14231 9911
rect 15025 9877 15059 9911
rect 17877 9877 17911 9911
rect 2605 9673 2639 9707
rect 4629 9673 4663 9707
rect 6101 9673 6135 9707
rect 1685 9605 1719 9639
rect 1869 9605 1903 9639
rect 6653 9605 6687 9639
rect 8953 9605 8987 9639
rect 9505 9605 9539 9639
rect 9965 9605 9999 9639
rect 10767 9605 10801 9639
rect 11621 9605 11655 9639
rect 13185 9605 13219 9639
rect 16129 9605 16163 9639
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 4813 9537 4847 9571
rect 5273 9537 5307 9571
rect 6469 9537 6503 9571
rect 7389 9537 7423 9571
rect 7757 9537 7791 9571
rect 8217 9537 8251 9571
rect 8861 9537 8895 9571
rect 9873 9537 9907 9571
rect 10057 9537 10091 9571
rect 10670 9537 10704 9571
rect 12357 9537 12391 9571
rect 13460 9537 13494 9571
rect 13553 9537 13587 9571
rect 14013 9537 14047 9571
rect 14565 9537 14599 9571
rect 15025 9537 15059 9571
rect 15209 9537 15243 9571
rect 15491 9537 15525 9571
rect 15669 9537 15703 9571
rect 16037 9537 16071 9571
rect 16221 9537 16255 9571
rect 17601 9537 17635 9571
rect 1593 9469 1627 9503
rect 3801 9469 3835 9503
rect 4261 9469 4295 9503
rect 4353 9469 4387 9503
rect 9137 9469 9171 9503
rect 11161 9469 11195 9503
rect 12449 9469 12483 9503
rect 12541 9469 12575 9503
rect 16773 9469 16807 9503
rect 17325 9469 17359 9503
rect 18153 9469 18187 9503
rect 5089 9401 5123 9435
rect 5641 9401 5675 9435
rect 10517 9401 10551 9435
rect 17233 9401 17267 9435
rect 18061 9401 18095 9435
rect 2145 9333 2179 9367
rect 6009 9333 6043 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 11069 9333 11103 9367
rect 11989 9333 12023 9367
rect 14105 9333 14139 9367
rect 15117 9333 15151 9367
rect 15577 9333 15611 9367
rect 7021 9129 7055 9163
rect 7941 9129 7975 9163
rect 9045 9129 9079 9163
rect 12817 9129 12851 9163
rect 14289 9129 14323 9163
rect 15485 9129 15519 9163
rect 18337 9129 18371 9163
rect 8585 9061 8619 9095
rect 15945 9061 15979 9095
rect 17693 9061 17727 9095
rect 9597 8993 9631 9027
rect 12081 8993 12115 9027
rect 1777 8925 1811 8959
rect 3249 8925 3283 8959
rect 4813 8925 4847 8959
rect 5825 8925 5859 8959
rect 6745 8925 6779 8959
rect 7205 8925 7239 8959
rect 7849 8925 7883 8959
rect 8033 8925 8067 8959
rect 8493 8925 8527 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 11345 8925 11379 8959
rect 12265 8925 12299 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 13553 8925 13587 8959
rect 13737 8925 13771 8959
rect 14197 8925 14231 8959
rect 14841 8925 14875 8959
rect 15393 8925 15427 8959
rect 15577 8925 15611 8959
rect 15853 8925 15887 8959
rect 16405 8925 16439 8959
rect 17877 8925 17911 8959
rect 18245 8925 18279 8959
rect 3341 8857 3375 8891
rect 3893 8857 3927 8891
rect 4077 8857 4111 8891
rect 5181 8857 5215 8891
rect 10609 8857 10643 8891
rect 11897 8857 11931 8891
rect 11989 8857 12023 8891
rect 14749 8857 14783 8891
rect 9413 8789 9447 8823
rect 9505 8789 9539 8823
rect 11161 8789 11195 8823
rect 13553 8789 13587 8823
rect 7389 8585 7423 8619
rect 11713 8585 11747 8619
rect 13737 8585 13771 8619
rect 18153 8585 18187 8619
rect 2697 8517 2731 8551
rect 3249 8517 3283 8551
rect 4169 8517 4203 8551
rect 6469 8517 6503 8551
rect 9597 8517 9631 8551
rect 11069 8517 11103 8551
rect 17693 8517 17727 8551
rect 1777 8449 1811 8483
rect 2237 8449 2271 8483
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 3617 8449 3651 8483
rect 4077 8449 4111 8483
rect 4629 8449 4663 8483
rect 5917 8449 5951 8483
rect 7021 8449 7055 8483
rect 7481 8449 7515 8483
rect 8493 8449 8527 8483
rect 9413 8449 9447 8483
rect 10333 8449 10367 8483
rect 11161 8449 11195 8483
rect 11989 8449 12023 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 13001 8449 13035 8483
rect 13093 8449 13127 8483
rect 13645 8449 13679 8483
rect 13829 8449 13863 8483
rect 14197 8449 14231 8483
rect 14565 8449 14599 8483
rect 15025 8449 15059 8483
rect 15209 8449 15243 8483
rect 15945 8449 15979 8483
rect 16129 8449 16163 8483
rect 16957 8449 16991 8483
rect 17877 8449 17911 8483
rect 18337 8449 18371 8483
rect 6561 8381 6595 8415
rect 7849 8381 7883 8415
rect 9045 8381 9079 8415
rect 10609 8381 10643 8415
rect 12817 8381 12851 8415
rect 14381 8381 14415 8415
rect 1869 8313 1903 8347
rect 4445 8313 4479 8347
rect 8953 8313 8987 8347
rect 12265 8313 12299 8347
rect 14473 8313 14507 8347
rect 15577 8313 15611 8347
rect 5733 8245 5767 8279
rect 15117 8245 15151 8279
rect 16129 8245 16163 8279
rect 1593 8041 1627 8075
rect 1961 8041 1995 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 6377 8041 6411 8075
rect 9505 8041 9539 8075
rect 12817 8041 12851 8075
rect 13369 8041 13403 8075
rect 17417 8041 17451 8075
rect 18245 8041 18279 8075
rect 3157 7973 3191 8007
rect 7665 7905 7699 7939
rect 13553 7905 13587 7939
rect 17601 7905 17635 7939
rect 4353 7837 4387 7871
rect 5733 7837 5767 7871
rect 6377 7837 6411 7871
rect 6745 7837 6779 7871
rect 7389 7837 7423 7871
rect 8217 7837 8251 7871
rect 8401 7837 8435 7871
rect 10241 7837 10275 7871
rect 10333 7837 10367 7871
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 11621 7837 11655 7871
rect 11805 7827 11839 7861
rect 12173 7837 12207 7871
rect 12449 7837 12483 7871
rect 12725 7837 12759 7871
rect 13277 7837 13311 7871
rect 14197 7837 14231 7871
rect 16497 7837 16531 7871
rect 17693 7837 17727 7871
rect 18337 7837 18371 7871
rect 6101 7769 6135 7803
rect 7481 7769 7515 7803
rect 8033 7769 8067 7803
rect 9597 7769 9631 7803
rect 13553 7769 13587 7803
rect 14473 7769 14507 7803
rect 16221 7769 16255 7803
rect 4261 7701 4295 7735
rect 7021 7701 7055 7735
rect 11621 7701 11655 7735
rect 12173 7701 12207 7735
rect 16589 7701 16623 7735
rect 17049 7701 17083 7735
rect 12081 7497 12115 7531
rect 15577 7497 15611 7531
rect 18061 7497 18095 7531
rect 10793 7429 10827 7463
rect 16037 7429 16071 7463
rect 16865 7429 16899 7463
rect 1961 7361 1995 7395
rect 2881 7361 2915 7395
rect 5181 7361 5215 7395
rect 5365 7361 5399 7395
rect 6101 7361 6135 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 9137 7361 9171 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12633 7361 12667 7395
rect 13185 7361 13219 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 16129 7361 16163 7395
rect 16773 7361 16807 7395
rect 16957 7361 16991 7395
rect 17417 7361 17451 7395
rect 17601 7361 17635 7395
rect 18245 7361 18279 7395
rect 2513 7293 2547 7327
rect 3157 7293 3191 7327
rect 13461 7293 13495 7327
rect 15209 7293 15243 7327
rect 5917 7225 5951 7259
rect 8953 7225 8987 7259
rect 4629 7157 4663 7191
rect 5273 7157 5307 7191
rect 6653 7157 6687 7191
rect 7205 7157 7239 7191
rect 10701 7157 10735 7191
rect 12725 7157 12759 7191
rect 17509 7157 17543 7191
rect 1961 6953 1995 6987
rect 3985 6953 4019 6987
rect 4077 6953 4111 6987
rect 6916 6953 6950 6987
rect 13277 6953 13311 6987
rect 15025 6953 15059 6987
rect 16865 6953 16899 6987
rect 4997 6885 5031 6919
rect 13185 6885 13219 6919
rect 17785 6885 17819 6919
rect 2605 6817 2639 6851
rect 2789 6817 2823 6851
rect 3893 6817 3927 6851
rect 6285 6817 6319 6851
rect 6653 6817 6687 6851
rect 10149 6817 10183 6851
rect 11897 6817 11931 6851
rect 12725 6817 12759 6851
rect 13369 6817 13403 6851
rect 14473 6817 14507 6851
rect 16957 6817 16991 6851
rect 18061 6817 18095 6851
rect 2145 6749 2179 6783
rect 2881 6749 2915 6783
rect 4169 6749 4203 6783
rect 4905 6749 4939 6783
rect 5089 6751 5123 6785
rect 5733 6749 5767 6783
rect 9781 6749 9815 6783
rect 10333 6749 10367 6783
rect 10517 6749 10551 6783
rect 10793 6749 10827 6783
rect 10977 6749 11011 6783
rect 11989 6749 12023 6783
rect 12633 6751 12667 6785
rect 12817 6749 12851 6783
rect 13093 6749 13127 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 15117 6749 15151 6783
rect 15393 6749 15427 6783
rect 15577 6749 15611 6783
rect 16681 6749 16715 6783
rect 16773 6749 16807 6783
rect 18153 6749 18187 6783
rect 4537 6681 4571 6715
rect 10885 6681 10919 6715
rect 2605 6613 2639 6647
rect 5365 6613 5399 6647
rect 8401 6613 8435 6647
rect 9045 6613 9079 6647
rect 9689 6613 9723 6647
rect 15485 6613 15519 6647
rect 3617 6409 3651 6443
rect 16313 6409 16347 6443
rect 17417 6409 17451 6443
rect 1777 6341 1811 6375
rect 5825 6341 5859 6375
rect 7205 6341 7239 6375
rect 11897 6341 11931 6375
rect 13645 6341 13679 6375
rect 14749 6341 14783 6375
rect 5641 6273 5675 6307
rect 6469 6273 6503 6307
rect 6653 6273 6687 6307
rect 7389 6273 7423 6307
rect 7481 6273 7515 6307
rect 7849 6273 7883 6307
rect 8585 6273 8619 6307
rect 9045 6273 9079 6307
rect 9229 6273 9263 6307
rect 9413 6273 9447 6307
rect 9965 6273 9999 6307
rect 10425 6273 10459 6307
rect 10793 6273 10827 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 15301 6273 15335 6307
rect 15485 6273 15519 6307
rect 16129 6273 16163 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 1501 6205 1535 6239
rect 5917 6205 5951 6239
rect 10287 6205 10321 6239
rect 11621 6205 11655 6239
rect 15945 6205 15979 6239
rect 17417 6205 17451 6239
rect 4261 6137 4295 6171
rect 5273 6137 5307 6171
rect 7205 6137 7239 6171
rect 3249 6069 3283 6103
rect 3893 6069 3927 6103
rect 6653 6069 6687 6103
rect 10057 6069 10091 6103
rect 10149 6069 10183 6103
rect 10977 6069 11011 6103
rect 15393 6069 15427 6103
rect 17601 6069 17635 6103
rect 18061 6069 18095 6103
rect 1777 5865 1811 5899
rect 6377 5865 6411 5899
rect 7021 5865 7055 5899
rect 7849 5865 7883 5899
rect 9137 5865 9171 5899
rect 10149 5865 10183 5899
rect 11713 5865 11747 5899
rect 11805 5865 11839 5899
rect 16681 5865 16715 5899
rect 2513 5797 2547 5831
rect 4169 5797 4203 5831
rect 15485 5797 15519 5831
rect 4813 5729 4847 5763
rect 5273 5729 5307 5763
rect 11897 5729 11931 5763
rect 12725 5729 12759 5763
rect 17693 5729 17727 5763
rect 17969 5729 18003 5763
rect 1685 5661 1719 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 4905 5661 4939 5695
rect 6653 5661 6687 5695
rect 6929 5661 6963 5695
rect 7113 5661 7147 5695
rect 7573 5661 7607 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 9045 5661 9079 5695
rect 9689 5661 9723 5695
rect 9873 5661 9907 5695
rect 10149 5661 10183 5695
rect 11621 5661 11655 5695
rect 12633 5661 12667 5695
rect 12817 5661 12851 5695
rect 13277 5661 13311 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 16589 5661 16623 5695
rect 18061 5661 18095 5695
rect 6377 5593 6411 5627
rect 7849 5593 7883 5627
rect 10241 5593 10275 5627
rect 10425 5593 10459 5627
rect 16037 5593 16071 5627
rect 2145 5525 2179 5559
rect 3525 5525 3559 5559
rect 6561 5525 6595 5559
rect 7665 5525 7699 5559
rect 8125 5525 8159 5559
rect 9873 5525 9907 5559
rect 13185 5525 13219 5559
rect 1869 5321 1903 5355
rect 2973 5321 3007 5355
rect 5549 5321 5583 5355
rect 9137 5321 9171 5355
rect 16221 5321 16255 5355
rect 17601 5321 17635 5355
rect 2237 5253 2271 5287
rect 6009 5253 6043 5287
rect 7665 5253 7699 5287
rect 10057 5253 10091 5287
rect 15393 5253 15427 5287
rect 1777 5185 1811 5219
rect 3065 5185 3099 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4721 5185 4755 5219
rect 5365 5185 5399 5219
rect 6101 5185 6135 5219
rect 6929 5185 6963 5219
rect 7113 5185 7147 5219
rect 9781 5185 9815 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 10977 5185 11011 5219
rect 11622 5175 11656 5209
rect 12449 5185 12483 5219
rect 12633 5185 12667 5219
rect 13369 5185 13403 5219
rect 15945 5185 15979 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 17417 5185 17451 5219
rect 17601 5185 17635 5219
rect 5181 5117 5215 5151
rect 7389 5117 7423 5151
rect 9689 5117 9723 5151
rect 11897 5117 11931 5151
rect 13645 5117 13679 5151
rect 15761 5117 15795 5151
rect 16313 5117 16347 5151
rect 10333 5049 10367 5083
rect 4077 4981 4111 5015
rect 4813 4981 4847 5015
rect 6929 4981 6963 5015
rect 10609 4981 10643 5015
rect 11069 4981 11103 5015
rect 11713 4981 11747 5015
rect 11805 4981 11839 5015
rect 12633 4981 12667 5015
rect 16865 4981 16899 5015
rect 1593 4777 1627 4811
rect 6285 4777 6319 4811
rect 7297 4777 7331 4811
rect 8493 4777 8527 4811
rect 9137 4777 9171 4811
rect 10627 4777 10661 4811
rect 13369 4777 13403 4811
rect 13461 4777 13495 4811
rect 4445 4709 4479 4743
rect 3985 4641 4019 4675
rect 5549 4641 5583 4675
rect 7113 4641 7147 4675
rect 8033 4641 8067 4675
rect 10885 4641 10919 4675
rect 11897 4641 11931 4675
rect 12173 4641 12207 4675
rect 13553 4641 13587 4675
rect 14473 4641 14507 4675
rect 17325 4641 17359 4675
rect 17969 4641 18003 4675
rect 2789 4573 2823 4607
rect 3249 4573 3283 4607
rect 3433 4573 3467 4607
rect 4077 4573 4111 4607
rect 5733 4573 5767 4607
rect 5825 4573 5859 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 6994 4573 7028 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8585 4573 8619 4607
rect 11345 4573 11379 4607
rect 11805 4573 11839 4607
rect 13277 4573 13311 4607
rect 14381 4573 14415 4607
rect 14565 4573 14599 4607
rect 14841 4573 14875 4607
rect 15025 4573 15059 4607
rect 15577 4573 15611 4607
rect 15761 4573 15795 4607
rect 17417 4573 17451 4607
rect 17877 4573 17911 4607
rect 18061 4573 18095 4607
rect 5549 4505 5583 4539
rect 2697 4437 2731 4471
rect 3249 4437 3283 4471
rect 11253 4437 11287 4471
rect 14933 4437 14967 4471
rect 15669 4437 15703 4471
rect 17049 4437 17083 4471
rect 3617 4233 3651 4267
rect 11161 4233 11195 4267
rect 7849 4165 7883 4199
rect 12449 4165 12483 4199
rect 13461 4165 13495 4199
rect 5273 4097 5307 4131
rect 5365 4097 5399 4131
rect 5549 4097 5583 4131
rect 6469 4097 6503 4131
rect 6653 4097 6687 4131
rect 7481 4097 7515 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 9321 4097 9355 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 11069 4097 11103 4131
rect 11897 4097 11931 4131
rect 12081 4097 12115 4131
rect 12357 4097 12391 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 13369 4097 13403 4131
rect 13553 4097 13587 4131
rect 14105 4097 14139 4131
rect 14565 4097 14599 4131
rect 14749 4097 14783 4131
rect 15485 4097 15519 4131
rect 16773 4097 16807 4131
rect 16957 4097 16991 4131
rect 1501 4029 1535 4063
rect 1777 4029 1811 4063
rect 3249 4029 3283 4063
rect 6837 4029 6871 4063
rect 7389 4029 7423 4063
rect 7757 4029 7791 4063
rect 10793 4029 10827 4063
rect 14657 4029 14691 4063
rect 15761 4029 15795 4063
rect 16865 4029 16899 4063
rect 4629 3961 4663 3995
rect 5549 3961 5583 3995
rect 14197 3961 14231 3995
rect 15577 3961 15611 3995
rect 15669 3961 15703 3995
rect 4997 3893 5031 3927
rect 7205 3893 7239 3927
rect 10701 3893 10735 3927
rect 13001 3893 13035 3927
rect 2789 3689 2823 3723
rect 8493 3689 8527 3723
rect 9321 3689 9355 3723
rect 9689 3689 9723 3723
rect 11805 3689 11839 3723
rect 16405 3689 16439 3723
rect 16957 3689 16991 3723
rect 1869 3621 1903 3655
rect 2881 3553 2915 3587
rect 5365 3553 5399 3587
rect 5825 3553 5859 3587
rect 7021 3553 7055 3587
rect 11161 3553 11195 3587
rect 11437 3553 11471 3587
rect 13185 3553 13219 3587
rect 14473 3553 14507 3587
rect 15393 3553 15427 3587
rect 15669 3553 15703 3587
rect 1777 3485 1811 3519
rect 2237 3485 2271 3519
rect 2605 3485 2639 3519
rect 2697 3485 2731 3519
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 5733 3485 5767 3519
rect 6745 3485 6779 3519
rect 11713 3485 11747 3519
rect 11897 3485 11931 3519
rect 12633 3485 12667 3519
rect 12909 3485 12943 3519
rect 13001 3485 13035 3519
rect 13737 3485 13771 3519
rect 13829 3485 13863 3519
rect 14381 3485 14415 3519
rect 14565 3485 14599 3519
rect 15761 3485 15795 3519
rect 16405 3485 16439 3519
rect 16589 3485 16623 3519
rect 16865 3485 16899 3519
rect 3341 3417 3375 3451
rect 12357 3417 12391 3451
rect 4353 3349 4387 3383
rect 13185 3349 13219 3383
rect 5089 3145 5123 3179
rect 7849 3145 7883 3179
rect 8769 3145 8803 3179
rect 10149 3145 10183 3179
rect 10885 3145 10919 3179
rect 11621 3145 11655 3179
rect 15485 3145 15519 3179
rect 6561 3077 6595 3111
rect 8493 3077 8527 3111
rect 12909 3077 12943 3111
rect 14657 3077 14691 3111
rect 2053 3009 2087 3043
rect 3249 3009 3283 3043
rect 3433 3009 3467 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 4813 3009 4847 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 6469 3009 6503 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 9413 3009 9447 3043
rect 9965 3009 9999 3043
rect 10149 3009 10183 3043
rect 10609 3009 10643 3043
rect 10793 3009 10827 3043
rect 10885 3009 10919 3043
rect 11989 3009 12023 3043
rect 12173 3009 12207 3043
rect 15301 3009 15335 3043
rect 15485 3009 15519 3043
rect 15853 3009 15887 3043
rect 15945 3009 15979 3043
rect 1961 2941 1995 2975
rect 5089 2941 5123 2975
rect 5457 2941 5491 2975
rect 7297 2941 7331 2975
rect 8033 2941 8067 2975
rect 9137 2941 9171 2975
rect 12633 2941 12667 2975
rect 3433 2873 3467 2907
rect 4905 2873 4939 2907
rect 9321 2873 9355 2907
rect 2421 2805 2455 2839
rect 4077 2805 4111 2839
rect 9229 2805 9263 2839
rect 12081 2805 12115 2839
rect 2881 2601 2915 2635
rect 4537 2601 4571 2635
rect 6837 2601 6871 2635
rect 9137 2601 9171 2635
rect 10425 2601 10459 2635
rect 10609 2601 10643 2635
rect 11253 2601 11287 2635
rect 2145 2533 2179 2567
rect 5825 2533 5859 2567
rect 11805 2533 11839 2567
rect 2513 2465 2547 2499
rect 3433 2465 3467 2499
rect 4353 2465 4387 2499
rect 8309 2465 8343 2499
rect 11437 2465 11471 2499
rect 13829 2465 13863 2499
rect 14197 2465 14231 2499
rect 1869 2397 1903 2431
rect 1961 2397 1995 2431
rect 2605 2397 2639 2431
rect 4261 2397 4295 2431
rect 7941 2397 7975 2431
rect 8033 2397 8067 2431
rect 9045 2397 9079 2431
rect 9689 2397 9723 2431
rect 10149 2397 10183 2431
rect 11161 2397 11195 2431
rect 5457 2329 5491 2363
rect 8401 2329 8435 2363
rect 9597 2329 9631 2363
rect 10793 2329 10827 2363
rect 11437 2329 11471 2363
rect 13553 2329 13587 2363
rect 14473 2329 14507 2363
rect 7205 2261 7239 2295
rect 7757 2261 7791 2295
rect 10057 2261 10091 2295
rect 10593 2261 10627 2295
rect 12081 2261 12115 2295
rect 15945 2261 15979 2295
rect 1685 2057 1719 2091
rect 11713 2057 11747 2091
rect 13737 2057 13771 2091
rect 5825 1989 5859 2023
rect 6745 1989 6779 2023
rect 7573 1989 7607 2023
rect 9321 1989 9355 2023
rect 10701 1989 10735 2023
rect 15209 1989 15243 2023
rect 15761 1989 15795 2023
rect 17601 1989 17635 2023
rect 3709 1921 3743 1955
rect 6929 1921 6963 1955
rect 7021 1921 7055 1955
rect 10057 1921 10091 1955
rect 10241 1921 10275 1955
rect 10517 1921 10551 1955
rect 10793 1921 10827 1955
rect 10885 1921 10919 1955
rect 13461 1921 13495 1955
rect 16865 1921 16899 1955
rect 3157 1853 3191 1887
rect 3433 1853 3467 1887
rect 4353 1853 4387 1887
rect 6101 1853 6135 1887
rect 6745 1853 6779 1887
rect 7297 1853 7331 1887
rect 13185 1853 13219 1887
rect 15485 1853 15519 1887
rect 9689 1785 9723 1819
rect 11069 1785 11103 1819
rect 3801 1717 3835 1751
rect 10149 1717 10183 1751
rect 2329 1513 2363 1547
rect 6009 1513 6043 1547
rect 8137 1513 8171 1547
rect 9137 1513 9171 1547
rect 12265 1513 12299 1547
rect 14644 1513 14678 1547
rect 16129 1513 16163 1547
rect 4353 1445 4387 1479
rect 5365 1445 5399 1479
rect 11713 1445 11747 1479
rect 3249 1377 3283 1411
rect 4169 1377 4203 1411
rect 6653 1377 6687 1411
rect 9689 1377 9723 1411
rect 14381 1377 14415 1411
rect 1777 1309 1811 1343
rect 2421 1309 2455 1343
rect 2697 1309 2731 1343
rect 3157 1309 3191 1343
rect 3341 1309 3375 1343
rect 4445 1309 4479 1343
rect 4721 1309 4755 1343
rect 5273 1309 5307 1343
rect 5917 1309 5951 1343
rect 6101 1309 6135 1343
rect 8401 1309 8435 1343
rect 9413 1309 9447 1343
rect 12173 1309 12207 1343
rect 13829 1241 13863 1275
rect 1869 1173 1903 1207
rect 4169 1173 4203 1207
rect 11161 1173 11195 1207
<< metal1 >>
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 15838 13920 15844 13932
rect 15068 13892 15844 13920
rect 15068 13880 15074 13892
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 15194 13784 15200 13796
rect 7248 13756 15200 13784
rect 7248 13744 7254 13756
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 1118 13676 1124 13728
rect 1176 13716 1182 13728
rect 4798 13716 4804 13728
rect 1176 13688 4804 13716
rect 1176 13676 1182 13688
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 17402 13716 17408 13728
rect 11296 13688 17408 13716
rect 11296 13676 11302 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 1104 13626 18860 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 18860 13626
rect 1104 13552 18860 13574
rect 7190 13472 7196 13524
rect 7248 13472 7254 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10100 13484 10701 13512
rect 10100 13472 10106 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 11149 13515 11207 13521
rect 11149 13481 11161 13515
rect 11195 13512 11207 13515
rect 16393 13515 16451 13521
rect 11195 13484 15240 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13444 3019 13447
rect 7006 13444 7012 13456
rect 3007 13416 7012 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 11238 13404 11244 13456
rect 11296 13404 11302 13456
rect 12084 13416 14964 13444
rect 1026 13336 1032 13388
rect 1084 13376 1090 13388
rect 1486 13376 1492 13388
rect 1084 13348 1492 13376
rect 1084 13336 1090 13348
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 3936 13348 4445 13376
rect 3936 13336 3942 13348
rect 4433 13345 4445 13348
rect 4479 13376 4491 13379
rect 7561 13379 7619 13385
rect 4479 13348 6868 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5074 13308 5080 13320
rect 5031 13280 5080 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 3252 13184 3280 13271
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13209 3939 13243
rect 3881 13203 3939 13209
rect 1854 13132 1860 13184
rect 1912 13132 1918 13184
rect 2498 13132 2504 13184
rect 2556 13132 2562 13184
rect 3234 13132 3240 13184
rect 3292 13132 3298 13184
rect 3421 13175 3479 13181
rect 3421 13141 3433 13175
rect 3467 13172 3479 13175
rect 3896 13172 3924 13203
rect 3970 13200 3976 13252
rect 4028 13200 4034 13252
rect 5445 13243 5503 13249
rect 5445 13209 5457 13243
rect 5491 13209 5503 13243
rect 5445 13203 5503 13209
rect 5537 13243 5595 13249
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 5813 13243 5871 13249
rect 5813 13240 5825 13243
rect 5583 13212 5825 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 5813 13209 5825 13212
rect 5859 13209 5871 13243
rect 6840 13240 6868 13348
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 7607 13348 8493 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 10594 13376 10600 13388
rect 9539 13348 10600 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 7926 13268 7932 13320
rect 7984 13268 7990 13320
rect 9758 13289 9816 13295
rect 9758 13255 9770 13289
rect 9804 13255 9816 13289
rect 9950 13268 9956 13320
rect 10008 13268 10014 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10502 13308 10508 13320
rect 10459 13280 10508 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 11256 13317 11284 13404
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 8389 13243 8447 13249
rect 6840 13212 8248 13240
rect 5813 13203 5871 13209
rect 3467 13144 3924 13172
rect 5460 13172 5488 13203
rect 5626 13172 5632 13184
rect 5460 13144 5632 13172
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 5994 13132 6000 13184
rect 6052 13132 6058 13184
rect 6641 13175 6699 13181
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 6914 13172 6920 13184
rect 6687 13144 6920 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7653 13175 7711 13181
rect 7653 13141 7665 13175
rect 7699 13172 7711 13175
rect 8110 13172 8116 13184
rect 7699 13144 8116 13172
rect 7699 13141 7711 13144
rect 7653 13135 7711 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8220 13172 8248 13212
rect 8389 13209 8401 13243
rect 8435 13240 8447 13243
rect 8754 13240 8760 13252
rect 8435 13212 8760 13240
rect 8435 13209 8447 13212
rect 8389 13203 8447 13209
rect 8754 13200 8760 13212
rect 8812 13240 8818 13252
rect 9758 13249 9816 13255
rect 9309 13243 9367 13249
rect 9309 13240 9321 13243
rect 8812 13212 9321 13240
rect 8812 13200 8818 13212
rect 9309 13209 9321 13212
rect 9355 13209 9367 13243
rect 9309 13203 9367 13209
rect 9398 13172 9404 13184
rect 8220 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9784 13172 9812 13249
rect 9861 13243 9919 13249
rect 9861 13209 9873 13243
rect 9907 13240 9919 13243
rect 10134 13240 10140 13252
rect 9907 13212 10140 13240
rect 9907 13209 9919 13212
rect 9861 13203 9919 13209
rect 10134 13200 10140 13212
rect 10192 13240 10198 13252
rect 11624 13240 11652 13271
rect 12084 13249 12112 13416
rect 12986 13376 12992 13388
rect 12636 13348 12992 13376
rect 12636 13317 12664 13348
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13170 13336 13176 13388
rect 13228 13376 13234 13388
rect 13228 13348 14688 13376
rect 13228 13336 13234 13348
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 12851 13280 13676 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 10192 13212 11652 13240
rect 11808 13212 12081 13240
rect 10192 13200 10198 13212
rect 10410 13172 10416 13184
rect 9784 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11808 13172 11836 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 12069 13203 12127 13209
rect 12161 13243 12219 13249
rect 12161 13209 12173 13243
rect 12207 13240 12219 13243
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 12207 13212 13185 13240
rect 12207 13209 12219 13212
rect 12161 13203 12219 13209
rect 13173 13209 13185 13212
rect 13219 13209 13231 13243
rect 13648 13240 13676 13280
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 14384 13317 14412 13348
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 13648 13212 14412 13240
rect 13173 13203 13231 13209
rect 11296 13144 11836 13172
rect 11296 13132 11302 13144
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12032 13144 12633 13172
rect 12032 13132 12038 13144
rect 12621 13141 12633 13144
rect 12667 13141 12679 13175
rect 12621 13135 12679 13141
rect 13078 13132 13084 13184
rect 13136 13132 13142 13184
rect 13538 13132 13544 13184
rect 13596 13132 13602 13184
rect 14384 13181 14412 13212
rect 14369 13175 14427 13181
rect 14369 13141 14381 13175
rect 14415 13141 14427 13175
rect 14568 13172 14596 13271
rect 14660 13252 14688 13348
rect 14936 13317 14964 13416
rect 15105 13379 15163 13385
rect 15105 13345 15117 13379
rect 15151 13345 15163 13379
rect 15212 13376 15240 13484
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16574 13512 16580 13524
rect 16439 13484 16580 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16574 13472 16580 13484
rect 16632 13512 16638 13524
rect 17310 13512 17316 13524
rect 16632 13484 17316 13512
rect 16632 13472 16638 13484
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 17681 13379 17739 13385
rect 17681 13376 17693 13379
rect 15212 13348 17693 13376
rect 15105 13339 15163 13345
rect 17681 13345 17693 13348
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13277 14979 13311
rect 15120 13308 15148 13339
rect 15562 13308 15568 13320
rect 15120 13280 15568 13308
rect 14921 13271 14979 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 15712 13280 16773 13308
rect 15712 13268 15718 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 17920 13280 18061 13308
rect 17920 13268 17926 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 14642 13200 14648 13252
rect 14700 13200 14706 13252
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 15841 13243 15899 13249
rect 15841 13240 15853 13243
rect 15160 13212 15853 13240
rect 15160 13200 15166 13212
rect 15841 13209 15853 13212
rect 15887 13209 15899 13243
rect 15841 13203 15899 13209
rect 17586 13200 17592 13252
rect 17644 13200 17650 13252
rect 15194 13172 15200 13184
rect 14568 13144 15200 13172
rect 14369 13135 14427 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 15378 13132 15384 13184
rect 15436 13132 15442 13184
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 17957 13175 18015 13181
rect 17957 13172 17969 13175
rect 17000 13144 17969 13172
rect 17000 13132 17006 13144
rect 17957 13141 17969 13144
rect 18003 13141 18015 13175
rect 17957 13135 18015 13141
rect 1104 13082 18860 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 18860 13082
rect 1104 13008 18860 13030
rect 6454 12968 6460 12980
rect 6196 12940 6460 12968
rect 3050 12860 3056 12912
rect 3108 12900 3114 12912
rect 3970 12900 3976 12912
rect 3108 12872 3976 12900
rect 3108 12860 3114 12872
rect 3970 12860 3976 12872
rect 4028 12860 4034 12912
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12900 4215 12903
rect 5626 12900 5632 12912
rect 4203 12872 5632 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 5626 12860 5632 12872
rect 5684 12900 5690 12912
rect 6089 12903 6147 12909
rect 6089 12900 6101 12903
rect 5684 12872 6101 12900
rect 5684 12860 5690 12872
rect 6089 12869 6101 12872
rect 6135 12869 6147 12903
rect 6089 12863 6147 12869
rect 6196 12844 6224 12940
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 7006 12928 7012 12980
rect 7064 12928 7070 12980
rect 8754 12928 8760 12980
rect 8812 12928 8818 12980
rect 10134 12928 10140 12980
rect 10192 12928 10198 12980
rect 10594 12928 10600 12980
rect 10652 12928 10658 12980
rect 13722 12928 13728 12980
rect 13780 12928 13786 12980
rect 13998 12968 14004 12980
rect 13924 12940 14004 12968
rect 7024 12900 7052 12928
rect 6472 12872 7052 12900
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3878 12832 3884 12844
rect 3743 12804 3884 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 2516 12764 2544 12795
rect 2682 12764 2688 12776
rect 2516 12736 2688 12764
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 2792 12764 2820 12795
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6178 12832 6184 12844
rect 6043 12804 6184 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 3234 12764 3240 12776
rect 2792 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12764 3298 12776
rect 3786 12764 3792 12776
rect 3292 12736 3792 12764
rect 3292 12724 3298 12736
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 4540 12764 4568 12795
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6472 12841 6500 12872
rect 7926 12860 7932 12912
rect 7984 12860 7990 12912
rect 8772 12900 8800 12928
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 8772 12872 8953 12900
rect 8941 12869 8953 12872
rect 8987 12869 8999 12903
rect 8941 12863 8999 12869
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6604 12804 6929 12832
rect 6604 12792 6610 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7944 12832 7972 12860
rect 7432 12804 7972 12832
rect 7432 12792 7438 12804
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8628 12804 8861 12832
rect 8628 12792 8634 12804
rect 8849 12801 8861 12804
rect 8895 12832 8907 12835
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8895 12804 9413 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9683 12835 9741 12841
rect 9683 12801 9695 12835
rect 9729 12832 9741 12835
rect 10152 12832 10180 12928
rect 10612 12900 10640 12928
rect 12713 12903 12771 12909
rect 10612 12872 12434 12900
rect 10612 12841 10640 12872
rect 9729 12804 10180 12832
rect 10597 12835 10655 12841
rect 9729 12801 9741 12804
rect 9683 12795 9741 12801
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 5074 12764 5080 12776
rect 4540 12736 5080 12764
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 10318 12764 10324 12776
rect 6380 12736 10324 12764
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 6380 12696 6408 12736
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 11238 12724 11244 12776
rect 11296 12724 11302 12776
rect 12406 12764 12434 12872
rect 12713 12869 12725 12903
rect 12759 12900 12771 12903
rect 12802 12900 12808 12912
rect 12759 12872 12808 12900
rect 12759 12869 12771 12872
rect 12713 12863 12771 12869
rect 12802 12860 12808 12872
rect 12860 12900 12866 12912
rect 13078 12900 13084 12912
rect 12860 12872 13084 12900
rect 12860 12860 12866 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12912 12764 12940 12795
rect 13446 12792 13452 12844
rect 13504 12832 13510 12844
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13504 12804 13645 12832
rect 13504 12792 13510 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13740 12764 13768 12928
rect 13924 12909 13952 12940
rect 13998 12928 14004 12940
rect 14056 12968 14062 12980
rect 15654 12968 15660 12980
rect 14056 12940 15660 12968
rect 14056 12928 14062 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 13817 12903 13875 12909
rect 13817 12869 13829 12903
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 13909 12903 13967 12909
rect 13909 12869 13921 12903
rect 13955 12869 13967 12903
rect 13909 12863 13967 12869
rect 12406 12736 13768 12764
rect 11606 12696 11612 12708
rect 2455 12668 6408 12696
rect 6564 12668 11612 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 1670 12588 1676 12640
rect 1728 12588 1734 12640
rect 2041 12631 2099 12637
rect 2041 12597 2053 12631
rect 2087 12628 2099 12631
rect 3326 12628 3332 12640
rect 2087 12600 3332 12628
rect 2087 12597 2099 12600
rect 2041 12591 2099 12597
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 6564 12637 6592 12668
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12894 12696 12900 12708
rect 11747 12668 12900 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12894 12656 12900 12668
rect 12952 12696 12958 12708
rect 13630 12696 13636 12708
rect 12952 12668 13636 12696
rect 12952 12656 12958 12668
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13832 12696 13860 12863
rect 15102 12860 15108 12912
rect 15160 12900 15166 12912
rect 15197 12903 15255 12909
rect 15197 12900 15209 12903
rect 15160 12872 15209 12900
rect 15160 12860 15166 12872
rect 15197 12869 15209 12872
rect 15243 12869 15255 12903
rect 15948 12900 15976 12928
rect 16209 12903 16267 12909
rect 16209 12900 16221 12903
rect 15948 12872 16221 12900
rect 15197 12863 15255 12869
rect 16209 12869 16221 12872
rect 16255 12869 16267 12903
rect 16209 12863 16267 12869
rect 17402 12860 17408 12912
rect 17460 12860 17466 12912
rect 18233 12903 18291 12909
rect 18233 12900 18245 12903
rect 17696 12872 18245 12900
rect 17696 12844 17724 12872
rect 18233 12869 18245 12872
rect 18279 12869 18291 12903
rect 18233 12863 18291 12869
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14734 12832 14740 12844
rect 14507 12804 14740 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15562 12832 15568 12844
rect 15427 12804 15568 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15562 12792 15568 12804
rect 15620 12832 15626 12844
rect 15838 12832 15844 12844
rect 15620 12804 15844 12832
rect 15620 12792 15626 12804
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 16758 12792 16764 12844
rect 16816 12792 16822 12844
rect 17678 12792 17684 12844
rect 17736 12792 17742 12844
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15344 12736 15669 12764
rect 15344 12724 15350 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 17770 12764 17776 12776
rect 16163 12736 17776 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 17770 12724 17776 12736
rect 17828 12764 17834 12776
rect 18064 12764 18092 12795
rect 17828 12736 18092 12764
rect 17828 12724 17834 12736
rect 16574 12696 16580 12708
rect 13832 12668 16580 12696
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 4065 12631 4123 12637
rect 4065 12628 4077 12631
rect 3936 12600 4077 12628
rect 3936 12588 3942 12600
rect 4065 12597 4077 12600
rect 4111 12597 4123 12631
rect 4065 12591 4123 12597
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7926 12628 7932 12640
rect 7055 12600 7932 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 9456 12600 13369 12628
rect 9456 12588 9462 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 13357 12591 13415 12597
rect 1104 12538 18860 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 18860 12538
rect 1104 12464 18860 12486
rect 5074 12384 5080 12436
rect 5132 12384 5138 12436
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 9217 12427 9275 12433
rect 6604 12396 7236 12424
rect 6604 12384 6610 12396
rect 2590 12316 2596 12368
rect 2648 12356 2654 12368
rect 7208 12356 7236 12396
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9674 12424 9680 12436
rect 9263 12396 9680 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 13173 12427 13231 12433
rect 13173 12424 13185 12427
rect 9784 12396 13185 12424
rect 9784 12356 9812 12396
rect 13173 12393 13185 12396
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 13538 12384 13544 12436
rect 13596 12384 13602 12436
rect 13078 12356 13084 12368
rect 2648 12328 4568 12356
rect 7208 12328 9812 12356
rect 9968 12328 13084 12356
rect 2648 12316 2654 12328
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 3142 12288 3148 12300
rect 1636 12260 3148 12288
rect 1636 12248 1642 12260
rect 1670 12180 1676 12232
rect 1728 12180 1734 12232
rect 1872 12229 1900 12260
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4540 12297 4568 12328
rect 7300 12297 7328 12328
rect 4525 12291 4583 12297
rect 3252 12260 4200 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3050 12220 3056 12232
rect 3007 12192 3056 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 1688 12152 1716 12180
rect 1688 12124 2452 12152
rect 1670 12044 1676 12096
rect 1728 12044 1734 12096
rect 2424 12093 2452 12124
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 3252 12152 3280 12260
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 4062 12220 4068 12232
rect 3384 12192 4068 12220
rect 3384 12180 3390 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4172 12220 4200 12260
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 7285 12291 7343 12297
rect 4755 12260 7144 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 5537 12223 5595 12229
rect 4172 12192 4660 12220
rect 2556 12124 3280 12152
rect 2556 12112 2562 12124
rect 3970 12112 3976 12164
rect 4028 12112 4034 12164
rect 4632 12161 4660 12192
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 6178 12220 6184 12232
rect 5583 12192 6184 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12220 6515 12223
rect 6546 12220 6552 12232
rect 6503 12192 6552 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12222 6791 12223
rect 6914 12222 6920 12232
rect 6779 12194 6920 12222
rect 6779 12189 6791 12194
rect 6733 12183 6791 12189
rect 6914 12180 6920 12194
rect 6972 12180 6978 12232
rect 4157 12155 4215 12161
rect 4157 12121 4169 12155
rect 4203 12121 4215 12155
rect 4157 12115 4215 12121
rect 4617 12155 4675 12161
rect 4617 12121 4629 12155
rect 4663 12121 4675 12155
rect 4617 12115 4675 12121
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12152 5871 12155
rect 5994 12152 6000 12164
rect 5859 12124 6000 12152
rect 5859 12121 5871 12124
rect 5813 12115 5871 12121
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2590 12084 2596 12096
rect 2455 12056 2596 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 3418 12044 3424 12096
rect 3476 12044 3482 12096
rect 4172 12084 4200 12115
rect 5994 12112 6000 12124
rect 6052 12152 6058 12164
rect 6638 12152 6644 12164
rect 6052 12124 6644 12152
rect 6052 12112 6058 12124
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 6822 12112 6828 12164
rect 6880 12112 6886 12164
rect 7116 12152 7144 12260
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 9582 12288 9588 12300
rect 8076 12260 9588 12288
rect 8076 12248 8082 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9968 12297 9996 12328
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 13556 12356 13584 12384
rect 13188 12328 13584 12356
rect 9953 12291 10011 12297
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 7650 12180 7656 12232
rect 7708 12180 7714 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8168 12192 8309 12220
rect 8168 12180 8174 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8496 12192 8708 12220
rect 8496 12152 8524 12192
rect 7116 12124 8524 12152
rect 8570 12112 8576 12164
rect 8628 12112 8634 12164
rect 8588 12084 8616 12112
rect 4172 12056 8616 12084
rect 8680 12084 8708 12192
rect 9122 12180 9128 12232
rect 9180 12229 9186 12232
rect 9180 12220 9189 12229
rect 9309 12223 9367 12229
rect 9180 12192 9260 12220
rect 9180 12183 9189 12192
rect 9180 12180 9186 12183
rect 9232 12152 9260 12192
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9968 12220 9996 12251
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 12032 12260 12173 12288
rect 12032 12248 12038 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13188 12288 13216 12328
rect 17402 12316 17408 12368
rect 17460 12356 17466 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 17460 12328 17693 12356
rect 17460 12316 17466 12328
rect 17681 12325 17693 12328
rect 17727 12325 17739 12359
rect 17681 12319 17739 12325
rect 12759 12260 13216 12288
rect 15197 12291 15255 12297
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 15197 12257 15209 12291
rect 15243 12288 15255 12291
rect 15378 12288 15384 12300
rect 15243 12260 15384 12288
rect 15243 12257 15255 12260
rect 15197 12251 15255 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17770 12288 17776 12300
rect 17359 12260 17776 12288
rect 17359 12257 17371 12260
rect 17313 12251 17371 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 9355 12192 9996 12220
rect 10781 12223 10839 12229
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 10781 12189 10793 12223
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 9858 12152 9864 12164
rect 9232 12124 9864 12152
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10686 12152 10692 12164
rect 10183 12124 10692 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10686 12112 10692 12124
rect 10744 12112 10750 12164
rect 10796 12152 10824 12183
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 10928 12192 11253 12220
rect 10928 12180 10934 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 11388 12192 11437 12220
rect 11388 12180 11394 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 12802 12220 12808 12232
rect 12667 12192 12808 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13449 12223 13507 12229
rect 13070 12201 13128 12207
rect 13070 12167 13082 12201
rect 13116 12167 13128 12201
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 11146 12152 11152 12164
rect 10796 12124 11152 12152
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 11698 12112 11704 12164
rect 11756 12112 11762 12164
rect 11790 12112 11796 12164
rect 11848 12112 11854 12164
rect 13070 12161 13128 12167
rect 13096 12096 13124 12161
rect 9950 12084 9956 12096
rect 8680 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 10318 12084 10324 12096
rect 10091 12056 10324 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10502 12044 10508 12096
rect 10560 12044 10566 12096
rect 10962 12044 10968 12096
rect 11020 12044 11026 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13464 12084 13492 12183
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13688 12192 14197 12220
rect 13688 12180 13694 12192
rect 14185 12189 14197 12192
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 14734 12220 14740 12232
rect 14691 12192 14740 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15102 12180 15108 12232
rect 15160 12180 15166 12232
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15344 12192 15761 12220
rect 15344 12180 15350 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 15896 12192 16681 12220
rect 15896 12180 15902 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 16816 12192 18153 12220
rect 16816 12180 16822 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 17589 12155 17647 12161
rect 17589 12152 17601 12155
rect 14608 12124 17601 12152
rect 14608 12112 14614 12124
rect 17589 12121 17601 12124
rect 17635 12121 17647 12155
rect 17589 12115 17647 12121
rect 13412 12056 13492 12084
rect 13412 12044 13418 12056
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 16574 12084 16580 12096
rect 13688 12056 16580 12084
rect 13688 12044 13694 12056
rect 16574 12044 16580 12056
rect 16632 12084 16638 12096
rect 17126 12084 17132 12096
rect 16632 12056 17132 12084
rect 16632 12044 16638 12056
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 1104 11994 18860 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 18860 11994
rect 1104 11920 18860 11942
rect 1670 11840 1676 11892
rect 1728 11840 1734 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 4028 11852 4261 11880
rect 4028 11840 4034 11852
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6178 11880 6184 11892
rect 6043 11852 6184 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 7064 11852 8861 11880
rect 7064 11840 7070 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9401 11883 9459 11889
rect 8996 11852 9352 11880
rect 8996 11840 9002 11852
rect 1688 11753 1716 11840
rect 2041 11815 2099 11821
rect 2041 11781 2053 11815
rect 2087 11812 2099 11815
rect 8018 11812 8024 11824
rect 2087 11784 2452 11812
rect 2087 11781 2099 11784
rect 2041 11775 2099 11781
rect 2424 11756 2452 11784
rect 7576 11784 8024 11812
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 2148 11540 2176 11707
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 5718 11744 5724 11756
rect 5491 11716 5724 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 4448 11676 4476 11707
rect 5718 11704 5724 11716
rect 5776 11744 5782 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5776 11716 5917 11744
rect 5776 11704 5782 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11742 6791 11747
rect 7006 11744 7012 11756
rect 6840 11742 7012 11744
rect 6779 11716 7012 11742
rect 6779 11714 6868 11716
rect 6779 11713 6791 11714
rect 6733 11707 6791 11713
rect 3712 11648 4476 11676
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 3712 11617 3740 11648
rect 4982 11636 4988 11688
rect 5040 11636 5046 11688
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 6564 11620 6592 11707
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7369 11753 7427 11759
rect 7576 11753 7604 11784
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 8168 11784 8309 11812
rect 8168 11772 8174 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8297 11775 8355 11781
rect 8389 11815 8447 11821
rect 8389 11781 8401 11815
rect 8435 11812 8447 11815
rect 9214 11812 9220 11824
rect 8435 11784 9220 11812
rect 8435 11781 8447 11784
rect 8389 11775 8447 11781
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 9324 11812 9352 11852
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 9858 11880 9864 11892
rect 9447 11852 9864 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 11609 11883 11667 11889
rect 10244 11852 11376 11880
rect 10244 11812 10272 11852
rect 11348 11824 11376 11852
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 11790 11880 11796 11892
rect 11655 11852 11796 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12986 11880 12992 11892
rect 12406 11852 12992 11880
rect 9324 11784 9904 11812
rect 7369 11750 7381 11753
rect 7208 11744 7381 11750
rect 7156 11722 7381 11744
rect 7156 11716 7236 11722
rect 7369 11719 7381 11722
rect 7415 11719 7427 11753
rect 7156 11704 7162 11716
rect 7369 11713 7427 11719
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 6748 11648 7481 11676
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 3016 11580 3709 11608
rect 3016 11568 3022 11580
rect 3697 11577 3709 11580
rect 3743 11577 3755 11611
rect 3697 11571 3755 11577
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 6748 11608 6776 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7576 11676 7604 11707
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8849 11747 8907 11753
rect 8849 11744 8861 11747
rect 7984 11716 8861 11744
rect 7984 11704 7990 11716
rect 8849 11713 8861 11716
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 7576 11648 7696 11676
rect 7469 11639 7527 11645
rect 6604 11580 6776 11608
rect 6604 11568 6610 11580
rect 6822 11540 6828 11552
rect 2148 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7668 11540 7696 11648
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7800 11648 7849 11676
rect 7800 11636 7806 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 9048 11608 9076 11707
rect 9324 11676 9352 11707
rect 9674 11676 9680 11688
rect 9324 11648 9680 11676
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9769 11679 9827 11685
rect 9769 11645 9781 11679
rect 9815 11645 9827 11679
rect 9876 11676 9904 11784
rect 9968 11784 10272 11812
rect 10321 11815 10379 11821
rect 9968 11753 9996 11784
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 10502 11812 10508 11824
rect 10367 11784 10508 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 10612 11784 11161 11812
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10612 11744 10640 11784
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 11330 11772 11336 11824
rect 11388 11772 11394 11824
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 12406 11812 12434 11852
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 13596 11852 14013 11880
rect 13596 11840 13602 11852
rect 14001 11849 14013 11852
rect 14047 11849 14059 11883
rect 15286 11880 15292 11892
rect 14001 11843 14059 11849
rect 14108 11852 15292 11880
rect 14108 11812 14136 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15841 11883 15899 11889
rect 15841 11849 15853 11883
rect 15887 11880 15899 11883
rect 16758 11880 16764 11892
rect 15887 11852 16764 11880
rect 15887 11849 15899 11852
rect 15841 11843 15899 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 15010 11812 15016 11824
rect 11756 11784 12434 11812
rect 12912 11784 14136 11812
rect 14325 11784 15016 11812
rect 11756 11772 11762 11784
rect 10100 11716 10640 11744
rect 10781 11747 10839 11753
rect 10100 11704 10106 11716
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 10870 11744 10876 11756
rect 10827 11716 10876 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11744 11299 11747
rect 11974 11744 11980 11756
rect 11287 11716 11980 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12912 11744 12940 11784
rect 12176 11716 12940 11744
rect 12989 11747 13047 11753
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 9876 11648 12081 11676
rect 9769 11639 9827 11645
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 9784 11608 9812 11639
rect 10229 11611 10287 11617
rect 9048 11580 9674 11608
rect 9784 11580 10180 11608
rect 7147 11512 7696 11540
rect 9646 11540 9674 11580
rect 10042 11540 10048 11552
rect 9646 11512 10048 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10152 11540 10180 11580
rect 10229 11577 10241 11611
rect 10275 11608 10287 11611
rect 12176 11608 12204 11716
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 13078 11744 13084 11756
rect 13035 11716 13084 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13538 11744 13544 11756
rect 13219 11716 13544 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 13998 11744 14004 11756
rect 13688 11716 14004 11744
rect 13688 11704 13694 11716
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14185 11737 14243 11743
rect 14185 11703 14197 11737
rect 14231 11734 14243 11737
rect 14325 11734 14353 11784
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 16574 11772 16580 11824
rect 16632 11772 16638 11824
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 18417 11815 18475 11821
rect 18417 11812 18429 11815
rect 17644 11784 18429 11812
rect 17644 11772 17650 11784
rect 18417 11781 18429 11784
rect 18463 11781 18475 11815
rect 18417 11775 18475 11781
rect 14231 11706 14353 11734
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11713 14519 11747
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14461 11707 14519 11713
rect 14568 11716 15485 11744
rect 14231 11703 14243 11706
rect 14185 11697 14243 11703
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12618 11676 12624 11688
rect 12299 11648 12624 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 10275 11580 12204 11608
rect 12636 11608 12664 11636
rect 14366 11608 14372 11620
rect 12636 11580 14372 11608
rect 10275 11577 10287 11580
rect 10229 11571 10287 11577
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 10502 11540 10508 11552
rect 10152 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10686 11500 10692 11552
rect 10744 11500 10750 11552
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11540 12771 11543
rect 13170 11540 13176 11552
rect 12759 11512 13176 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 13170 11500 13176 11512
rect 13228 11540 13234 11552
rect 13630 11540 13636 11552
rect 13228 11512 13636 11540
rect 13228 11500 13234 11512
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14476 11540 14504 11707
rect 14568 11552 14596 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16592 11744 16620 11772
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16592 11716 16865 11744
rect 16117 11707 16175 11713
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14700 11648 15209 11676
rect 14700 11636 14706 11648
rect 15197 11645 15209 11648
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 15212 11608 15240 11639
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15344 11648 15393 11676
rect 15344 11636 15350 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 15838 11676 15844 11688
rect 15427 11648 15844 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16132 11676 16160 11707
rect 17770 11704 17776 11756
rect 17828 11704 17834 11756
rect 16080 11648 16160 11676
rect 16080 11636 16086 11648
rect 16209 11611 16267 11617
rect 16209 11608 16221 11611
rect 15212 11580 16221 11608
rect 16209 11577 16221 11580
rect 16255 11577 16267 11611
rect 16209 11571 16267 11577
rect 13872 11512 14504 11540
rect 13872 11500 13878 11512
rect 14550 11500 14556 11552
rect 14608 11500 14614 11552
rect 1104 11450 18860 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 18860 11450
rect 1104 11376 18860 11398
rect 1854 11296 1860 11348
rect 1912 11296 1918 11348
rect 2406 11296 2412 11348
rect 2464 11296 2470 11348
rect 2866 11296 2872 11348
rect 2924 11296 2930 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 5534 11336 5540 11348
rect 4019 11308 5540 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6273 11339 6331 11345
rect 5776 11308 5856 11336
rect 5776 11296 5782 11308
rect 1872 11200 1900 11296
rect 1688 11172 1900 11200
rect 2317 11203 2375 11209
rect 1688 11144 1716 11172
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 2424 11200 2452 11296
rect 2884 11209 2912 11296
rect 5828 11277 5856 11308
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6454 11336 6460 11348
rect 6319 11308 6460 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 7650 11336 7656 11348
rect 6687 11308 7656 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 7984 11308 8585 11336
rect 7984 11296 7990 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 10410 11336 10416 11348
rect 9447 11308 10416 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 10689 11339 10747 11345
rect 10689 11305 10701 11339
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 11563 11308 14688 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 5813 11271 5871 11277
rect 5813 11237 5825 11271
rect 5859 11237 5871 11271
rect 6472 11268 6500 11296
rect 6730 11268 6736 11280
rect 6472 11240 6736 11268
rect 5813 11231 5871 11237
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 6822 11228 6828 11280
rect 6880 11268 6886 11280
rect 10704 11268 10732 11299
rect 6880 11240 10732 11268
rect 6880 11228 6886 11240
rect 12618 11228 12624 11280
rect 12676 11228 12682 11280
rect 14185 11271 14243 11277
rect 14185 11268 14197 11271
rect 13464 11240 14197 11268
rect 2363 11172 2452 11200
rect 2869 11203 2927 11209
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 2869 11169 2881 11203
rect 2915 11169 2927 11203
rect 4614 11200 4620 11212
rect 2869 11163 2927 11169
rect 4356 11172 4620 11200
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2590 11132 2596 11144
rect 1903 11104 2596 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2590 11092 2596 11104
rect 2648 11132 2654 11144
rect 3694 11132 3700 11144
rect 2648 11104 3700 11132
rect 2648 11092 2654 11104
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 4356 11141 4384 11172
rect 4614 11160 4620 11172
rect 4672 11200 4678 11212
rect 4982 11200 4988 11212
rect 4672 11172 4988 11200
rect 4672 11160 4678 11172
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 7006 11200 7012 11212
rect 6840 11172 7012 11200
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 5534 11092 5540 11144
rect 5592 11092 5598 11144
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 6840 11132 6868 11172
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 11149 11203 11207 11209
rect 7116 11172 8892 11200
rect 6779 11104 6868 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7116 11141 7144 11172
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6972 11104 7113 11132
rect 6972 11092 6978 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7558 11132 7564 11144
rect 7331 11104 7564 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 8570 11132 8576 11144
rect 8527 11104 8576 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 1765 11067 1823 11073
rect 1765 11033 1777 11067
rect 1811 11064 1823 11067
rect 2777 11067 2835 11073
rect 1811 11036 2728 11064
rect 1811 11033 1823 11036
rect 1765 11027 1823 11033
rect 2700 10996 2728 11036
rect 2777 11033 2789 11067
rect 2823 11064 2835 11067
rect 2866 11064 2872 11076
rect 2823 11036 2872 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 3326 11024 3332 11076
rect 3384 11024 3390 11076
rect 7374 11024 7380 11076
rect 7432 11024 7438 11076
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 8036 11064 8064 11095
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 8711 11104 8800 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 8772 11064 8800 11104
rect 7800 11036 8800 11064
rect 8864 11064 8892 11172
rect 9508 11172 10824 11200
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9398 11132 9404 11144
rect 9355 11104 9404 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9508 11141 9536 11172
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 9582 11092 9588 11144
rect 9640 11092 9646 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 9600 11064 9628 11092
rect 8864 11036 9628 11064
rect 7800 11024 7806 11036
rect 8772 11008 8800 11036
rect 9968 11008 9996 11095
rect 10042 11024 10048 11076
rect 10100 11024 10106 11076
rect 10152 11064 10180 11095
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10796 11141 10824 11172
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 12636 11200 12664 11228
rect 11195 11172 12020 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10376 11104 10609 11132
rect 10376 11092 10382 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 10827 11104 11008 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 10152 11036 10916 11064
rect 10888 11008 10916 11036
rect 10980 11008 11008 11104
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11624 11064 11652 11095
rect 11112 11036 11652 11064
rect 11112 11024 11118 11036
rect 3418 10996 3424 11008
rect 2700 10968 3424 10996
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 3513 10999 3571 11005
rect 3513 10965 3525 10999
rect 3559 10996 3571 10999
rect 3970 10996 3976 11008
rect 3559 10968 3976 10996
rect 3559 10965 3571 10968
rect 3513 10959 3571 10965
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 4065 10999 4123 11005
rect 4065 10965 4077 10999
rect 4111 10996 4123 10999
rect 5350 10996 5356 11008
rect 4111 10968 5356 10996
rect 4111 10965 4123 10968
rect 4065 10959 4123 10965
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 7929 10999 7987 11005
rect 7929 10965 7941 10999
rect 7975 10996 7987 10999
rect 8110 10996 8116 11008
rect 7975 10968 8116 10996
rect 7975 10965 7987 10968
rect 7929 10959 7987 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 9950 10956 9956 11008
rect 10008 10956 10014 11008
rect 10870 10956 10876 11008
rect 10928 10956 10934 11008
rect 10962 10956 10968 11008
rect 11020 10956 11026 11008
rect 11992 10996 12020 11172
rect 12360 11172 12664 11200
rect 12360 11141 12388 11172
rect 13354 11160 13360 11212
rect 13412 11160 13418 11212
rect 13464 11209 13492 11240
rect 14185 11237 14197 11240
rect 14231 11237 14243 11271
rect 14185 11231 14243 11237
rect 14366 11228 14372 11280
rect 14424 11228 14430 11280
rect 14660 11268 14688 11308
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15197 11339 15255 11345
rect 15197 11336 15209 11339
rect 14792 11308 15209 11336
rect 14792 11296 14798 11308
rect 15197 11305 15209 11308
rect 15243 11305 15255 11339
rect 15197 11299 15255 11305
rect 15494 11308 16896 11336
rect 15494 11268 15522 11308
rect 14660 11240 15522 11268
rect 16117 11271 16175 11277
rect 16117 11237 16129 11271
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 13538 11160 13544 11212
rect 13596 11160 13602 11212
rect 14384 11200 14412 11228
rect 16132 11200 16160 11231
rect 14384 11172 16160 11200
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12084 11064 12112 11095
rect 12618 11092 12624 11104
rect 12676 11132 12682 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12676 11104 12817 11132
rect 12676 11092 12682 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 12084 11036 12449 11064
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 13556 11064 13584 11160
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 12437 11027 12495 11033
rect 12544 11036 13584 11064
rect 13740 11064 13768 11095
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14310 11135 14368 11141
rect 14310 11132 14322 11135
rect 14056 11104 14322 11132
rect 14056 11092 14062 11104
rect 14310 11101 14322 11104
rect 14356 11101 14368 11135
rect 14310 11095 14368 11101
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14608 11104 14749 11132
rect 14608 11092 14614 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15580 11141 15608 11172
rect 16758 11160 16764 11212
rect 16816 11200 16822 11212
rect 16868 11200 16896 11308
rect 16942 11228 16948 11280
rect 17000 11228 17006 11280
rect 17954 11268 17960 11280
rect 17052 11240 17960 11268
rect 17052 11209 17080 11240
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 17037 11203 17095 11209
rect 16816 11172 16988 11200
rect 16816 11160 16822 11172
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 14976 11104 15393 11132
rect 14976 11092 14982 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 14182 11064 14188 11076
rect 13740 11036 14188 11064
rect 12544 10996 12572 11036
rect 14182 11024 14188 11036
rect 14240 11064 14246 11076
rect 14936 11064 14964 11092
rect 14240 11036 14964 11064
rect 15672 11064 15700 11095
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16172 11104 16497 11132
rect 16172 11092 16178 11104
rect 16485 11101 16497 11104
rect 16531 11101 16543 11135
rect 16960 11132 16988 11172
rect 17037 11169 17049 11203
rect 17083 11169 17095 11203
rect 17037 11163 17095 11169
rect 17862 11160 17868 11212
rect 17920 11160 17926 11212
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 16960 11104 17325 11132
rect 16485 11095 16543 11101
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 17644 11104 18337 11132
rect 17644 11092 17650 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 17773 11067 17831 11073
rect 15672 11036 17724 11064
rect 14240 11024 14246 11036
rect 11992 10968 12572 10996
rect 14369 10999 14427 11005
rect 14369 10965 14381 10999
rect 14415 10996 14427 10999
rect 14458 10996 14464 11008
rect 14415 10968 14464 10996
rect 14415 10965 14427 10968
rect 14369 10959 14427 10965
rect 14458 10956 14464 10968
rect 14516 10996 14522 11008
rect 15102 10996 15108 11008
rect 14516 10968 15108 10996
rect 14516 10956 14522 10968
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 17696 10996 17724 11036
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 18046 11064 18052 11076
rect 17819 11036 18052 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 18156 11036 18460 11064
rect 18156 10996 18184 11036
rect 18432 11008 18460 11036
rect 17696 10968 18184 10996
rect 18230 10956 18236 11008
rect 18288 10956 18294 11008
rect 18414 10956 18420 11008
rect 18472 10956 18478 11008
rect 1104 10906 18860 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 18860 10906
rect 1104 10832 18860 10854
rect 1486 10752 1492 10804
rect 1544 10752 1550 10804
rect 3160 10764 6684 10792
rect 1504 10665 1532 10752
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 2004 10628 2053 10656
rect 2004 10616 2010 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2314 10616 2320 10668
rect 2372 10616 2378 10668
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10557 2835 10591
rect 2777 10551 2835 10557
rect 2222 10480 2228 10532
rect 2280 10520 2286 10532
rect 2792 10520 2820 10551
rect 2280 10492 2820 10520
rect 2280 10480 2286 10492
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 3160 10452 3188 10764
rect 3326 10684 3332 10736
rect 3384 10684 3390 10736
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 4614 10724 4620 10736
rect 4387 10696 4620 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 5169 10727 5227 10733
rect 5169 10724 5181 10727
rect 4724 10696 5181 10724
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 4724 10665 4752 10696
rect 5169 10693 5181 10696
rect 5215 10724 5227 10727
rect 5534 10724 5540 10736
rect 5215 10696 5540 10724
rect 5215 10693 5227 10696
rect 5169 10687 5227 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 5644 10696 6561 10724
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3476 10628 3985 10656
rect 3476 10616 3482 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4709 10659 4767 10665
rect 4295 10628 4660 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3283 10492 3556 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3528 10464 3556 10492
rect 1627 10424 3188 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 3510 10412 3516 10464
rect 3568 10412 3574 10464
rect 3694 10412 3700 10464
rect 3752 10412 3758 10464
rect 4632 10452 4660 10628
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5644 10656 5672 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6656 10724 6684 10764
rect 7558 10752 7564 10804
rect 7616 10752 7622 10804
rect 8662 10792 8668 10804
rect 7668 10764 8668 10792
rect 7668 10724 7696 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 11422 10792 11428 10804
rect 11195 10764 11428 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 12529 10795 12587 10801
rect 12529 10792 12541 10795
rect 12406 10764 12541 10792
rect 6656 10696 7696 10724
rect 6549 10687 6607 10693
rect 8018 10684 8024 10736
rect 8076 10724 8082 10736
rect 9309 10727 9367 10733
rect 9309 10724 9321 10727
rect 8076 10696 9321 10724
rect 8076 10684 8082 10696
rect 9309 10693 9321 10696
rect 9355 10693 9367 10727
rect 10686 10724 10692 10736
rect 9309 10687 9367 10693
rect 9876 10696 10692 10724
rect 5408 10628 5672 10656
rect 6089 10659 6147 10665
rect 5408 10616 5414 10628
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6135 10628 7052 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 4908 10560 6469 10588
rect 4908 10529 4936 10560
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 6457 10551 6515 10557
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7024 10597 7052 10628
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 8570 10656 8576 10668
rect 7883 10628 8576 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8662 10616 8668 10668
rect 8720 10616 8726 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 7926 10588 7932 10600
rect 7607 10560 7932 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 4893 10523 4951 10529
rect 4893 10489 4905 10523
rect 4939 10489 4951 10523
rect 4893 10483 4951 10489
rect 5902 10480 5908 10532
rect 5960 10520 5966 10532
rect 6822 10520 6828 10532
rect 5960 10492 6828 10520
rect 5960 10480 5966 10492
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 6932 10452 6960 10548
rect 4632 10424 6960 10452
rect 7024 10452 7052 10551
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8864 10588 8892 10619
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 8938 10588 8944 10600
rect 8864 10560 8944 10588
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9416 10588 9444 10619
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9876 10665 9904 10696
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 12253 10727 12311 10733
rect 11020 10696 12020 10724
rect 11020 10684 11026 10696
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9824 10628 9873 10656
rect 9824 10616 9830 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9950 10616 9956 10668
rect 10008 10616 10014 10668
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 11072 10665 11100 10696
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11790 10656 11796 10668
rect 11287 10628 11796 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11992 10656 12020 10696
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12406 10724 12434 10764
rect 12529 10761 12541 10764
rect 12575 10761 12587 10795
rect 12529 10755 12587 10761
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 14274 10792 14280 10804
rect 13035 10764 14280 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 14918 10792 14924 10804
rect 14691 10764 14924 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15010 10752 15016 10804
rect 15068 10752 15074 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15160 10764 16313 10792
rect 15160 10752 15166 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 13078 10724 13084 10736
rect 12299 10696 12434 10724
rect 12820 10696 13084 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 12820 10656 12848 10696
rect 13078 10684 13084 10696
rect 13136 10724 13142 10736
rect 13136 10696 13676 10724
rect 13136 10684 13142 10696
rect 11992 10628 12848 10656
rect 11885 10619 11943 10625
rect 10612 10588 10640 10616
rect 9416 10560 10640 10588
rect 9876 10532 9904 10560
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11480 10560 11713 10588
rect 11480 10548 11486 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11900 10588 11928 10619
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13648 10665 13676 10696
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 13633 10659 13691 10665
rect 12952 10628 13491 10656
rect 12952 10616 12958 10628
rect 11900 10560 12434 10588
rect 11701 10551 11759 10557
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 8113 10523 8171 10529
rect 8113 10520 8125 10523
rect 7156 10492 8125 10520
rect 7156 10480 7162 10492
rect 8113 10489 8125 10492
rect 8159 10489 8171 10523
rect 8113 10483 8171 10489
rect 8849 10523 8907 10529
rect 8849 10489 8861 10523
rect 8895 10520 8907 10523
rect 9582 10520 9588 10532
rect 8895 10492 9588 10520
rect 8895 10489 8907 10492
rect 8849 10483 8907 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 9858 10480 9864 10532
rect 9916 10480 9922 10532
rect 11885 10523 11943 10529
rect 11885 10520 11897 10523
rect 9968 10492 11897 10520
rect 7926 10452 7932 10464
rect 7024 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9968 10452 9996 10492
rect 11885 10489 11897 10492
rect 11931 10489 11943 10523
rect 12406 10520 12434 10560
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 13463 10588 13491 10628
rect 13633 10625 13645 10659
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13832 10588 13860 10684
rect 14384 10665 14412 10752
rect 15212 10696 15608 10724
rect 15212 10668 15240 10696
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 15194 10616 15200 10668
rect 15252 10616 15258 10668
rect 15378 10616 15384 10668
rect 15436 10616 15442 10668
rect 15580 10665 15608 10696
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 18325 10727 18383 10733
rect 18325 10724 18337 10727
rect 18104 10696 18337 10724
rect 18104 10684 18110 10696
rect 18325 10693 18337 10696
rect 18371 10693 18383 10727
rect 18325 10687 18383 10693
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10625 15623 10659
rect 16022 10656 16028 10668
rect 15565 10619 15623 10625
rect 15672 10628 16028 10656
rect 13463 10560 13860 10588
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 14691 10560 15485 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 15672 10520 15700 10628
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 16758 10656 16764 10668
rect 16719 10628 16764 10656
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 18230 10616 18236 10668
rect 18288 10616 18294 10668
rect 12406 10492 14504 10520
rect 11885 10483 11943 10489
rect 14476 10464 14504 10492
rect 15488 10492 15700 10520
rect 15488 10464 15516 10492
rect 9088 10424 9996 10452
rect 9088 10412 9094 10424
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13078 10452 13084 10464
rect 11848 10424 13084 10452
rect 11848 10412 11854 10424
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13228 10424 14013 10452
rect 13228 10412 13234 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 14458 10412 14464 10464
rect 14516 10412 14522 10464
rect 15470 10412 15476 10464
rect 15528 10412 15534 10464
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15712 10424 15945 10452
rect 15712 10412 15718 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 1104 10362 18860 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 18860 10362
rect 1104 10288 18860 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2004 10220 4936 10248
rect 2004 10208 2010 10220
rect 2222 10140 2228 10192
rect 2280 10140 2286 10192
rect 4908 10180 4936 10220
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 7834 10248 7840 10260
rect 5644 10220 7840 10248
rect 5644 10180 5672 10220
rect 7834 10208 7840 10220
rect 7892 10248 7898 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 7892 10220 8125 10248
rect 7892 10208 7898 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8754 10248 8760 10260
rect 8619 10220 8760 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9030 10248 9036 10260
rect 8864 10220 9036 10248
rect 8864 10180 8892 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 9272 10220 9321 10248
rect 9272 10208 9278 10220
rect 9309 10217 9321 10220
rect 9355 10217 9367 10251
rect 9309 10211 9367 10217
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 13265 10251 13323 10257
rect 10008 10220 13216 10248
rect 10008 10208 10014 10220
rect 4908 10152 5672 10180
rect 6656 10152 8892 10180
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1360 10084 1593 10112
rect 1360 10072 1366 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2240 10044 2268 10140
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 3568 10084 5488 10112
rect 3568 10072 3574 10084
rect 1995 10016 2268 10044
rect 3421 10047 3479 10053
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3436 9976 3464 10007
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 5460 10053 5488 10084
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 3436 9948 3893 9976
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 3881 9939 3939 9945
rect 3896 9908 3924 9939
rect 4062 9908 4068 9920
rect 3896 9880 4068 9908
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 4816 9908 4844 10007
rect 6178 9936 6184 9988
rect 6236 9936 6242 9988
rect 6270 9936 6276 9988
rect 6328 9936 6334 9988
rect 6656 9908 6684 10152
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 11333 10183 11391 10189
rect 11333 10180 11345 10183
rect 8996 10152 11345 10180
rect 8996 10140 9002 10152
rect 11333 10149 11345 10152
rect 11379 10149 11391 10183
rect 11790 10180 11796 10192
rect 11333 10143 11391 10149
rect 11716 10152 11796 10180
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 10226 10112 10232 10124
rect 7515 10084 8340 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 6748 10044 6776 10075
rect 7006 10044 7012 10056
rect 6748 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8110 10044 8116 10056
rect 8067 10016 8116 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 7098 9976 7104 9988
rect 6788 9948 7104 9976
rect 6788 9936 6794 9948
rect 7098 9936 7104 9948
rect 7156 9976 7162 9988
rect 7392 9976 7420 10007
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8312 10044 8340 10084
rect 9416 10084 10232 10112
rect 8662 10044 8668 10056
rect 8312 10016 8668 10044
rect 8205 10007 8263 10013
rect 7156 9948 7420 9976
rect 8220 9976 8248 10007
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9306 10044 9312 10056
rect 9263 10016 9312 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9416 10053 9444 10084
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 11716 10121 11744 10152
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12618 10180 12624 10192
rect 11940 10152 12624 10180
rect 11940 10140 11946 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13188 10180 13216 10220
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13446 10248 13452 10260
rect 13311 10220 13452 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13446 10208 13452 10220
rect 13504 10248 13510 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13504 10220 14381 10248
rect 13504 10208 13510 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 18414 10208 18420 10260
rect 18472 10208 18478 10260
rect 13998 10180 14004 10192
rect 13188 10152 14004 10180
rect 13998 10140 14004 10152
rect 14056 10180 14062 10192
rect 14056 10152 14412 10180
rect 14056 10140 14062 10152
rect 11701 10115 11759 10121
rect 10560 10084 11284 10112
rect 10560 10072 10566 10084
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9582 10004 9588 10056
rect 9640 10044 9646 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9640 10016 9689 10044
rect 9640 10004 9646 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9766 10004 9772 10056
rect 9824 10004 9830 10056
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10962 10053 10968 10056
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10468 10016 10793 10044
rect 10468 10004 10474 10016
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10958 10044 10968 10053
rect 10923 10016 10968 10044
rect 10781 10007 10839 10013
rect 10958 10007 10968 10016
rect 10962 10004 10968 10007
rect 11020 10004 11026 10056
rect 11256 10053 11284 10084
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 14182 10072 14188 10124
rect 14240 10072 14246 10124
rect 14384 10112 14412 10152
rect 15749 10115 15807 10121
rect 14384 10084 14504 10112
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11848 10016 11897 10044
rect 11848 10004 11854 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12115 10016 12449 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12802 10044 12808 10056
rect 12667 10016 12808 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13219 10016 13584 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 9784 9976 9812 10004
rect 8220 9948 9812 9976
rect 9953 9979 10011 9985
rect 7156 9936 7162 9948
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10134 9976 10140 9988
rect 9999 9948 10140 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10134 9936 10140 9948
rect 10192 9976 10198 9988
rect 10873 9979 10931 9985
rect 10873 9976 10885 9979
rect 10192 9948 10885 9976
rect 10192 9936 10198 9948
rect 10873 9945 10885 9948
rect 10919 9945 10931 9979
rect 13354 9976 13360 9988
rect 10873 9939 10931 9945
rect 10980 9948 13360 9976
rect 4764 9880 6684 9908
rect 4764 9868 4770 9880
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 10980 9908 11008 9948
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 13556 9976 13584 10016
rect 13630 10004 13636 10056
rect 13688 10004 13694 10056
rect 14476 10053 14504 10084
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 18322 10112 18328 10124
rect 15795 10084 16160 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 16132 10056 16160 10084
rect 17144 10084 18328 10112
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 15304 9976 15332 10007
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 15528 10016 15669 10044
rect 15528 10004 15534 10016
rect 15657 10013 15669 10016
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 15378 9976 15384 9988
rect 13556 9948 14504 9976
rect 15304 9948 15384 9976
rect 14476 9920 14504 9948
rect 15378 9936 15384 9948
rect 15436 9976 15442 9988
rect 16040 9976 16068 10007
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 16172 10016 16313 10044
rect 16172 10004 16178 10016
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17144 9976 17172 10084
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10044 18015 10047
rect 18046 10044 18052 10056
rect 18003 10016 18052 10044
rect 18003 10013 18015 10016
rect 17957 10007 18015 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 15436 9948 15792 9976
rect 16040 9948 17172 9976
rect 17221 9979 17279 9985
rect 15436 9936 15442 9948
rect 15764 9920 15792 9948
rect 17221 9945 17233 9979
rect 17267 9976 17279 9979
rect 18230 9976 18236 9988
rect 17267 9948 18236 9976
rect 17267 9945 17279 9948
rect 17221 9939 17279 9945
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 7984 9880 11008 9908
rect 7984 9868 7990 9880
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12032 9880 12541 9908
rect 12032 9868 12038 9880
rect 12529 9877 12541 9880
rect 12575 9908 12587 9911
rect 12618 9908 12624 9920
rect 12575 9880 12624 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13228 9880 13737 9908
rect 13228 9868 13234 9880
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 13964 9880 14197 9908
rect 13964 9868 13970 9880
rect 14185 9877 14197 9880
rect 14231 9877 14243 9911
rect 14185 9871 14243 9877
rect 14458 9868 14464 9920
rect 14516 9868 14522 9920
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9908 15071 9911
rect 15562 9908 15568 9920
rect 15059 9880 15568 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 15746 9868 15752 9920
rect 15804 9868 15810 9920
rect 17862 9868 17868 9920
rect 17920 9868 17926 9920
rect 1104 9818 18860 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 18860 9818
rect 1104 9744 18860 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 1360 9676 1808 9704
rect 1360 9664 1366 9676
rect 1210 9596 1216 9648
rect 1268 9636 1274 9648
rect 1670 9636 1676 9648
rect 1268 9608 1676 9636
rect 1268 9596 1274 9608
rect 1670 9596 1676 9608
rect 1728 9596 1734 9648
rect 1780 9568 1808 9676
rect 2314 9664 2320 9716
rect 2372 9704 2378 9716
rect 2593 9707 2651 9713
rect 2593 9704 2605 9707
rect 2372 9676 2605 9704
rect 2372 9664 2378 9676
rect 2593 9673 2605 9676
rect 2639 9673 2651 9707
rect 2593 9667 2651 9673
rect 4617 9707 4675 9713
rect 4617 9673 4629 9707
rect 4663 9674 4675 9707
rect 4663 9673 4752 9674
rect 4617 9667 4752 9673
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 3878 9636 3884 9648
rect 1903 9608 3884 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 3970 9596 3976 9648
rect 4028 9596 4034 9648
rect 4632 9646 4752 9667
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 6089 9707 6147 9713
rect 4856 9676 6040 9704
rect 4856 9664 4862 9676
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 1780 9540 2513 9568
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2501 9531 2559 9537
rect 2608 9540 2697 9568
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 2406 9500 2412 9512
rect 1627 9472 2412 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 2608 9500 2636 9540
rect 2685 9537 2697 9540
rect 2731 9568 2743 9571
rect 3050 9568 3056 9580
rect 2731 9540 3056 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3252 9500 3280 9531
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 2464 9472 2636 9500
rect 2700 9472 3280 9500
rect 3789 9503 3847 9509
rect 2464 9460 2470 9472
rect 2700 9376 2728 9472
rect 3789 9469 3801 9503
rect 3835 9469 3847 9503
rect 3988 9500 4016 9596
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 4724 9568 4752 9646
rect 6012 9636 6040 9676
rect 6089 9673 6101 9707
rect 6135 9704 6147 9707
rect 6270 9704 6276 9716
rect 6135 9676 6276 9704
rect 6135 9673 6147 9676
rect 6089 9667 6147 9673
rect 6270 9664 6276 9676
rect 6328 9704 6334 9716
rect 9122 9704 9128 9716
rect 6328 9676 6684 9704
rect 6328 9664 6334 9676
rect 6656 9645 6684 9676
rect 6748 9676 9128 9704
rect 6641 9639 6699 9645
rect 6012 9608 6592 9636
rect 4672 9540 4752 9568
rect 4672 9528 4678 9540
rect 4798 9528 4804 9580
rect 4856 9528 4862 9580
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 6454 9528 6460 9580
rect 6512 9528 6518 9580
rect 6564 9568 6592 9608
rect 6641 9605 6653 9639
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 6748 9568 6776 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 9582 9704 9588 9716
rect 9364 9676 9588 9704
rect 9364 9664 9370 9676
rect 9582 9664 9588 9676
rect 9640 9704 9646 9716
rect 15654 9704 15660 9716
rect 9640 9676 15660 9704
rect 9640 9664 9646 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 7006 9596 7012 9648
rect 7064 9636 7070 9648
rect 8018 9636 8024 9648
rect 7064 9608 8024 9636
rect 7064 9596 7070 9608
rect 7392 9577 7420 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8996 9608 9505 9636
rect 8996 9596 9002 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 9953 9639 10011 9645
rect 9953 9636 9965 9639
rect 9732 9608 9965 9636
rect 9732 9596 9738 9608
rect 9953 9605 9965 9608
rect 9999 9636 10011 9639
rect 10318 9636 10324 9648
rect 9999 9608 10324 9636
rect 9999 9605 10011 9608
rect 9953 9599 10011 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 10755 9639 10813 9645
rect 10755 9605 10767 9639
rect 10801 9636 10813 9639
rect 11514 9636 11520 9648
rect 10801 9608 11520 9636
rect 10801 9605 10813 9608
rect 10755 9599 10813 9605
rect 11514 9596 11520 9608
rect 11572 9636 11578 9648
rect 11609 9639 11667 9645
rect 11609 9636 11621 9639
rect 11572 9608 11621 9636
rect 11572 9596 11578 9608
rect 11609 9605 11621 9608
rect 11655 9605 11667 9639
rect 11609 9599 11667 9605
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 12768 9608 13185 9636
rect 12768 9596 12774 9608
rect 13173 9605 13185 9608
rect 13219 9605 13231 9639
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 13173 9599 13231 9605
rect 13280 9608 16129 9636
rect 6564 9540 6776 9568
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7926 9568 7932 9580
rect 7791 9540 7932 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 8662 9568 8668 9580
rect 8251 9540 8668 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9692 9568 9720 9596
rect 13280 9580 13308 9608
rect 8895 9540 9720 9568
rect 9861 9571 9919 9577
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 10045 9574 10103 9577
rect 10045 9571 10180 9574
rect 10045 9537 10057 9571
rect 10091 9568 10180 9571
rect 10658 9571 10716 9577
rect 10091 9546 10624 9568
rect 10091 9537 10103 9546
rect 10152 9540 10624 9546
rect 10045 9531 10103 9537
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3988 9472 4261 9500
rect 3789 9463 3847 9469
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 9030 9500 9036 9512
rect 4387 9472 5120 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 3804 9432 3832 9463
rect 4706 9432 4712 9444
rect 3804 9404 4712 9432
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 5092 9441 5120 9472
rect 6564 9472 9036 9500
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 5629 9435 5687 9441
rect 5629 9401 5641 9435
rect 5675 9432 5687 9435
rect 6564 9432 6592 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9766 9500 9772 9512
rect 9180 9472 9772 9500
rect 9180 9460 9186 9472
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9876 9500 9904 9531
rect 10410 9500 10416 9512
rect 9876 9472 10416 9500
rect 10060 9444 10088 9472
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 10596 9500 10624 9540
rect 10658 9537 10670 9571
rect 10704 9568 10716 9571
rect 11330 9568 11336 9580
rect 10704 9540 11336 9568
rect 10704 9537 10716 9540
rect 10658 9531 10716 9537
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 12032 9540 12357 9568
rect 12032 9528 12038 9540
rect 12345 9537 12357 9540
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 13556 9577 13584 9608
rect 13448 9571 13506 9577
rect 13448 9537 13460 9571
rect 13494 9537 13506 9571
rect 13448 9531 13506 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 10870 9500 10876 9512
rect 10596 9472 10876 9500
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 11112 9472 11161 9500
rect 11112 9460 11118 9472
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 11664 9472 12449 9500
rect 11664 9460 11670 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9469 12587 9503
rect 13464 9500 13492 9531
rect 13998 9528 14004 9580
rect 14056 9528 14062 9580
rect 14553 9571 14611 9577
rect 14553 9537 14565 9571
rect 14599 9568 14611 9571
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14599 9540 15025 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 14274 9500 14280 9512
rect 13464 9472 14280 9500
rect 12529 9463 12587 9469
rect 5675 9404 6592 9432
rect 5675 9401 5687 9404
rect 5629 9395 5687 9401
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 2682 9324 2688 9376
rect 2740 9324 2746 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3694 9364 3700 9376
rect 3108 9336 3700 9364
rect 3108 9324 3114 9336
rect 3694 9324 3700 9336
rect 3752 9364 3758 9376
rect 5644 9364 5672 9395
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 7800 9404 7972 9432
rect 7800 9392 7806 9404
rect 3752 9336 5672 9364
rect 3752 9324 3758 9336
rect 5994 9324 6000 9376
rect 6052 9324 6058 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7340 9336 7849 9364
rect 7340 9324 7346 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7944 9364 7972 9404
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 8904 9404 9674 9432
rect 8904 9392 8910 9404
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 7944 9336 8493 9364
rect 7837 9327 7895 9333
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 9646 9364 9674 9404
rect 10042 9392 10048 9444
rect 10100 9392 10106 9444
rect 10505 9435 10563 9441
rect 10505 9401 10517 9435
rect 10551 9432 10563 9435
rect 10594 9432 10600 9444
rect 10551 9404 10600 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 11882 9392 11888 9444
rect 11940 9432 11946 9444
rect 12544 9432 12572 9463
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 13262 9432 13268 9444
rect 11940 9404 13268 9432
rect 11940 9392 11946 9404
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14568 9432 14596 9531
rect 15028 9500 15056 9531
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 15470 9528 15476 9580
rect 15528 9577 15534 9580
rect 15672 9577 15700 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 15528 9568 15537 9577
rect 15657 9571 15715 9577
rect 15528 9540 15573 9568
rect 15528 9531 15537 9540
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 15528 9528 15534 9531
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15804 9540 16037 9568
rect 15804 9528 15810 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9537 16267 9571
rect 16942 9568 16948 9580
rect 16209 9531 16267 9537
rect 16500 9540 16948 9568
rect 15378 9500 15384 9512
rect 15028 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 16224 9432 16252 9531
rect 13780 9404 14596 9432
rect 14647 9404 16252 9432
rect 13780 9392 13786 9404
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 9646 9336 11069 9364
rect 8481 9327 8539 9333
rect 11057 9333 11069 9336
rect 11103 9364 11115 9367
rect 11422 9364 11428 9376
rect 11103 9336 11428 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11756 9336 11989 9364
rect 11756 9324 11762 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 11977 9327 12035 9333
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 12618 9364 12624 9376
rect 12124 9336 12624 9364
rect 12124 9324 12130 9336
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14090 9364 14096 9376
rect 13872 9336 14096 9364
rect 13872 9324 13878 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14647 9364 14675 9404
rect 14424 9336 14675 9364
rect 14424 9324 14430 9336
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 15068 9336 15117 9364
rect 15068 9324 15074 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 16500 9364 16528 9540
rect 16942 9528 16948 9540
rect 17000 9568 17006 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 17000 9540 17601 9568
rect 17000 9528 17006 9540
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16632 9472 16773 9500
rect 16632 9460 16638 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 17218 9392 17224 9444
rect 17276 9392 17282 9444
rect 15611 9336 16528 9364
rect 17328 9364 17356 9463
rect 18138 9460 18144 9512
rect 18196 9460 18202 9512
rect 18046 9392 18052 9444
rect 18104 9392 18110 9444
rect 17328 9336 18920 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 1104 9274 18860 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 18860 9274
rect 1104 9200 18860 9222
rect 2130 9120 2136 9172
rect 2188 9120 2194 9172
rect 3878 9120 3884 9172
rect 3936 9120 3942 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6236 9132 7021 9160
rect 6236 9120 6242 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 7009 9123 7067 9129
rect 7926 9120 7932 9172
rect 7984 9120 7990 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8720 9132 9045 9160
rect 8720 9120 8726 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9122 9120 9128 9172
rect 9180 9120 9186 9172
rect 11330 9160 11336 9172
rect 9646 9132 11336 9160
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2148 8956 2176 9120
rect 3896 9092 3924 9120
rect 8573 9095 8631 9101
rect 3896 9064 8524 9092
rect 7282 9024 7288 9036
rect 6748 8996 7288 9024
rect 1811 8928 2176 8956
rect 3237 8959 3295 8965
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3283 8928 3924 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3896 8897 3924 8928
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 6748 8965 6776 8996
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 8496 9024 8524 9064
rect 8573 9061 8585 9095
rect 8619 9092 8631 9095
rect 9140 9092 9168 9120
rect 8619 9064 9168 9092
rect 8619 9061 8631 9064
rect 8573 9055 8631 9061
rect 9214 9052 9220 9104
rect 9272 9092 9278 9104
rect 9646 9092 9674 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12710 9160 12716 9172
rect 12084 9132 12716 9160
rect 9272 9064 9674 9092
rect 9272 9052 9278 9064
rect 10594 9052 10600 9104
rect 10652 9052 10658 9104
rect 12084 9092 12112 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 12805 9163 12863 9169
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 12894 9160 12900 9172
rect 12851 9132 12900 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13814 9160 13820 9172
rect 13372 9132 13820 9160
rect 13372 9092 13400 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14274 9120 14280 9172
rect 14332 9120 14338 9172
rect 15194 9120 15200 9172
rect 15252 9120 15258 9172
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 18046 9120 18052 9172
rect 18104 9120 18110 9172
rect 18325 9163 18383 9169
rect 18325 9129 18337 9163
rect 18371 9160 18383 9163
rect 18892 9160 18920 9336
rect 18371 9132 18920 9160
rect 18371 9129 18383 9132
rect 18325 9123 18383 9129
rect 15212 9092 15240 9120
rect 15933 9095 15991 9101
rect 15933 9092 15945 9095
rect 10704 9064 12112 9092
rect 12268 9064 13400 9092
rect 13464 9064 15148 9092
rect 15212 9064 15945 9092
rect 9398 9024 9404 9036
rect 7484 8996 8156 9024
rect 8496 8996 9404 9024
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4028 8928 4813 8956
rect 4028 8916 4034 8928
rect 4801 8925 4813 8928
rect 4847 8956 4859 8959
rect 5813 8959 5871 8965
rect 4847 8928 5764 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 3329 8891 3387 8897
rect 3329 8888 3341 8891
rect 2746 8860 3341 8888
rect 2746 8832 2774 8860
rect 3329 8857 3341 8860
rect 3375 8857 3387 8891
rect 3329 8851 3387 8857
rect 3881 8891 3939 8897
rect 3881 8857 3893 8891
rect 3927 8857 3939 8891
rect 3881 8851 3939 8857
rect 2682 8780 2688 8832
rect 2740 8792 2774 8832
rect 3896 8820 3924 8851
rect 4062 8848 4068 8900
rect 4120 8848 4126 8900
rect 5169 8891 5227 8897
rect 5169 8857 5181 8891
rect 5215 8888 5227 8891
rect 5215 8860 5488 8888
rect 5215 8857 5227 8860
rect 5169 8851 5227 8857
rect 5460 8832 5488 8860
rect 4798 8820 4804 8832
rect 3896 8792 4804 8820
rect 2740 8780 2746 8792
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 5736 8820 5764 8928
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7239 8928 7420 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 5828 8888 5856 8919
rect 7392 8900 7420 8928
rect 6454 8888 6460 8900
rect 5828 8860 6460 8888
rect 6454 8848 6460 8860
rect 6512 8888 6518 8900
rect 7374 8888 7380 8900
rect 6512 8860 7380 8888
rect 6512 8848 6518 8860
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 7484 8820 7512 8996
rect 7834 8916 7840 8968
rect 7892 8916 7898 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 5736 8792 7512 8820
rect 8036 8820 8064 8919
rect 8128 8888 8156 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8956 8539 8959
rect 8662 8956 8668 8968
rect 8527 8928 8668 8956
rect 8527 8925 8539 8928
rect 8481 8919 8539 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 10612 8956 10640 9052
rect 10704 8965 10732 9064
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 10551 8928 10640 8956
rect 10689 8959 10747 8965
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10689 8919 10747 8925
rect 10796 8928 11345 8956
rect 10597 8891 10655 8897
rect 10597 8888 10609 8891
rect 8128 8860 10609 8888
rect 10597 8857 10609 8860
rect 10643 8857 10655 8891
rect 10597 8851 10655 8857
rect 10796 8832 10824 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 8846 8820 8852 8832
rect 8036 8792 8852 8820
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9398 8780 9404 8832
rect 9456 8780 9462 8832
rect 9490 8780 9496 8832
rect 9548 8780 9554 8832
rect 10778 8780 10784 8832
rect 10836 8780 10842 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 11348 8820 11376 8919
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 12268 8965 12296 9064
rect 13464 9024 13492 9064
rect 13906 9024 13912 9036
rect 12820 8996 13492 9024
rect 13556 8996 13912 9024
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11480 8928 12265 8956
rect 11480 8916 11486 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11885 8891 11943 8897
rect 11885 8888 11897 8891
rect 11756 8860 11897 8888
rect 11756 8848 11762 8860
rect 11885 8857 11897 8860
rect 11931 8857 11943 8891
rect 11885 8851 11943 8857
rect 11977 8891 12035 8897
rect 11977 8857 11989 8891
rect 12023 8888 12035 8891
rect 12618 8888 12624 8900
rect 12023 8860 12624 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 12820 8820 12848 8996
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13446 8956 13452 8968
rect 12943 8928 13452 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 13556 8965 13584 8996
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 15120 9024 15148 9064
rect 15933 9061 15945 9064
rect 15979 9061 15991 9095
rect 15933 9055 15991 9061
rect 17681 9095 17739 9101
rect 17681 9061 17693 9095
rect 17727 9061 17739 9095
rect 17681 9055 17739 9061
rect 17218 9024 17224 9036
rect 15120 8996 17224 9024
rect 17218 8984 17224 8996
rect 17276 9024 17282 9036
rect 17696 9024 17724 9055
rect 17276 8996 17724 9024
rect 17276 8984 17282 8996
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13722 8916 13728 8968
rect 13780 8916 13786 8968
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 13872 8928 14197 8956
rect 13872 8916 13878 8928
rect 14185 8925 14197 8928
rect 14231 8925 14243 8959
rect 14185 8919 14243 8925
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8956 14887 8959
rect 15286 8956 15292 8968
rect 14875 8928 15292 8956
rect 14875 8925 14887 8928
rect 14829 8919 14887 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15470 8956 15476 8968
rect 15427 8928 15476 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 15654 8956 15660 8968
rect 15611 8928 15660 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15764 8928 15853 8956
rect 14734 8888 14740 8900
rect 13372 8860 14740 8888
rect 13372 8832 13400 8860
rect 14734 8848 14740 8860
rect 14792 8888 14798 8900
rect 15764 8888 15792 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15988 8928 16405 8956
rect 15988 8916 15994 8928
rect 16393 8925 16405 8928
rect 16439 8956 16451 8959
rect 16574 8956 16580 8968
rect 16439 8928 16580 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 18064 8956 18092 9120
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18064 8928 18245 8956
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 14792 8860 15792 8888
rect 14792 8848 14798 8860
rect 11348 8792 12848 8820
rect 13354 8780 13360 8832
rect 13412 8780 13418 8832
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 1104 8730 18860 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 18860 8730
rect 1104 8656 18860 8678
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 4614 8576 4620 8628
rect 4672 8576 4678 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 7282 8616 7288 8628
rect 7024 8588 7288 8616
rect 1118 8508 1124 8560
rect 1176 8508 1182 8560
rect 1136 8480 1164 8508
rect 1578 8480 1584 8492
rect 1136 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8480 1642 8492
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1636 8452 1777 8480
rect 1636 8440 1642 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 2148 8480 2176 8576
rect 2682 8508 2688 8560
rect 2740 8508 2746 8560
rect 3237 8551 3295 8557
rect 3237 8517 3249 8551
rect 3283 8548 3295 8551
rect 4080 8548 4108 8576
rect 3283 8520 4108 8548
rect 3283 8517 3295 8520
rect 3237 8511 3295 8517
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 2148 8452 2237 8480
rect 1765 8443 1823 8449
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 2823 8452 3065 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3970 8480 3976 8492
rect 3651 8452 3976 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4080 8489 4108 8520
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 4632 8548 4660 8576
rect 4203 8520 4660 8548
rect 6012 8548 6040 8576
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6012 8520 6469 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 6457 8517 6469 8520
rect 6503 8517 6515 8551
rect 6457 8511 6515 8517
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 4632 8412 4660 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 7024 8489 7052 8588
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7374 8576 7380 8628
rect 7432 8576 7438 8628
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 11388 8588 11713 8616
rect 11388 8576 11394 8588
rect 11701 8585 11713 8588
rect 11747 8616 11759 8619
rect 13170 8616 13176 8628
rect 11747 8588 13176 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13722 8576 13728 8628
rect 13780 8576 13786 8628
rect 13832 8588 15884 8616
rect 9508 8548 9536 8576
rect 7116 8520 9536 8548
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 5442 8412 5448 8424
rect 1872 8384 2774 8412
rect 4632 8384 5448 8412
rect 1872 8353 1900 8384
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8313 1915 8347
rect 2746 8344 2774 8384
rect 5442 8372 5448 8384
rect 5500 8412 5506 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 5500 8384 6561 8412
rect 5500 8372 5506 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 4433 8347 4491 8353
rect 2746 8316 4384 8344
rect 1857 8307 1915 8313
rect 4356 8276 4384 8316
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 4798 8344 4804 8356
rect 4479 8316 4804 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 7116 8344 7144 8520
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 11057 8551 11115 8557
rect 11057 8548 11069 8551
rect 9640 8520 11069 8548
rect 9640 8508 9646 8520
rect 11057 8517 11069 8520
rect 11103 8517 11115 8551
rect 11057 8511 11115 8517
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7484 8356 7512 8443
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7800 8452 8493 8480
rect 7800 8440 7806 8452
rect 8481 8449 8493 8452
rect 8527 8480 8539 8483
rect 8570 8480 8576 8492
rect 8527 8452 8576 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 11164 8489 11192 8576
rect 12084 8520 13768 8548
rect 12084 8492 12112 8520
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9180 8452 9413 8480
rect 9180 8440 9186 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 11149 8483 11207 8489
rect 10367 8452 10640 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 7834 8372 7840 8424
rect 7892 8372 7898 8424
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 10612 8421 10640 8452
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11940 8452 11989 8480
rect 11940 8440 11946 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 13004 8489 13032 8520
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12989 8483 13047 8489
rect 12299 8452 12572 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 4908 8316 7144 8344
rect 4908 8276 4936 8316
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 8938 8344 8944 8356
rect 7524 8316 8944 8344
rect 7524 8304 7530 8316
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 4356 8248 4936 8276
rect 5718 8236 5724 8288
rect 5776 8236 5782 8288
rect 10612 8276 10640 8375
rect 11974 8304 11980 8356
rect 12032 8344 12038 8356
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 12032 8316 12265 8344
rect 12032 8304 12038 8316
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 12544 8344 12572 8452
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13320 8452 13645 8480
rect 13320 8440 13326 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12676 8384 12817 8412
rect 12676 8372 12682 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 13740 8412 13768 8520
rect 13832 8489 13860 8588
rect 15856 8560 15884 8588
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18138 8576 18144 8628
rect 18196 8576 18202 8628
rect 13924 8520 14596 8548
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 13924 8412 13952 8520
rect 14568 8489 14596 8520
rect 15838 8508 15844 8560
rect 15896 8508 15902 8560
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 14553 8483 14611 8489
rect 14231 8452 14504 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 13740 8384 13952 8412
rect 12805 8375 12863 8381
rect 13446 8344 13452 8356
rect 12544 8316 13452 8344
rect 12253 8307 12311 8313
rect 13446 8304 13452 8316
rect 13504 8344 13510 8356
rect 14200 8344 14228 8443
rect 14366 8372 14372 8424
rect 14424 8372 14430 8424
rect 14476 8412 14504 8452
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14700 8452 15025 8480
rect 14700 8440 14706 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15930 8480 15936 8492
rect 15344 8452 15936 8480
rect 15344 8440 15350 8452
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16022 8440 16028 8492
rect 16080 8480 16086 8492
rect 16960 8489 16988 8576
rect 17681 8551 17739 8557
rect 17681 8517 17693 8551
rect 17727 8548 17739 8551
rect 18064 8548 18092 8576
rect 17727 8520 18092 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 16080 8452 16129 8480
rect 16080 8440 16086 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 17920 8452 18337 8480
rect 17920 8440 17926 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 15304 8412 15332 8440
rect 14476 8384 15332 8412
rect 13504 8316 14228 8344
rect 13504 8304 13510 8316
rect 14458 8304 14464 8356
rect 14516 8304 14522 8356
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 15838 8344 15844 8356
rect 15611 8316 15844 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 13538 8276 13544 8288
rect 10612 8248 13544 8276
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 15102 8236 15108 8288
rect 15160 8236 15166 8288
rect 16114 8236 16120 8288
rect 16172 8236 16178 8288
rect 1104 8186 18860 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 18860 8186
rect 1104 8112 18860 8134
rect 1578 8032 1584 8084
rect 1636 8032 1642 8084
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1728 8044 1961 8072
rect 1728 8032 1734 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2406 8032 2412 8084
rect 2464 8032 2470 8084
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6914 8072 6920 8084
rect 6411 8044 6920 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6914 8032 6920 8044
rect 6972 8072 6978 8084
rect 7466 8072 7472 8084
rect 6972 8044 7472 8072
rect 6972 8032 6978 8044
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9088 8044 9505 8072
rect 9088 8032 9094 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 12802 8032 12808 8084
rect 12860 8032 12866 8084
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 13446 8032 13452 8084
rect 13504 8032 13510 8084
rect 15102 8072 15108 8084
rect 13648 8044 15108 8072
rect 3142 7964 3148 8016
rect 3200 7964 3206 8016
rect 11790 8004 11796 8016
rect 11624 7976 11796 8004
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 7098 7936 7104 7948
rect 4120 7908 7104 7936
rect 4120 7896 4126 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 8110 7936 8116 7948
rect 7699 7908 8116 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 8110 7896 8116 7908
rect 8168 7936 8174 7948
rect 8662 7936 8668 7948
rect 8168 7908 8668 7936
rect 8168 7896 8174 7908
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4387 7840 4752 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4724 7744 4752 7840
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6604 7840 6745 7868
rect 6604 7828 6610 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7834 7868 7840 7880
rect 7423 7840 7840 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 6638 7800 6644 7812
rect 6135 7772 6644 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6748 7800 6776 7831
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7944 7840 8217 7868
rect 7469 7803 7527 7809
rect 7469 7800 7481 7803
rect 6748 7772 7481 7800
rect 7469 7769 7481 7772
rect 7515 7800 7527 7803
rect 7944 7800 7972 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8570 7868 8576 7880
rect 8435 7840 8576 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9180 7840 10241 7868
rect 9180 7828 9186 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10367 7840 10701 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 11624 7877 11652 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 13464 8004 13492 8032
rect 12636 7976 13492 8004
rect 12636 7936 12664 7976
rect 11716 7908 12664 7936
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11716 7858 11744 7908
rect 11793 7861 11851 7867
rect 11793 7858 11805 7861
rect 11716 7830 11805 7858
rect 11793 7827 11805 7830
rect 11839 7827 11851 7861
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11940 7840 12173 7868
rect 11940 7828 11946 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12636 7868 12664 7908
rect 13541 7944 13599 7945
rect 13648 7944 13676 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 15252 8044 17417 8072
rect 15252 8032 15258 8044
rect 17405 8041 17417 8044
rect 17451 8041 17463 8075
rect 17405 8035 17463 8041
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18322 8072 18328 8084
rect 18279 8044 18328 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 13541 7939 13676 7944
rect 13541 7905 13553 7939
rect 13587 7916 13676 7939
rect 14550 7936 14556 7948
rect 13587 7905 13599 7916
rect 13541 7899 13599 7905
rect 13740 7908 14556 7936
rect 12483 7840 12664 7868
rect 12713 7871 12771 7877
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13740 7868 13768 7908
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 17586 7896 17592 7948
rect 17644 7896 17650 7948
rect 13311 7840 13768 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 11793 7821 11851 7827
rect 7515 7772 7972 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 8018 7760 8024 7812
rect 8076 7760 8082 7812
rect 9582 7760 9588 7812
rect 9640 7760 9646 7812
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 12728 7800 12756 7831
rect 14182 7828 14188 7880
rect 14240 7828 14246 7880
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 16172 7840 16497 7868
rect 16172 7828 16178 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 16908 7840 17693 7868
rect 16908 7828 16914 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 17681 7831 17739 7837
rect 17880 7840 18337 7868
rect 12032 7772 12756 7800
rect 13541 7803 13599 7809
rect 12032 7760 12038 7772
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 13587 7772 14473 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 14568 7772 14950 7800
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4614 7732 4620 7744
rect 4295 7704 4620 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 4706 7692 4712 7744
rect 4764 7692 4770 7744
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11112 7704 11621 7732
rect 11112 7692 11118 7704
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 11609 7695 11667 7701
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 11756 7704 12173 7732
rect 11756 7692 11762 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12161 7695 12219 7701
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14568 7732 14596 7772
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 15988 7772 16221 7800
rect 15988 7760 15994 7772
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16209 7763 16267 7769
rect 17880 7744 17908 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 14148 7704 14596 7732
rect 14148 7692 14154 7704
rect 16574 7692 16580 7744
rect 16632 7692 16638 7744
rect 17037 7735 17095 7741
rect 17037 7701 17049 7735
rect 17083 7732 17095 7735
rect 17862 7732 17868 7744
rect 17083 7704 17868 7732
rect 17083 7701 17095 7704
rect 17037 7695 17095 7701
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 1104 7642 18860 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 18860 7642
rect 1104 7568 18860 7590
rect 2746 7500 6684 7528
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 2746 7460 2774 7500
rect 6656 7472 6684 7500
rect 7006 7488 7012 7540
rect 7064 7488 7070 7540
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 10796 7500 12081 7528
rect 1544 7432 2774 7460
rect 1544 7420 1550 7432
rect 1946 7352 1952 7404
rect 2004 7352 2010 7404
rect 2746 7392 2774 7432
rect 3602 7420 3608 7472
rect 3660 7420 3666 7472
rect 5184 7432 6040 7460
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2746 7364 2881 7392
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5184 7401 5212 7432
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4856 7364 5181 7392
rect 4856 7352 4862 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 2774 7324 2780 7336
rect 2547 7296 2780 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 5368 7324 5396 7355
rect 5184 7296 5396 7324
rect 5184 7200 5212 7296
rect 5902 7216 5908 7268
rect 5960 7216 5966 7268
rect 6012 7256 6040 7432
rect 6638 7420 6644 7472
rect 6696 7420 6702 7472
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7024 7392 7052 7488
rect 6779 7364 7052 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6104 7324 6132 7355
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7392 7711 7395
rect 8036 7392 8064 7488
rect 9398 7420 9404 7472
rect 9456 7460 9462 7472
rect 10796 7469 10824 7500
rect 12069 7497 12081 7500
rect 12115 7528 12127 7531
rect 13722 7528 13728 7540
rect 12115 7500 13728 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14182 7528 14188 7540
rect 13832 7500 14188 7528
rect 10781 7463 10839 7469
rect 10781 7460 10793 7463
rect 9456 7432 10793 7460
rect 9456 7420 9462 7432
rect 10781 7429 10793 7432
rect 10827 7429 10839 7463
rect 10781 7423 10839 7429
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 11698 7460 11704 7472
rect 10928 7432 11704 7460
rect 10928 7420 10934 7432
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 13354 7460 13360 7472
rect 11940 7432 12664 7460
rect 11940 7420 11946 7432
rect 7699 7364 8064 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 6914 7324 6920 7336
rect 6104 7296 6920 7324
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7392 7256 7420 7355
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10888 7392 10916 7420
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 10643 7364 10916 7392
rect 11716 7364 11989 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10226 7284 10232 7336
rect 10284 7324 10290 7336
rect 10612 7324 10640 7355
rect 10284 7296 10640 7324
rect 10284 7284 10290 7296
rect 6012 7228 7420 7256
rect 8938 7216 8944 7268
rect 8996 7216 9002 7268
rect 11716 7256 11744 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12636 7401 12664 7432
rect 13188 7432 13360 7460
rect 13188 7401 13216 7432
rect 13354 7420 13360 7432
rect 13412 7460 13418 7472
rect 13832 7460 13860 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 14424 7500 14780 7528
rect 14424 7488 14430 7500
rect 13412 7432 13860 7460
rect 13412 7420 13418 7432
rect 14090 7420 14096 7472
rect 14148 7420 14154 7472
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 12124 7364 12173 7392
rect 12124 7352 12130 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 13173 7395 13231 7401
rect 12667 7364 13124 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12986 7256 12992 7268
rect 11716 7228 12992 7256
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7188 4675 7191
rect 4706 7188 4712 7200
rect 4663 7160 4712 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 6914 7188 6920 7200
rect 6687 7160 6920 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 7064 7160 7205 7188
rect 7064 7148 7070 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 10686 7148 10692 7200
rect 10744 7148 10750 7200
rect 12713 7191 12771 7197
rect 12713 7157 12725 7191
rect 12759 7188 12771 7191
rect 12802 7188 12808 7200
rect 12759 7160 12808 7188
rect 12759 7157 12771 7160
rect 12713 7151 12771 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13096 7188 13124 7364
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7324 13507 7327
rect 13538 7324 13544 7336
rect 13495 7296 13544 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 14752 7324 14780 7500
rect 15010 7488 15016 7540
rect 15068 7488 15074 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15746 7528 15752 7540
rect 15611 7500 15752 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 16632 7500 16988 7528
rect 16632 7488 16638 7500
rect 15028 7392 15056 7488
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 16071 7432 16804 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15028 7364 15485 7392
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15930 7352 15936 7404
rect 15988 7352 15994 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16776 7401 16804 7432
rect 16850 7420 16856 7472
rect 16908 7420 16914 7472
rect 16960 7401 16988 7500
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 18012 7500 18061 7528
rect 18012 7488 18018 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17092 7364 17417 7392
rect 17092 7352 17098 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 15194 7324 15200 7336
rect 14752 7296 15200 7324
rect 14752 7188 14780 7296
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 17604 7324 17632 7355
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 16080 7296 17632 7324
rect 16080 7284 16086 7296
rect 13096 7160 14780 7188
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 17954 7188 17960 7200
rect 17543 7160 17960 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 1104 7098 18860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 18860 7098
rect 1104 7024 18860 7046
rect 1946 6944 1952 6996
rect 2004 6944 2010 6996
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 3200 6956 3985 6984
rect 3200 6944 3206 6956
rect 3973 6953 3985 6956
rect 4019 6953 4031 6987
rect 3973 6947 4031 6953
rect 4065 6987 4123 6993
rect 4065 6953 4077 6987
rect 4111 6984 4123 6987
rect 4798 6984 4804 6996
rect 4111 6956 4804 6984
rect 4111 6953 4123 6956
rect 4065 6947 4123 6953
rect 4080 6916 4108 6947
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 5258 6984 5264 6996
rect 4908 6956 5264 6984
rect 3804 6888 4108 6916
rect 3804 6860 3832 6888
rect 2590 6808 2596 6860
rect 2648 6808 2654 6860
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 3786 6848 3792 6860
rect 2823 6820 3792 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4908 6848 4936 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 6904 6987 6962 6993
rect 6904 6953 6916 6987
rect 6950 6984 6962 6987
rect 7006 6984 7012 6996
rect 6950 6956 7012 6984
rect 6950 6953 6962 6956
rect 6904 6947 6962 6953
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 13265 6987 13323 6993
rect 13265 6953 13277 6987
rect 13311 6984 13323 6987
rect 13538 6984 13544 6996
rect 13311 6956 13544 6984
rect 13311 6953 13323 6956
rect 13265 6947 13323 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 15013 6987 15071 6993
rect 15013 6953 15025 6987
rect 15059 6984 15071 6987
rect 16022 6984 16028 6996
rect 15059 6956 16028 6984
rect 15059 6953 15071 6956
rect 15013 6947 15071 6953
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 16853 6987 16911 6993
rect 16853 6953 16865 6987
rect 16899 6984 16911 6987
rect 17586 6984 17592 6996
rect 16899 6956 17592 6984
rect 16899 6953 16911 6956
rect 16853 6947 16911 6953
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 4985 6919 5043 6925
rect 4985 6885 4997 6919
rect 5031 6916 5043 6919
rect 6546 6916 6552 6928
rect 5031 6888 6552 6916
rect 5031 6885 5043 6888
rect 4985 6879 5043 6885
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 10100 6888 12664 6916
rect 10100 6876 10106 6888
rect 3927 6820 4936 6848
rect 6273 6851 6331 6857
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 6362 6848 6368 6860
rect 6319 6820 6368 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6638 6808 6644 6860
rect 6696 6808 6702 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7650 6848 7656 6860
rect 6972 6820 7656 6848
rect 6972 6808 6978 6820
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 2958 6780 2964 6792
rect 2915 6752 2964 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 2148 6712 2176 6743
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4614 6780 4620 6792
rect 4203 6752 4620 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6749 4951 6783
rect 5077 6785 5135 6791
rect 5077 6780 5089 6785
rect 4893 6743 4951 6749
rect 5000 6752 5089 6780
rect 2148 6684 2774 6712
rect 1762 6604 1768 6656
rect 1820 6644 1826 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 1820 6616 2605 6644
rect 1820 6604 1826 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2746 6644 2774 6684
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4525 6715 4583 6721
rect 4525 6712 4537 6715
rect 3936 6684 4537 6712
rect 3936 6672 3942 6684
rect 4525 6681 4537 6684
rect 4571 6712 4583 6715
rect 4908 6712 4936 6743
rect 5000 6724 5028 6752
rect 5077 6751 5089 6752
rect 5123 6780 5135 6785
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5123 6752 5733 6780
rect 5123 6751 5135 6752
rect 5077 6745 5135 6751
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 10060 6780 10088 6876
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10226 6848 10232 6860
rect 10183 6820 10232 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 11698 6848 11704 6860
rect 10336 6820 11704 6848
rect 10336 6789 10364 6820
rect 11698 6808 11704 6820
rect 11756 6848 11762 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 11756 6820 11897 6848
rect 11756 6808 11762 6820
rect 11885 6817 11897 6820
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 12636 6792 12664 6888
rect 12802 6876 12808 6928
rect 12860 6916 12866 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 12860 6888 13185 6916
rect 12860 6876 12866 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 17773 6919 17831 6925
rect 17773 6916 17785 6919
rect 13173 6879 13231 6885
rect 14568 6888 17785 6916
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 9815 6752 10088 6780
rect 10321 6783 10379 6789
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10594 6780 10600 6792
rect 10551 6752 10600 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10744 6752 10793 6780
rect 10744 6740 10750 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 4571 6684 4936 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 4982 6672 4988 6724
rect 5040 6672 5046 6724
rect 7374 6712 7380 6724
rect 7208 6684 7380 6712
rect 2866 6644 2872 6656
rect 2746 6616 2872 6644
rect 2593 6607 2651 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 3660 6616 5365 6644
rect 3660 6604 3666 6616
rect 5353 6613 5365 6616
rect 5399 6644 5411 6647
rect 7208 6644 7236 6684
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 9858 6672 9864 6724
rect 9916 6712 9922 6724
rect 10873 6715 10931 6721
rect 10873 6712 10885 6715
rect 9916 6684 10885 6712
rect 9916 6672 9922 6684
rect 10873 6681 10885 6684
rect 10919 6681 10931 6715
rect 10873 6675 10931 6681
rect 10980 6656 11008 6743
rect 11992 6712 12020 6743
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 12820 6789 12848 6876
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 13403 6820 14473 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 14568 6789 14596 6888
rect 17773 6885 17785 6888
rect 17819 6885 17831 6919
rect 17773 6879 17831 6885
rect 14642 6808 14648 6860
rect 14700 6808 14706 6860
rect 16942 6808 16948 6860
rect 17000 6808 17006 6860
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13136 6752 14381 6780
rect 13136 6740 13142 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 12066 6712 12072 6724
rect 11992 6684 12072 6712
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 14384 6712 14412 6743
rect 14660 6712 14688 6808
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 14384 6684 14688 6712
rect 15120 6712 15148 6743
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15252 6752 15393 6780
rect 15252 6740 15258 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 16114 6780 16120 6792
rect 15620 6752 16120 6780
rect 15620 6740 15626 6752
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 16758 6740 16764 6792
rect 16816 6740 16822 6792
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18012 6752 18153 6780
rect 18012 6740 18018 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 15120 6684 15516 6712
rect 5399 6616 7236 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 7340 6616 8401 6644
rect 7340 6604 7346 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8628 6616 9045 6644
rect 8628 6604 8634 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 9950 6644 9956 6656
rect 9723 6616 9956 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10962 6604 10968 6656
rect 11020 6604 11026 6656
rect 15488 6653 15516 6684
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 15930 6644 15936 6656
rect 15519 6616 15936 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 1104 6554 18860 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 18860 6554
rect 1104 6480 18860 6502
rect 3602 6400 3608 6452
rect 3660 6400 3666 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 7282 6440 7288 6452
rect 5224 6412 7288 6440
rect 5224 6400 5230 6412
rect 1762 6332 1768 6384
rect 1820 6332 1826 6384
rect 3620 6372 3648 6400
rect 7208 6381 7236 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 8570 6440 8576 6452
rect 7432 6412 8576 6440
rect 7432 6400 7438 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 11848 6412 11928 6440
rect 11848 6400 11854 6412
rect 11900 6381 11928 6412
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 16301 6443 16359 6449
rect 12124 6412 13676 6440
rect 12124 6400 12130 6412
rect 13648 6381 13676 6412
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 16942 6440 16948 6452
rect 16347 6412 16948 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17405 6443 17463 6449
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 18046 6440 18052 6452
rect 17451 6412 18052 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 2990 6358 3648 6372
rect 2976 6344 3648 6358
rect 5813 6375 5871 6381
rect 1486 6196 1492 6248
rect 1544 6196 1550 6248
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 2976 6236 3004 6344
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 7193 6375 7251 6381
rect 5859 6344 7144 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 4062 6264 4068 6316
rect 4120 6264 4126 6316
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 5675 6276 6469 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 2464 6208 3004 6236
rect 2464 6196 2470 6208
rect 4706 6196 4712 6248
rect 4764 6196 4770 6248
rect 3970 6168 3976 6180
rect 3160 6140 3976 6168
rect 2498 6060 2504 6112
rect 2556 6100 2562 6112
rect 3160 6100 3188 6140
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 5166 6168 5172 6180
rect 4295 6140 5172 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 5261 6171 5319 6177
rect 5261 6137 5273 6171
rect 5307 6168 5319 6171
rect 5644 6168 5672 6267
rect 6638 6264 6644 6316
rect 6696 6264 6702 6316
rect 7116 6304 7144 6344
rect 7193 6341 7205 6375
rect 7239 6341 7251 6375
rect 11885 6375 11943 6381
rect 7193 6335 7251 6341
rect 7300 6344 10824 6372
rect 7300 6304 7328 6344
rect 7116 6276 7328 6304
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 7484 6236 7512 6267
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7708 6276 7849 6304
rect 7708 6264 7714 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 5951 6208 6408 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 5307 6140 5672 6168
rect 5307 6137 5319 6140
rect 5261 6131 5319 6137
rect 6380 6112 6408 6208
rect 6472 6208 7512 6236
rect 6472 6112 6500 6208
rect 7190 6128 7196 6180
rect 7248 6128 7254 6180
rect 7852 6168 7880 6267
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 9048 6313 9076 6344
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9447 6276 9965 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10410 6264 10416 6316
rect 10468 6264 10474 6316
rect 10796 6313 10824 6344
rect 11885 6341 11897 6375
rect 11931 6341 11943 6375
rect 11885 6335 11943 6341
rect 13633 6375 13691 6381
rect 13633 6341 13645 6375
rect 13679 6372 13691 6375
rect 14737 6375 14795 6381
rect 13679 6344 14688 6372
rect 13679 6341 13691 6344
rect 13633 6335 13691 6341
rect 14660 6316 14688 6344
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 14783 6344 17448 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 14090 6304 14096 6316
rect 13044 6276 14096 6304
rect 13044 6264 13050 6276
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14752 6276 14841 6304
rect 10275 6239 10333 6245
rect 10275 6205 10287 6239
rect 10321 6236 10333 6239
rect 11054 6236 11060 6248
rect 10321 6208 11060 6236
rect 10321 6205 10333 6208
rect 10275 6199 10333 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11296 6208 11621 6236
rect 11296 6196 11302 6208
rect 11609 6205 11621 6208
rect 11655 6236 11667 6239
rect 13354 6236 13360 6248
rect 11655 6208 13360 6236
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 10870 6168 10876 6180
rect 7852 6140 10876 6168
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 14752 6168 14780 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15252 6276 15301 6304
rect 15252 6264 15258 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15562 6304 15568 6316
rect 15519 6276 15568 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15286 6168 15292 6180
rect 14752 6140 15292 6168
rect 2556 6072 3188 6100
rect 2556 6060 2562 6072
rect 3234 6060 3240 6112
rect 3292 6060 3298 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 4798 6100 4804 6112
rect 3927 6072 4804 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 6362 6060 6368 6112
rect 6420 6060 6426 6112
rect 6454 6060 6460 6112
rect 6512 6060 6518 6112
rect 6641 6103 6699 6109
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 7926 6100 7932 6112
rect 6687 6072 7932 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 10042 6060 10048 6112
rect 10100 6060 10106 6112
rect 10134 6060 10140 6112
rect 10192 6060 10198 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 12618 6100 12624 6112
rect 11020 6072 12624 6100
rect 11020 6060 11026 6072
rect 12618 6060 12624 6072
rect 12676 6100 12682 6112
rect 14752 6100 14780 6140
rect 15286 6128 15292 6140
rect 15344 6168 15350 6180
rect 15488 6168 15516 6267
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 16132 6313 16160 6344
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 15933 6239 15991 6245
rect 15933 6205 15945 6239
rect 15979 6236 15991 6239
rect 17052 6236 17080 6264
rect 17420 6248 17448 6344
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17957 6307 18015 6313
rect 17957 6304 17969 6307
rect 17727 6276 17969 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 17957 6273 17969 6276
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 15979 6208 17080 6236
rect 15979 6205 15991 6208
rect 15933 6199 15991 6205
rect 15344 6140 15516 6168
rect 15344 6128 15350 6140
rect 12676 6072 14780 6100
rect 15381 6103 15439 6109
rect 12676 6060 12682 6072
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15948 6100 15976 6199
rect 17402 6196 17408 6248
rect 17460 6196 17466 6248
rect 17696 6168 17724 6267
rect 16132 6140 17724 6168
rect 16132 6112 16160 6140
rect 15427 6072 15976 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 16114 6060 16120 6112
rect 16172 6060 16178 6112
rect 16758 6060 16764 6112
rect 16816 6100 16822 6112
rect 17586 6100 17592 6112
rect 16816 6072 17592 6100
rect 16816 6060 16822 6072
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17828 6072 18061 6100
rect 17828 6060 17834 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 1104 6010 18860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 18860 6010
rect 1104 5936 18860 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 4062 5896 4068 5908
rect 1811 5868 4068 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 6362 5856 6368 5908
rect 6420 5856 6426 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6696 5868 7021 5896
rect 6696 5856 6702 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 7282 5856 7288 5908
rect 7340 5856 7346 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7708 5868 7849 5896
rect 7708 5856 7714 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 7926 5856 7932 5908
rect 7984 5856 7990 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9214 5896 9220 5908
rect 9171 5868 9220 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 10042 5856 10048 5908
rect 10100 5856 10106 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 11698 5856 11704 5908
rect 11756 5856 11762 5908
rect 11790 5856 11796 5908
rect 11848 5856 11854 5908
rect 12820 5868 16252 5896
rect 2498 5788 2504 5840
rect 2556 5788 2562 5840
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 4157 5831 4215 5837
rect 4157 5828 4169 5831
rect 2648 5800 4169 5828
rect 2648 5788 2654 5800
rect 4157 5797 4169 5800
rect 4203 5797 4215 5831
rect 6454 5828 6460 5840
rect 4157 5791 4215 5797
rect 4632 5800 6460 5828
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 1360 5732 1716 5760
rect 1360 5720 1366 5732
rect 1688 5704 1716 5732
rect 3234 5720 3240 5772
rect 3292 5720 3298 5772
rect 3786 5720 3792 5772
rect 3844 5720 3850 5772
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4028 5732 4292 5760
rect 4028 5720 4034 5732
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 2774 5652 2780 5704
rect 2832 5652 2838 5704
rect 3804 5692 3832 5720
rect 4264 5701 4292 5732
rect 4632 5704 4660 5800
rect 6454 5788 6460 5800
rect 6512 5828 6518 5840
rect 6512 5800 7236 5828
rect 6512 5788 6518 5800
rect 4798 5720 4804 5772
rect 4856 5720 4862 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5307 5732 7144 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3804 5664 4077 5692
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4614 5692 4620 5704
rect 4295 5664 4620 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4890 5692 4896 5704
rect 4724 5664 4896 5692
rect 4724 5624 4752 5664
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 6656 5701 6684 5732
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7116 5701 7144 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 3528 5596 4752 5624
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 3418 5556 3424 5568
rect 2179 5528 3424 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3528 5565 3556 5596
rect 6362 5584 6368 5636
rect 6420 5584 6426 5636
rect 7208 5624 7236 5800
rect 7300 5760 7328 5856
rect 7944 5760 7972 5856
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 9766 5828 9772 5840
rect 8076 5800 9772 5828
rect 8076 5788 8082 5800
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 10060 5760 10088 5856
rect 7300 5732 7696 5760
rect 7944 5732 9076 5760
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7668 5692 7696 5732
rect 9048 5701 9076 5732
rect 9692 5732 10088 5760
rect 11885 5763 11943 5769
rect 9692 5701 9720 5732
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 11931 5732 12725 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7668 5664 8125 5692
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 7837 5627 7895 5633
rect 7208 5596 7788 5624
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5525 3571 5559
rect 3513 5519 3571 5525
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 5684 5528 6561 5556
rect 5684 5516 5690 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7524 5528 7665 5556
rect 7524 5516 7530 5528
rect 7653 5525 7665 5528
rect 7699 5525 7711 5559
rect 7760 5556 7788 5596
rect 7837 5593 7849 5627
rect 7883 5624 7895 5627
rect 7926 5624 7932 5636
rect 7883 5596 7932 5624
rect 7883 5593 7895 5596
rect 7837 5587 7895 5593
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 8312 5624 8340 5655
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 10008 5664 10149 5692
rect 10008 5652 10014 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 12820 5701 12848 5868
rect 14642 5788 14648 5840
rect 14700 5788 14706 5840
rect 15286 5788 15292 5840
rect 15344 5788 15350 5840
rect 15473 5831 15531 5837
rect 15473 5797 15485 5831
rect 15519 5828 15531 5831
rect 16114 5828 16120 5840
rect 15519 5800 16120 5828
rect 15519 5797 15531 5800
rect 15473 5791 15531 5797
rect 16114 5788 16120 5800
rect 16172 5788 16178 5840
rect 13078 5720 13084 5772
rect 13136 5720 13142 5772
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11664 5664 12633 5692
rect 11664 5652 11670 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 9122 5624 9128 5636
rect 8036 5596 9128 5624
rect 8036 5556 8064 5596
rect 9122 5584 9128 5596
rect 9180 5584 9186 5636
rect 10226 5584 10232 5636
rect 10284 5584 10290 5636
rect 10413 5627 10471 5633
rect 10413 5593 10425 5627
rect 10459 5624 10471 5627
rect 10594 5624 10600 5636
rect 10459 5596 10600 5624
rect 10459 5593 10471 5596
rect 10413 5587 10471 5593
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 12636 5624 12664 5655
rect 13096 5624 13124 5720
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 13228 5664 13277 5692
rect 13228 5652 13234 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 14660 5692 14688 5788
rect 15304 5760 15332 5788
rect 15304 5732 15516 5760
rect 15488 5701 15516 5732
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14660 5664 15301 5692
rect 13265 5655 13323 5661
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 12636 5596 13124 5624
rect 13280 5624 13308 5655
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16132 5701 16160 5788
rect 16224 5760 16252 5868
rect 16666 5856 16672 5908
rect 16724 5856 16730 5908
rect 17586 5856 17592 5908
rect 17644 5856 17650 5908
rect 17604 5828 17632 5856
rect 17604 5800 18000 5828
rect 17972 5769 18000 5800
rect 17681 5763 17739 5769
rect 17681 5760 17693 5763
rect 16224 5732 17693 5760
rect 17681 5729 17693 5732
rect 17727 5729 17739 5763
rect 17681 5723 17739 5729
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 15378 5624 15384 5636
rect 13280 5596 15384 5624
rect 15378 5584 15384 5596
rect 15436 5584 15442 5636
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5624 16083 5627
rect 16592 5624 16620 5655
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 18049 5695 18107 5701
rect 18049 5692 18061 5695
rect 17644 5664 18061 5692
rect 17644 5652 17650 5664
rect 18049 5661 18061 5664
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 16071 5596 16620 5624
rect 16071 5593 16083 5596
rect 16025 5587 16083 5593
rect 7760 5528 8064 5556
rect 7653 5519 7711 5525
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 9861 5559 9919 5565
rect 9861 5525 9873 5559
rect 9907 5556 9919 5559
rect 10318 5556 10324 5568
rect 9907 5528 10324 5556
rect 9907 5525 9919 5528
rect 9861 5519 9919 5525
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 13170 5516 13176 5568
rect 13228 5516 13234 5568
rect 1104 5466 18860 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 18860 5466
rect 1104 5392 18860 5414
rect 1670 5312 1676 5364
rect 1728 5312 1734 5364
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 2774 5352 2780 5364
rect 1903 5324 2780 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 2958 5312 2964 5364
rect 3016 5312 3022 5364
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 4614 5312 4620 5364
rect 4672 5312 4678 5364
rect 4890 5312 4896 5364
rect 4948 5312 4954 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 6362 5352 6368 5364
rect 5583 5324 6368 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 8628 5324 8800 5352
rect 8628 5312 8634 5324
rect 1688 5284 1716 5312
rect 2225 5287 2283 5293
rect 2225 5284 2237 5287
rect 1688 5256 2237 5284
rect 2225 5253 2237 5256
rect 2271 5253 2283 5287
rect 2225 5247 2283 5253
rect 1118 5176 1124 5228
rect 1176 5216 1182 5228
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1176 5188 1777 5216
rect 1176 5176 1182 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3252 5216 3280 5312
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 3878 5284 3884 5296
rect 3476 5256 3884 5284
rect 3476 5244 3482 5256
rect 3878 5244 3884 5256
rect 3936 5284 3942 5296
rect 3936 5256 4200 5284
rect 3936 5244 3942 5256
rect 3099 5188 3280 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 4172 5225 4200 5256
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3660 5188 3985 5216
rect 3660 5176 3666 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4632 5216 4660 5312
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4632 5188 4721 5216
rect 4157 5179 4215 5185
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 4908 5216 4936 5312
rect 5997 5287 6055 5293
rect 5997 5253 6009 5287
rect 6043 5284 6055 5287
rect 7392 5284 7420 5312
rect 6043 5256 7420 5284
rect 6043 5253 6055 5256
rect 5997 5247 6055 5253
rect 7650 5244 7656 5296
rect 7708 5244 7714 5296
rect 8772 5228 8800 5324
rect 9122 5312 9128 5364
rect 9180 5312 9186 5364
rect 10226 5352 10232 5364
rect 10060 5324 10232 5352
rect 10060 5293 10088 5324
rect 10226 5312 10232 5324
rect 10284 5352 10290 5364
rect 13998 5352 14004 5364
rect 10284 5324 14004 5352
rect 10284 5312 10290 5324
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 16758 5352 16764 5364
rect 16255 5324 16764 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 17402 5312 17408 5364
rect 17460 5312 17466 5364
rect 17586 5312 17592 5364
rect 17644 5312 17650 5364
rect 17770 5312 17776 5364
rect 17828 5312 17834 5364
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5253 10103 5287
rect 10045 5247 10103 5253
rect 11440 5256 12480 5284
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4908 5188 5365 5216
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7006 5216 7012 5228
rect 6963 5188 7012 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 4816 5148 4844 5176
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4816 5120 5181 5148
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 6104 5080 6132 5179
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7282 5216 7288 5228
rect 7147 5188 7288 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 8754 5176 8760 5228
rect 8812 5176 8818 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10226 5216 10232 5228
rect 9815 5188 10232 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10594 5216 10600 5228
rect 10367 5188 10600 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 10594 5176 10600 5188
rect 10652 5216 10658 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10652 5188 10977 5216
rect 10652 5176 10658 5188
rect 10965 5185 10977 5188
rect 11011 5216 11023 5219
rect 11440 5216 11468 5256
rect 11011 5188 11560 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11532 5160 11560 5188
rect 11606 5176 11612 5228
rect 11664 5206 11670 5228
rect 12452 5225 12480 5256
rect 14090 5244 14096 5296
rect 14148 5244 14154 5296
rect 15378 5244 15384 5296
rect 15436 5244 15442 5296
rect 12437 5219 12495 5225
rect 11664 5178 11699 5206
rect 12437 5185 12449 5219
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 12621 5219 12679 5225
rect 12621 5185 12633 5219
rect 12667 5216 12679 5219
rect 12710 5216 12716 5228
rect 12667 5188 12716 5216
rect 12667 5185 12679 5188
rect 12621 5179 12679 5185
rect 11664 5176 11670 5178
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13354 5176 13360 5228
rect 13412 5176 13418 5228
rect 15396 5216 15424 5244
rect 15396 5188 15884 5216
rect 11610 5175 11622 5176
rect 11656 5175 11668 5176
rect 11610 5169 11668 5175
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6696 5120 7389 5148
rect 6696 5108 6702 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 10410 5148 10416 5160
rect 9723 5120 10416 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 10410 5108 10416 5120
rect 10468 5148 10474 5160
rect 10468 5120 11468 5148
rect 10468 5108 10474 5120
rect 11440 5092 11468 5120
rect 11514 5108 11520 5160
rect 11572 5108 11578 5160
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 11974 5148 11980 5160
rect 11931 5120 11980 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 13630 5108 13636 5160
rect 13688 5108 13694 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 14240 5120 15761 5148
rect 14240 5108 14246 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15856 5148 15884 5188
rect 15930 5176 15936 5228
rect 15988 5176 15994 5228
rect 17420 5225 17448 5312
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16040 5188 16773 5216
rect 16040 5148 16068 5188
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17589 5219 17647 5225
rect 17589 5185 17601 5219
rect 17635 5216 17647 5219
rect 17788 5216 17816 5312
rect 17635 5188 17816 5216
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 15856 5120 16068 5148
rect 15749 5111 15807 5117
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16301 5151 16359 5157
rect 16301 5148 16313 5151
rect 16172 5120 16313 5148
rect 16172 5108 16178 5120
rect 16301 5117 16313 5120
rect 16347 5117 16359 5151
rect 16301 5111 16359 5117
rect 7190 5080 7196 5092
rect 6104 5052 7196 5080
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10502 5080 10508 5092
rect 10367 5052 10508 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 11422 5040 11428 5092
rect 11480 5040 11486 5092
rect 16022 5040 16028 5092
rect 16080 5080 16086 5092
rect 16960 5080 16988 5179
rect 16080 5052 16988 5080
rect 16080 5040 16086 5052
rect 4062 4972 4068 5024
rect 4120 4972 4126 5024
rect 4798 4972 4804 5024
rect 4856 4972 4862 5024
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 7466 5012 7472 5024
rect 6963 4984 7472 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 9364 4984 10609 5012
rect 9364 4972 9370 4984
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11103 4984 11713 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11790 4972 11796 5024
rect 11848 4972 11854 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12066 5012 12072 5024
rect 11940 4984 12072 5012
rect 11940 4972 11946 4984
rect 12066 4972 12072 4984
rect 12124 5012 12130 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12124 4984 12633 5012
rect 12124 4972 12130 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 16850 4972 16856 5024
rect 16908 4972 16914 5024
rect 1104 4922 18860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 18860 4922
rect 1104 4848 18860 4870
rect 1118 4768 1124 4820
rect 1176 4808 1182 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1176 4780 1593 4808
rect 1176 4768 1182 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 3786 4768 3792 4820
rect 3844 4768 3850 4820
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 6273 4811 6331 4817
rect 4856 4780 6224 4808
rect 4856 4768 4862 4780
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 3804 4672 3832 4768
rect 2924 4644 3832 4672
rect 2924 4632 2930 4644
rect 3252 4613 3280 4644
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3936 4644 3985 4672
rect 3936 4632 3942 4644
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 4080 4672 4108 4768
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 4479 4712 5856 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 5537 4675 5595 4681
rect 5537 4672 5549 4675
rect 4080 4644 5549 4672
rect 3973 4635 4031 4641
rect 5537 4641 5549 4644
rect 5583 4641 5595 4675
rect 5537 4635 5595 4641
rect 5626 4632 5632 4684
rect 5684 4632 5690 4684
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3237 4607 3295 4613
rect 2823 4576 3096 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3068 4480 3096 4576
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3660 4576 4077 4604
rect 3660 4564 3666 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 5537 4539 5595 4545
rect 5537 4505 5549 4539
rect 5583 4536 5595 4539
rect 5644 4536 5672 4632
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 5828 4613 5856 4712
rect 6196 4672 6224 4780
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 6914 4808 6920 4820
rect 6319 4780 6920 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 7558 4808 7564 4820
rect 7331 4780 7564 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8662 4808 8668 4820
rect 8527 4780 8668 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 10502 4808 10508 4820
rect 9171 4780 10508 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10615 4811 10673 4817
rect 10615 4777 10627 4811
rect 10661 4808 10673 4811
rect 11790 4808 11796 4820
rect 10661 4780 11796 4808
rect 10661 4777 10673 4780
rect 10615 4771 10673 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 13170 4808 13176 4820
rect 12406 4780 13176 4808
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 12406 4740 12434 4780
rect 13170 4768 13176 4780
rect 13228 4808 13234 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 13228 4780 13369 4808
rect 13228 4768 13234 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 13357 4771 13415 4777
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 13630 4808 13636 4820
rect 13495 4780 13636 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13998 4768 14004 4820
rect 14056 4768 14062 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 14700 4780 15056 4808
rect 14700 4768 14706 4780
rect 6696 4712 9628 4740
rect 6696 4700 6702 4712
rect 7101 4675 7159 4681
rect 6196 4644 6408 4672
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4604 5871 4607
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5859 4576 6101 4604
rect 5859 4573 5871 4576
rect 5813 4567 5871 4573
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 6380 4604 6408 4644
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 6982 4607 7040 4613
rect 6982 4604 6994 4607
rect 6380 4576 6994 4604
rect 6982 4573 6994 4576
rect 7028 4573 7040 4607
rect 7116 4604 7144 4635
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7340 4644 8033 4672
rect 7340 4632 7346 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 9600 4672 9628 4712
rect 11164 4712 12434 4740
rect 10873 4675 10931 4681
rect 10873 4672 10885 4675
rect 9600 4644 10885 4672
rect 8021 4635 8079 4641
rect 10873 4641 10885 4644
rect 10919 4672 10931 4675
rect 11054 4672 11060 4684
rect 10919 4644 11060 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 7190 4604 7196 4616
rect 7116 4576 7196 4604
rect 6982 4567 7040 4573
rect 7190 4564 7196 4576
rect 7248 4604 7254 4616
rect 7926 4604 7932 4616
rect 7248 4576 7932 4604
rect 7248 4564 7254 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 5583 4508 5672 4536
rect 8588 4536 8616 4567
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9306 4604 9312 4616
rect 8812 4576 9312 4604
rect 8812 4564 8818 4576
rect 9306 4564 9312 4576
rect 9364 4604 9370 4616
rect 9364 4576 9522 4604
rect 9364 4564 9370 4576
rect 8588 4508 9352 4536
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 2648 4440 2697 4468
rect 2648 4428 2654 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 2685 4431 2743 4437
rect 3050 4428 3056 4480
rect 3108 4428 3114 4480
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 9324 4468 9352 4508
rect 11164 4468 11192 4712
rect 13078 4700 13084 4752
rect 13136 4700 13142 4752
rect 14016 4740 14044 4768
rect 14550 4740 14556 4752
rect 14016 4712 14556 4740
rect 14550 4700 14556 4712
rect 14608 4740 14614 4752
rect 14608 4712 14872 4740
rect 14608 4700 14614 4712
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12207 4644 12664 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11348 4536 11376 4567
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11790 4604 11796 4616
rect 11480 4576 11796 4604
rect 11480 4564 11486 4576
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 11900 4604 11928 4635
rect 11900 4576 12572 4604
rect 11882 4536 11888 4548
rect 11348 4508 11888 4536
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 9324 4440 11192 4468
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 12544 4468 12572 4576
rect 12636 4548 12664 4644
rect 13096 4604 13124 4700
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 14461 4675 14519 4681
rect 14461 4672 14473 4675
rect 13587 4644 14473 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 14461 4641 14473 4644
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 13096 4576 13277 4604
rect 13265 4573 13277 4576
rect 13311 4604 13323 4607
rect 14366 4604 14372 4616
rect 13311 4576 14372 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14844 4613 14872 4712
rect 15028 4672 15056 4780
rect 16022 4672 16028 4684
rect 15028 4644 16028 4672
rect 15028 4613 15056 4644
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 12618 4496 12624 4548
rect 12676 4496 12682 4548
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 14568 4536 14596 4567
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15764 4613 15792 4644
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 17310 4632 17316 4684
rect 17368 4632 17374 4684
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17420 4644 17969 4672
rect 15565 4607 15623 4613
rect 15565 4604 15577 4607
rect 15436 4576 15577 4604
rect 15436 4564 15442 4576
rect 15565 4573 15577 4576
rect 15611 4573 15623 4607
rect 15565 4567 15623 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 16850 4564 16856 4616
rect 16908 4604 16914 4616
rect 17420 4613 17448 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 17405 4607 17463 4613
rect 16908 4576 17356 4604
rect 16908 4564 16914 4576
rect 17328 4536 17356 4576
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17862 4564 17868 4616
rect 17920 4564 17926 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18064 4536 18092 4567
rect 12768 4508 14504 4536
rect 14568 4508 17080 4536
rect 17328 4508 18092 4536
rect 12768 4496 12774 4508
rect 13170 4468 13176 4480
rect 12544 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14476 4468 14504 4508
rect 14642 4468 14648 4480
rect 14476 4440 14648 4468
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 14918 4428 14924 4480
rect 14976 4428 14982 4480
rect 15654 4428 15660 4480
rect 15712 4428 15718 4480
rect 17052 4477 17080 4508
rect 17037 4471 17095 4477
rect 17037 4437 17049 4471
rect 17083 4437 17095 4471
rect 17037 4431 17095 4437
rect 1104 4378 18860 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 18860 4378
rect 1104 4304 18860 4326
rect 3602 4224 3608 4276
rect 3660 4224 3666 4276
rect 7926 4224 7932 4276
rect 7984 4224 7990 4276
rect 11149 4267 11207 4273
rect 11149 4233 11161 4267
rect 11195 4264 11207 4267
rect 11606 4264 11612 4276
rect 11195 4236 11612 4264
rect 11195 4233 11207 4236
rect 11149 4227 11207 4233
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 14182 4264 14188 4276
rect 12268 4236 14188 4264
rect 2406 4156 2412 4208
rect 2464 4156 2470 4208
rect 7837 4199 7895 4205
rect 5184 4168 6868 4196
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3200 4100 3818 4128
rect 3200 4088 3206 4100
rect 1486 4020 1492 4072
rect 1544 4020 1550 4072
rect 1762 4020 1768 4072
rect 1820 4020 1826 4072
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3108 4032 3249 4060
rect 3108 4020 3114 4032
rect 3237 4029 3249 4032
rect 3283 4060 3295 4063
rect 3283 4032 3910 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 1504 3924 1532 4020
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 4617 3995 4675 4001
rect 4617 3992 4629 3995
rect 3476 3964 4629 3992
rect 3476 3952 3482 3964
rect 4617 3961 4629 3964
rect 4663 3992 4675 3995
rect 5184 3992 5212 4168
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5442 4128 5448 4140
rect 5399 4100 5448 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5276 4060 5304 4091
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5583 4100 6469 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6840 4128 6868 4168
rect 7392 4168 7696 4196
rect 7392 4128 7420 4168
rect 6687 4100 6776 4128
rect 6840 4100 7420 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 5276 4032 5396 4060
rect 5368 4004 5396 4032
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 4663 3964 5212 3992
rect 4663 3961 4675 3964
rect 4617 3955 4675 3961
rect 5350 3952 5356 4004
rect 5408 3952 5414 4004
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 5736 3992 5764 4020
rect 6748 4004 6776 4100
rect 7466 4088 7472 4140
rect 7524 4088 7530 4140
rect 7668 4128 7696 4168
rect 7837 4165 7849 4199
rect 7883 4196 7895 4199
rect 7944 4196 7972 4224
rect 7883 4168 8432 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 8110 4128 8116 4140
rect 7668 4100 8116 4128
rect 8110 4088 8116 4100
rect 8168 4128 8174 4140
rect 8404 4137 8432 4168
rect 10226 4156 10232 4208
rect 10284 4196 10290 4208
rect 10284 4168 10548 4196
rect 10284 4156 10290 4168
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8168 4100 8309 4128
rect 8168 4088 8174 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8570 4088 8576 4140
rect 8628 4088 8634 4140
rect 8662 4088 8668 4140
rect 8720 4088 8726 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 6822 4020 6828 4072
rect 6880 4020 6886 4072
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7064 4032 7389 4060
rect 7064 4020 7070 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 7742 4020 7748 4072
rect 7800 4020 7806 4072
rect 8588 4060 8616 4088
rect 8772 4060 8800 4091
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 10520 4137 10548 4168
rect 11790 4156 11796 4208
rect 11848 4196 11854 4208
rect 11848 4168 11928 4196
rect 11848 4156 11854 4168
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10870 4128 10876 4140
rect 10643 4100 10876 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10870 4088 10876 4100
rect 10928 4128 10934 4140
rect 11900 4137 11928 4168
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10928 4100 11069 4128
rect 10928 4088 10934 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12066 4088 12072 4140
rect 12124 4088 12130 4140
rect 12268 4128 12296 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 14642 4224 14648 4276
rect 14700 4224 14706 4276
rect 16850 4224 16856 4276
rect 16908 4224 16914 4276
rect 12437 4199 12495 4205
rect 12437 4165 12449 4199
rect 12483 4165 12495 4199
rect 12437 4159 12495 4165
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 12268 4100 12357 4128
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 8588 4032 8800 4060
rect 10778 4020 10784 4072
rect 10836 4020 10842 4072
rect 11238 4020 11244 4072
rect 11296 4020 11302 4072
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12452 4060 12480 4159
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13449 4199 13507 4205
rect 13449 4196 13461 4199
rect 13228 4168 13461 4196
rect 13228 4156 13234 4168
rect 13449 4165 13461 4168
rect 13495 4165 13507 4199
rect 13449 4159 13507 4165
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12676 4100 12909 4128
rect 12676 4088 12682 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 13357 4091 13415 4097
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14200 4128 14228 4224
rect 14568 4137 14596 4224
rect 14139 4100 14228 4128
rect 14553 4131 14611 4137
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14553 4097 14565 4131
rect 14599 4097 14611 4131
rect 14660 4128 14688 4224
rect 14918 4156 14924 4208
rect 14976 4156 14982 4208
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14660 4100 14749 4128
rect 14553 4091 14611 4097
rect 14737 4097 14749 4100
rect 14783 4097 14795 4131
rect 14936 4128 14964 4156
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 14936 4100 15485 4128
rect 14737 4091 14795 4097
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 15473 4091 15531 4097
rect 15764 4100 16773 4128
rect 13372 4060 13400 4091
rect 11848 4032 12480 4060
rect 12728 4032 13400 4060
rect 11848 4020 11854 4032
rect 5583 3964 5764 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6730 3952 6736 4004
rect 6788 3952 6794 4004
rect 2498 3924 2504 3936
rect 1504 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 6840 3924 6868 4020
rect 11256 3992 11284 4020
rect 12728 3992 12756 4032
rect 11256 3964 12756 3992
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13556 3992 13584 4091
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 15286 4060 15292 4072
rect 14691 4032 15292 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 15286 4020 15292 4032
rect 15344 4060 15350 4072
rect 15764 4069 15792 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16868 4128 16896 4224
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16868 4100 16957 4128
rect 16761 4091 16819 4097
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15344 4032 15761 4060
rect 15344 4020 15350 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16172 4032 16865 4060
rect 16172 4020 16178 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 12860 3964 13584 3992
rect 14185 3995 14243 4001
rect 12860 3952 12866 3964
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15562 3992 15568 4004
rect 14231 3964 15568 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 15562 3952 15568 3964
rect 15620 3952 15626 4004
rect 15657 3995 15715 4001
rect 15657 3961 15669 3995
rect 15703 3992 15715 3995
rect 17328 3992 17356 4020
rect 15703 3964 17356 3992
rect 15703 3961 15715 3964
rect 15657 3955 15715 3961
rect 5031 3896 6868 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7156 3896 7205 3924
rect 7156 3884 7162 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 10502 3924 10508 3936
rect 9824 3896 10508 3924
rect 9824 3884 9830 3896
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10686 3884 10692 3936
rect 10744 3884 10750 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12032 3896 13001 3924
rect 12032 3884 12038 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 1104 3834 18860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 18860 3834
rect 1104 3760 18860 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 1820 3692 2789 3720
rect 1820 3680 1826 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 3142 3680 3148 3732
rect 3200 3680 3206 3732
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4028 3692 6500 3720
rect 4028 3680 4034 3692
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 3160 3652 3188 3680
rect 1903 3624 3188 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3252 3584 3280 3680
rect 6472 3664 6500 3692
rect 6822 3680 6828 3732
rect 6880 3680 6886 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8168 3692 8493 3720
rect 8168 3680 8174 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 9306 3680 9312 3732
rect 9364 3680 9370 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 10134 3720 10140 3732
rect 9723 3692 10140 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11204 3692 11468 3720
rect 11204 3680 11210 3692
rect 6362 3652 6368 3664
rect 2915 3556 3280 3584
rect 3344 3624 6368 3652
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 992 3488 1777 3516
rect 992 3476 998 3488
rect 1765 3485 1777 3488
rect 1811 3516 1823 3519
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1811 3488 2237 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2590 3476 2596 3528
rect 2648 3476 2654 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2774 3516 2780 3528
rect 2731 3488 2780 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3344 3516 3372 3624
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 6454 3612 6460 3664
rect 6512 3612 6518 3664
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5813 3587 5871 3593
rect 5408 3556 5580 3584
rect 5408 3544 5414 3556
rect 3292 3488 3372 3516
rect 4157 3519 4215 3525
rect 3292 3476 3298 3488
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4798 3516 4804 3528
rect 4387 3488 4804 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 3326 3448 3332 3460
rect 2464 3420 3332 3448
rect 2464 3408 2470 3420
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 4172 3448 4200 3479
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 4614 3448 4620 3460
rect 4172 3420 4620 3448
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 5552 3392 5580 3556
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 6840 3584 6868 3680
rect 5859 3556 6868 3584
rect 7009 3587 7067 3593
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7098 3584 7104 3596
rect 7055 3556 7104 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5736 3448 5764 3479
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6696 3488 6745 3516
rect 6696 3476 6702 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 8754 3516 8760 3528
rect 8142 3488 8760 3516
rect 6733 3479 6791 3485
rect 8754 3476 8760 3488
rect 8812 3516 8818 3528
rect 9324 3516 9352 3680
rect 11440 3652 11468 3692
rect 11790 3680 11796 3732
rect 11848 3720 11854 3732
rect 12802 3720 12808 3732
rect 11848 3692 12808 3720
rect 11848 3680 11854 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13078 3680 13084 3732
rect 13136 3680 13142 3732
rect 15562 3680 15568 3732
rect 15620 3680 15626 3732
rect 15654 3680 15660 3732
rect 15712 3680 15718 3732
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 15988 3692 16405 3720
rect 15988 3680 15994 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 16945 3723 17003 3729
rect 16945 3689 16957 3723
rect 16991 3720 17003 3723
rect 17862 3720 17868 3732
rect 16991 3692 17868 3720
rect 16991 3689 17003 3692
rect 16945 3683 17003 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 12618 3652 12624 3664
rect 11440 3624 12624 3652
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11440 3593 11468 3624
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10744 3556 11161 3584
rect 10744 3544 10750 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 11425 3587 11483 3593
rect 11425 3553 11437 3587
rect 11471 3553 11483 3587
rect 12710 3584 12716 3596
rect 11425 3547 11483 3553
rect 12406 3556 12716 3584
rect 8812 3502 10074 3516
rect 8812 3488 10088 3502
rect 8812 3476 8818 3488
rect 5736 3420 6776 3448
rect 6748 3392 6776 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3510 3380 3516 3392
rect 2924 3352 3516 3380
rect 2924 3340 2930 3352
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 4341 3383 4399 3389
rect 4341 3349 4353 3383
rect 4387 3380 4399 3383
rect 4890 3380 4896 3392
rect 4387 3352 4896 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5534 3340 5540 3392
rect 5592 3340 5598 3392
rect 6730 3340 6736 3392
rect 6788 3340 6794 3392
rect 10060 3380 10088 3488
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11572 3488 11713 3516
rect 11572 3476 11578 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11885 3519 11943 3525
rect 11885 3485 11897 3519
rect 11931 3516 11943 3519
rect 12406 3516 12434 3556
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 13096 3584 13124 3680
rect 12912 3556 13124 3584
rect 13173 3587 13231 3593
rect 12912 3525 12940 3556
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 13219 3556 14473 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 14461 3547 14519 3553
rect 14568 3556 15393 3584
rect 11931 3488 12434 3516
rect 12621 3519 12679 3525
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13035 3488 13737 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 13998 3516 14004 3528
rect 13863 3488 14004 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 12345 3451 12403 3457
rect 12345 3448 12357 3451
rect 12124 3420 12357 3448
rect 12124 3408 12130 3420
rect 12345 3417 12357 3420
rect 12391 3417 12403 3451
rect 12345 3411 12403 3417
rect 10962 3380 10968 3392
rect 10060 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 12636 3380 12664 3479
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14366 3476 14372 3528
rect 14424 3476 14430 3528
rect 14568 3525 14596 3556
rect 15381 3553 15393 3556
rect 15427 3553 15439 3587
rect 15580 3584 15608 3680
rect 15672 3652 15700 3680
rect 15672 3624 16620 3652
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15580 3556 15669 3584
rect 15381 3547 15439 3553
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14918 3476 14924 3528
rect 14976 3476 14982 3528
rect 15746 3476 15752 3528
rect 15804 3476 15810 3528
rect 16592 3525 16620 3624
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16623 3488 16865 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 14936 3448 14964 3476
rect 16408 3448 16436 3479
rect 13096 3420 13308 3448
rect 14936 3420 16436 3448
rect 13096 3380 13124 3420
rect 11296 3352 13124 3380
rect 11296 3340 11302 3352
rect 13170 3340 13176 3392
rect 13228 3340 13234 3392
rect 13280 3380 13308 3420
rect 17586 3380 17592 3392
rect 13280 3352 17592 3380
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 1104 3290 18860 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 18860 3290
rect 1104 3216 18860 3238
rect 5077 3179 5135 3185
rect 3436 3148 4936 3176
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 3436 3049 3464 3148
rect 4908 3108 4936 3148
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5442 3176 5448 3188
rect 5123 3148 5448 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 6420 3148 7236 3176
rect 6420 3136 6426 3148
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 3804 3080 4844 3108
rect 4908 3080 6561 3108
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 1854 2932 1860 2984
rect 1912 2972 1918 2984
rect 1949 2975 2007 2981
rect 1949 2972 1961 2975
rect 1912 2944 1961 2972
rect 1912 2932 1918 2944
rect 1949 2941 1961 2944
rect 1995 2941 2007 2975
rect 3252 2972 3280 3003
rect 3326 2972 3332 2984
rect 3252 2944 3332 2972
rect 1949 2935 2007 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3804 2972 3832 3080
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 3970 3040 3976 3052
rect 3927 3012 3976 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4816 3049 4844 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 3436 2944 3832 2972
rect 3436 2913 3464 2944
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2873 3479 2907
rect 4080 2904 4108 3003
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 4908 2972 4936 3000
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4908 2944 5089 2972
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 4614 2904 4620 2916
rect 4080 2876 4620 2904
rect 3421 2867 3479 2873
rect 4614 2864 4620 2876
rect 4672 2904 4678 2916
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 4672 2876 4905 2904
rect 4672 2864 4678 2876
rect 4893 2873 4905 2876
rect 4939 2873 4951 2907
rect 5368 2904 5396 3003
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 7208 3049 7236 3148
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7800 3148 7849 3176
rect 7800 3136 7806 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8168 3148 8524 3176
rect 8168 3136 8174 3148
rect 7466 3108 7472 3120
rect 7392 3080 7472 3108
rect 7392 3049 7420 3080
rect 7466 3068 7472 3080
rect 7524 3108 7530 3120
rect 8496 3117 8524 3148
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 10778 3176 10784 3188
rect 10183 3148 10784 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11020 3148 11621 3176
rect 11020 3136 11026 3148
rect 11609 3145 11621 3148
rect 11655 3176 11667 3179
rect 11790 3176 11796 3188
rect 11655 3148 11796 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 13170 3176 13176 3188
rect 12912 3148 13176 3176
rect 8481 3111 8539 3117
rect 7524 3080 8432 3108
rect 7524 3068 7530 3080
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7926 3040 7932 3052
rect 7377 3003 7435 3009
rect 7852 3012 7932 3040
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 6270 2972 6276 2984
rect 5491 2944 6276 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 4893 2867 4951 2873
rect 5000 2876 5396 2904
rect 2406 2796 2412 2848
rect 2464 2796 2470 2848
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 5000 2836 5028 2876
rect 4111 2808 5028 2836
rect 7208 2836 7236 3003
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7852 2972 7880 3012
rect 7926 3000 7932 3012
rect 7984 3040 7990 3052
rect 8404 3049 8432 3080
rect 8481 3077 8493 3111
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 9306 3108 9312 3120
rect 8628 3080 9312 3108
rect 8628 3068 8634 3080
rect 9306 3068 9312 3080
rect 9364 3108 9370 3120
rect 9364 3080 9444 3108
rect 9364 3068 9370 3080
rect 9416 3049 9444 3080
rect 10042 3068 10048 3120
rect 10100 3068 10106 3120
rect 10888 3108 10916 3136
rect 12912 3117 12940 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 14918 3136 14924 3188
rect 14976 3136 14982 3188
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 15746 3176 15752 3188
rect 15519 3148 15752 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 10152 3080 10916 3108
rect 12897 3111 12955 3117
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7984 3012 8125 3040
rect 7984 3000 7990 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 9401 3043 9459 3049
rect 8435 3012 9168 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 9140 2981 9168 3012
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10060 3040 10088 3068
rect 10152 3049 10180 3080
rect 12897 3077 12909 3111
rect 12943 3077 12955 3111
rect 12897 3071 12955 3077
rect 13906 3068 13912 3120
rect 13964 3068 13970 3120
rect 14550 3068 14556 3120
rect 14608 3108 14614 3120
rect 14645 3111 14703 3117
rect 14645 3108 14657 3111
rect 14608 3080 14657 3108
rect 14608 3068 14614 3080
rect 14645 3077 14657 3080
rect 14691 3077 14703 3111
rect 14936 3108 14964 3136
rect 14936 3080 15976 3108
rect 14645 3071 14703 3077
rect 9999 3012 10088 3040
rect 10137 3043 10195 3049
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 10594 3000 10600 3052
rect 10652 3000 10658 3052
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 10744 3012 10793 3040
rect 10744 3000 10750 3012
rect 10781 3009 10793 3012
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 7331 2944 7880 2972
rect 8021 2975 8079 2981
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 8021 2941 8033 2975
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 10336 2972 10364 3000
rect 10888 2972 10916 3003
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11756 3012 11989 3040
rect 11756 3000 11762 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 10336 2944 10916 2972
rect 9125 2935 9183 2941
rect 8036 2904 8064 2935
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 12066 2972 12072 2984
rect 11112 2944 12072 2972
rect 11112 2932 11118 2944
rect 12066 2932 12072 2944
rect 12124 2972 12130 2984
rect 12176 2972 12204 3003
rect 15286 3000 15292 3052
rect 15344 3000 15350 3052
rect 15948 3049 15976 3080
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3040 15531 3043
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 15519 3012 15853 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 12124 2944 12204 2972
rect 12124 2932 12130 2944
rect 12618 2932 12624 2984
rect 12676 2932 12682 2984
rect 9030 2904 9036 2916
rect 8036 2876 9036 2904
rect 9030 2864 9036 2876
rect 9088 2904 9094 2916
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 9088 2876 9321 2904
rect 9088 2864 9094 2876
rect 9309 2873 9321 2876
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 10686 2864 10692 2916
rect 10744 2904 10750 2916
rect 11238 2904 11244 2916
rect 10744 2876 11244 2904
rect 10744 2864 10750 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 8570 2836 8576 2848
rect 7208 2808 8576 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 9214 2796 9220 2848
rect 9272 2796 9278 2848
rect 12066 2796 12072 2848
rect 12124 2796 12130 2848
rect 1104 2746 18860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 18860 2746
rect 1104 2672 18860 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3878 2632 3884 2644
rect 2915 2604 3884 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4614 2632 4620 2644
rect 4571 2604 4620 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 6730 2592 6736 2644
rect 6788 2632 6794 2644
rect 6825 2635 6883 2641
rect 6825 2632 6837 2635
rect 6788 2604 6837 2632
rect 6788 2592 6794 2604
rect 6825 2601 6837 2604
rect 6871 2601 6883 2635
rect 6825 2595 6883 2601
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7064 2604 8984 2632
rect 7064 2592 7070 2604
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 4706 2564 4712 2576
rect 2179 2536 4712 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 2501 2499 2559 2505
rect 2501 2496 2513 2499
rect 2464 2468 2513 2496
rect 2464 2456 2470 2468
rect 2501 2465 2513 2468
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 3418 2456 3424 2508
rect 3476 2456 3482 2508
rect 1854 2388 1860 2440
rect 1912 2388 1918 2440
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2038 2428 2044 2440
rect 1995 2400 2044 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2038 2388 2044 2400
rect 2096 2428 2102 2440
rect 2593 2431 2651 2437
rect 2096 2400 2360 2428
rect 2096 2388 2102 2400
rect 2332 2304 2360 2400
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 3326 2428 3332 2440
rect 2639 2400 3332 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 4264 2437 4292 2536
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 5868 2536 6914 2564
rect 5868 2524 5874 2536
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4356 2360 4384 2459
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5500 2468 5750 2496
rect 5500 2456 5506 2468
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 6886 2428 6914 2536
rect 7926 2524 7932 2576
rect 7984 2524 7990 2576
rect 8956 2564 8984 2604
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 9088 2604 9137 2632
rect 9088 2592 9094 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 10597 2635 10655 2641
rect 10597 2601 10609 2635
rect 10643 2632 10655 2635
rect 10962 2632 10968 2644
rect 10643 2604 10968 2632
rect 10643 2601 10655 2604
rect 10597 2595 10655 2601
rect 8956 2536 9720 2564
rect 7944 2496 7972 2524
rect 8297 2499 8355 2505
rect 7944 2468 8064 2496
rect 8036 2437 8064 2468
rect 8297 2465 8309 2499
rect 8343 2496 8355 2499
rect 9214 2496 9220 2508
rect 8343 2468 9220 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9692 2440 9720 2536
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 6886 2400 7941 2428
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8662 2428 8668 2440
rect 8021 2391 8079 2397
rect 8128 2400 8668 2428
rect 4798 2360 4804 2372
rect 4356 2332 4804 2360
rect 4798 2320 4804 2332
rect 4856 2360 4862 2372
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 4856 2332 5457 2360
rect 4856 2320 4862 2332
rect 5445 2329 5457 2332
rect 5491 2329 5503 2363
rect 7944 2360 7972 2391
rect 8128 2360 8156 2400
rect 8662 2388 8668 2400
rect 8720 2428 8726 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8720 2400 9045 2428
rect 8720 2388 8726 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9674 2388 9680 2440
rect 9732 2388 9738 2440
rect 10137 2431 10195 2437
rect 10137 2397 10149 2431
rect 10183 2428 10195 2431
rect 10612 2428 10640 2595
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 12066 2592 12072 2644
rect 12124 2592 12130 2644
rect 11790 2524 11796 2576
rect 11848 2524 11854 2576
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12084 2496 12112 2592
rect 11471 2468 12112 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 13446 2496 13452 2508
rect 12860 2468 13452 2496
rect 12860 2456 12866 2468
rect 13446 2456 13452 2468
rect 13504 2496 13510 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13504 2468 13829 2496
rect 13504 2456 13510 2468
rect 13817 2465 13829 2468
rect 13863 2496 13875 2499
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13863 2468 14197 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 10183 2400 10640 2428
rect 10183 2397 10195 2400
rect 10137 2391 10195 2397
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11698 2428 11704 2440
rect 11256 2400 11704 2428
rect 7944 2332 8156 2360
rect 8389 2363 8447 2369
rect 5445 2323 5503 2329
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 9585 2363 9643 2369
rect 9585 2360 9597 2363
rect 8435 2332 9597 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 9585 2329 9597 2332
rect 9631 2360 9643 2363
rect 10226 2360 10232 2372
rect 9631 2332 10232 2360
rect 9631 2329 9643 2332
rect 9585 2323 9643 2329
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 10468 2332 10793 2360
rect 10468 2320 10474 2332
rect 10781 2329 10793 2332
rect 10827 2360 10839 2363
rect 11256 2360 11284 2400
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 10827 2332 11284 2360
rect 11425 2363 11483 2369
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11425 2329 11437 2363
rect 11471 2360 11483 2363
rect 11471 2332 12296 2360
rect 11471 2329 11483 2332
rect 11425 2323 11483 2329
rect 2314 2252 2320 2304
rect 2372 2252 2378 2304
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2292 7251 2295
rect 7650 2292 7656 2304
rect 7239 2264 7656 2292
rect 7239 2261 7251 2264
rect 7193 2255 7251 2261
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 10042 2252 10048 2304
rect 10100 2252 10106 2304
rect 10581 2295 10639 2301
rect 10581 2261 10593 2295
rect 10627 2292 10639 2295
rect 11974 2292 11980 2304
rect 10627 2264 11980 2292
rect 10627 2261 10639 2264
rect 10581 2255 10639 2261
rect 11974 2252 11980 2264
rect 12032 2292 12038 2304
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 12032 2264 12081 2292
rect 12032 2252 12038 2264
rect 12069 2261 12081 2264
rect 12115 2261 12127 2295
rect 12268 2292 12296 2332
rect 12894 2320 12900 2372
rect 12952 2320 12958 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 13556 2292 13584 2323
rect 14090 2320 14096 2372
rect 14148 2320 14154 2372
rect 14458 2320 14464 2372
rect 14516 2320 14522 2372
rect 14568 2332 14950 2360
rect 12268 2264 13584 2292
rect 14108 2292 14136 2320
rect 14568 2292 14596 2332
rect 14108 2264 14596 2292
rect 15933 2295 15991 2301
rect 12069 2255 12127 2261
rect 15933 2261 15945 2295
rect 15979 2292 15991 2295
rect 16942 2292 16948 2304
rect 15979 2264 16948 2292
rect 15979 2261 15991 2264
rect 15933 2255 15991 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 1104 2202 18860 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 18860 2202
rect 1104 2128 18860 2150
rect 1673 2091 1731 2097
rect 1673 2057 1685 2091
rect 1719 2088 1731 2091
rect 1854 2088 1860 2100
rect 1719 2060 1860 2088
rect 1719 2057 1731 2060
rect 1673 2051 1731 2057
rect 1854 2048 1860 2060
rect 1912 2088 1918 2100
rect 1912 2060 3740 2088
rect 1912 2048 1918 2060
rect 3418 2020 3424 2032
rect 2714 1992 3424 2020
rect 3418 1980 3424 1992
rect 3476 2020 3482 2032
rect 3476 1992 3648 2020
rect 3476 1980 3482 1992
rect 3142 1844 3148 1896
rect 3200 1844 3206 1896
rect 3421 1887 3479 1893
rect 3421 1884 3433 1887
rect 3344 1856 3433 1884
rect 3344 1816 3372 1856
rect 3421 1853 3433 1856
rect 3467 1853 3479 1887
rect 3620 1884 3648 1992
rect 3712 1961 3740 2060
rect 7006 2048 7012 2100
rect 7064 2048 7070 2100
rect 7926 2088 7932 2100
rect 7576 2060 7932 2088
rect 5813 2023 5871 2029
rect 5813 1989 5825 2023
rect 5859 2020 5871 2023
rect 6733 2023 6791 2029
rect 6733 2020 6745 2023
rect 5859 1992 6745 2020
rect 5859 1989 5871 1992
rect 5813 1983 5871 1989
rect 6733 1989 6745 1992
rect 6779 1989 6791 2023
rect 7024 2020 7052 2048
rect 7576 2029 7604 2060
rect 7926 2048 7932 2060
rect 7984 2048 7990 2100
rect 9674 2048 9680 2100
rect 9732 2048 9738 2100
rect 10042 2048 10048 2100
rect 10100 2048 10106 2100
rect 10226 2048 10232 2100
rect 10284 2088 10290 2100
rect 10284 2060 10732 2088
rect 10284 2048 10290 2060
rect 6733 1983 6791 1989
rect 6932 1992 7052 2020
rect 7561 2023 7619 2029
rect 6932 1964 6960 1992
rect 7561 1989 7573 2023
rect 7607 1989 7619 2023
rect 7561 1983 7619 1989
rect 9306 1980 9312 2032
rect 9364 1980 9370 2032
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 3988 1924 4738 1952
rect 3988 1884 4016 1924
rect 6914 1912 6920 1964
rect 6972 1912 6978 1964
rect 7006 1912 7012 1964
rect 7064 1912 7070 1964
rect 8694 1924 8800 1952
rect 3620 1856 4016 1884
rect 4341 1887 4399 1893
rect 3421 1847 3479 1853
rect 4341 1853 4353 1887
rect 4387 1884 4399 1887
rect 5442 1884 5448 1896
rect 4387 1856 5448 1884
rect 4387 1853 4399 1856
rect 4341 1847 4399 1853
rect 5442 1844 5448 1856
rect 5500 1844 5506 1896
rect 6089 1887 6147 1893
rect 6089 1853 6101 1887
rect 6135 1853 6147 1887
rect 6089 1847 6147 1853
rect 6104 1816 6132 1847
rect 6362 1844 6368 1896
rect 6420 1884 6426 1896
rect 6733 1887 6791 1893
rect 6733 1884 6745 1887
rect 6420 1856 6745 1884
rect 6420 1844 6426 1856
rect 6733 1853 6745 1856
rect 6779 1853 6791 1887
rect 7285 1887 7343 1893
rect 7285 1884 7297 1887
rect 6733 1847 6791 1853
rect 6886 1856 7297 1884
rect 6638 1816 6644 1828
rect 3344 1788 4844 1816
rect 3344 1760 3372 1788
rect 2774 1708 2780 1760
rect 2832 1748 2838 1760
rect 3326 1748 3332 1760
rect 2832 1720 3332 1748
rect 2832 1708 2838 1720
rect 3326 1708 3332 1720
rect 3384 1708 3390 1760
rect 3786 1708 3792 1760
rect 3844 1708 3850 1760
rect 4816 1748 4844 1788
rect 6104 1788 6644 1816
rect 6104 1748 6132 1788
rect 6638 1776 6644 1788
rect 6696 1816 6702 1828
rect 6886 1816 6914 1856
rect 7285 1853 7297 1856
rect 7331 1884 7343 1887
rect 8018 1884 8024 1896
rect 7331 1856 8024 1884
rect 7331 1853 7343 1856
rect 7285 1847 7343 1853
rect 8018 1844 8024 1856
rect 8076 1844 8082 1896
rect 8772 1828 8800 1924
rect 9692 1884 9720 2048
rect 10060 1961 10088 2048
rect 10244 1961 10272 2048
rect 10410 1980 10416 2032
rect 10468 1980 10474 2032
rect 10704 2029 10732 2060
rect 11698 2048 11704 2100
rect 11756 2048 11762 2100
rect 11790 2048 11796 2100
rect 11848 2088 11854 2100
rect 13725 2091 13783 2097
rect 11848 2060 12848 2088
rect 11848 2048 11854 2060
rect 10689 2023 10747 2029
rect 10689 1989 10701 2023
rect 10735 1989 10747 2023
rect 11054 2020 11060 2032
rect 10689 1983 10747 1989
rect 10796 1992 11060 2020
rect 10045 1955 10103 1961
rect 10045 1921 10057 1955
rect 10091 1921 10103 1955
rect 10045 1915 10103 1921
rect 10229 1955 10287 1961
rect 10229 1921 10241 1955
rect 10275 1921 10287 1955
rect 10428 1952 10456 1980
rect 10796 1961 10824 1992
rect 11054 1980 11060 1992
rect 11112 1980 11118 2032
rect 12820 2020 12848 2060
rect 13725 2057 13737 2091
rect 13771 2088 13783 2091
rect 14458 2088 14464 2100
rect 13771 2060 14464 2088
rect 13771 2057 13783 2060
rect 13725 2051 13783 2057
rect 14458 2048 14464 2060
rect 14516 2048 14522 2100
rect 12894 2020 12900 2032
rect 12742 1992 12900 2020
rect 12894 1980 12900 1992
rect 12952 2020 12958 2032
rect 13906 2020 13912 2032
rect 12952 1992 13912 2020
rect 12952 1980 12958 1992
rect 13906 1980 13912 1992
rect 13964 1980 13970 2032
rect 14918 1980 14924 2032
rect 14976 2020 14982 2032
rect 15197 2023 15255 2029
rect 15197 2020 15209 2023
rect 14976 1992 15209 2020
rect 14976 1980 14982 1992
rect 15197 1989 15209 1992
rect 15243 2020 15255 2023
rect 15749 2023 15807 2029
rect 15749 2020 15761 2023
rect 15243 1992 15761 2020
rect 15243 1989 15255 1992
rect 15197 1983 15255 1989
rect 15749 1989 15761 1992
rect 15795 1989 15807 2023
rect 15749 1983 15807 1989
rect 17586 1980 17592 2032
rect 17644 1980 17650 2032
rect 16948 1964 17000 1970
rect 10505 1955 10563 1961
rect 10505 1952 10517 1955
rect 10428 1924 10517 1952
rect 10229 1915 10287 1921
rect 10505 1921 10517 1924
rect 10551 1921 10563 1955
rect 10505 1915 10563 1921
rect 10781 1955 10839 1961
rect 10781 1921 10793 1955
rect 10827 1921 10839 1955
rect 10781 1915 10839 1921
rect 10873 1955 10931 1961
rect 10873 1921 10885 1955
rect 10919 1952 10931 1955
rect 10962 1952 10968 1964
rect 10919 1924 10968 1952
rect 10919 1921 10931 1924
rect 10873 1915 10931 1921
rect 10796 1884 10824 1915
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 13446 1912 13452 1964
rect 13504 1912 13510 1964
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 14090 1952 14096 1964
rect 13596 1924 14096 1952
rect 13596 1912 13602 1924
rect 14090 1912 14096 1924
rect 14148 1912 14154 1964
rect 16114 1912 16120 1964
rect 16172 1952 16178 1964
rect 16853 1955 16911 1961
rect 16853 1952 16865 1955
rect 16172 1924 16865 1952
rect 16172 1912 16178 1924
rect 16853 1921 16865 1924
rect 16899 1921 16911 1955
rect 16853 1915 16911 1921
rect 13173 1887 13231 1893
rect 13173 1884 13185 1887
rect 9692 1856 10824 1884
rect 11072 1856 13185 1884
rect 6696 1788 6914 1816
rect 6696 1776 6702 1788
rect 8754 1776 8760 1828
rect 8812 1816 8818 1828
rect 9674 1816 9680 1828
rect 8812 1788 9680 1816
rect 8812 1776 8818 1788
rect 9674 1776 9680 1788
rect 9732 1816 9738 1828
rect 11072 1825 11100 1856
rect 13173 1853 13185 1856
rect 13219 1853 13231 1887
rect 13464 1884 13492 1912
rect 16948 1906 17000 1912
rect 15473 1887 15531 1893
rect 15473 1884 15485 1887
rect 13464 1856 15485 1884
rect 13173 1847 13231 1853
rect 15473 1853 15485 1856
rect 15519 1853 15531 1887
rect 15473 1847 15531 1853
rect 11057 1819 11115 1825
rect 9732 1788 10272 1816
rect 9732 1776 9738 1788
rect 4816 1720 6132 1748
rect 10134 1708 10140 1760
rect 10192 1708 10198 1760
rect 10244 1748 10272 1788
rect 11057 1785 11069 1819
rect 11103 1785 11115 1819
rect 11057 1779 11115 1785
rect 11790 1776 11796 1828
rect 11848 1776 11854 1828
rect 11808 1748 11836 1776
rect 10244 1720 11836 1748
rect 1104 1658 18860 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 18860 1658
rect 1104 1584 18860 1606
rect 2314 1504 2320 1556
rect 2372 1504 2378 1556
rect 3234 1504 3240 1556
rect 3292 1504 3298 1556
rect 5997 1547 6055 1553
rect 5997 1513 6009 1547
rect 6043 1544 6055 1547
rect 6362 1544 6368 1556
rect 6043 1516 6368 1544
rect 6043 1513 6055 1516
rect 5997 1507 6055 1513
rect 6362 1504 6368 1516
rect 6420 1504 6426 1556
rect 7006 1544 7012 1556
rect 6886 1516 7012 1544
rect 3252 1476 3280 1504
rect 3160 1448 3280 1476
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 2409 1343 2467 1349
rect 2409 1309 2421 1343
rect 2455 1340 2467 1343
rect 2685 1343 2743 1349
rect 2685 1340 2697 1343
rect 2455 1312 2697 1340
rect 2455 1309 2467 1312
rect 2409 1303 2467 1309
rect 2685 1309 2697 1312
rect 2731 1340 2743 1343
rect 2866 1340 2872 1352
rect 2731 1312 2872 1340
rect 2731 1309 2743 1312
rect 2685 1303 2743 1309
rect 1780 1272 1808 1303
rect 2866 1300 2872 1312
rect 2924 1300 2930 1352
rect 3050 1300 3056 1352
rect 3108 1300 3114 1352
rect 3160 1349 3188 1448
rect 3510 1436 3516 1488
rect 3568 1476 3574 1488
rect 4341 1479 4399 1485
rect 4341 1476 4353 1479
rect 3568 1448 4353 1476
rect 3568 1436 3574 1448
rect 4341 1445 4353 1448
rect 4387 1476 4399 1479
rect 5353 1479 5411 1485
rect 4387 1448 4844 1476
rect 4387 1445 4399 1448
rect 4341 1439 4399 1445
rect 3237 1416 3295 1417
rect 3237 1411 3464 1416
rect 3237 1377 3249 1411
rect 3283 1408 3464 1411
rect 4157 1411 4215 1417
rect 4157 1408 4169 1411
rect 3283 1388 4169 1408
rect 3283 1377 3295 1388
rect 3436 1380 4169 1388
rect 3237 1371 3295 1377
rect 4157 1377 4169 1380
rect 4203 1377 4215 1411
rect 4157 1371 4215 1377
rect 4356 1380 4568 1408
rect 3145 1343 3203 1349
rect 3145 1309 3157 1343
rect 3191 1309 3203 1343
rect 3145 1303 3203 1309
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1340 3387 1343
rect 3418 1340 3424 1352
rect 3375 1312 3424 1340
rect 3375 1309 3387 1312
rect 3329 1303 3387 1309
rect 3418 1300 3424 1312
rect 3476 1300 3482 1352
rect 4356 1340 4384 1380
rect 3528 1312 4384 1340
rect 4433 1343 4491 1349
rect 3068 1272 3096 1300
rect 3528 1272 3556 1312
rect 4433 1309 4445 1343
rect 4479 1309 4491 1343
rect 4540 1340 4568 1380
rect 4709 1343 4767 1349
rect 4709 1340 4721 1343
rect 4540 1312 4721 1340
rect 4433 1303 4491 1309
rect 4709 1309 4721 1312
rect 4755 1309 4767 1343
rect 4709 1303 4767 1309
rect 1780 1244 3556 1272
rect 3786 1232 3792 1284
rect 3844 1272 3850 1284
rect 4448 1272 4476 1303
rect 3844 1244 4476 1272
rect 4816 1272 4844 1448
rect 5353 1445 5365 1479
rect 5399 1476 5411 1479
rect 6886 1476 6914 1516
rect 7006 1504 7012 1516
rect 7064 1504 7070 1556
rect 7742 1504 7748 1556
rect 7800 1544 7806 1556
rect 8125 1547 8183 1553
rect 8125 1544 8137 1547
rect 7800 1516 8137 1544
rect 7800 1504 7806 1516
rect 8125 1513 8137 1516
rect 8171 1513 8183 1547
rect 8125 1507 8183 1513
rect 9125 1547 9183 1553
rect 9125 1513 9137 1547
rect 9171 1544 9183 1547
rect 9674 1544 9680 1556
rect 9171 1516 9680 1544
rect 9171 1513 9183 1516
rect 9125 1507 9183 1513
rect 9674 1504 9680 1516
rect 9732 1504 9738 1556
rect 11146 1504 11152 1556
rect 11204 1544 11210 1556
rect 12253 1547 12311 1553
rect 12253 1544 12265 1547
rect 11204 1516 12265 1544
rect 11204 1504 11210 1516
rect 12253 1513 12265 1516
rect 12299 1513 12311 1547
rect 12253 1507 12311 1513
rect 14632 1547 14690 1553
rect 14632 1513 14644 1547
rect 14678 1544 14690 1547
rect 14678 1516 16068 1544
rect 14678 1513 14690 1516
rect 14632 1507 14690 1513
rect 5399 1448 6914 1476
rect 11701 1479 11759 1485
rect 5399 1445 5411 1448
rect 5353 1439 5411 1445
rect 11701 1445 11713 1479
rect 11747 1476 11759 1479
rect 11790 1476 11796 1488
rect 11747 1448 11796 1476
rect 11747 1445 11759 1448
rect 11701 1439 11759 1445
rect 11790 1436 11796 1448
rect 11848 1436 11854 1488
rect 11974 1436 11980 1488
rect 12032 1436 12038 1488
rect 16040 1476 16068 1516
rect 16114 1504 16120 1556
rect 16172 1504 16178 1556
rect 16942 1544 16948 1556
rect 16546 1516 16948 1544
rect 16546 1476 16574 1516
rect 16942 1504 16948 1516
rect 17000 1504 17006 1556
rect 16040 1448 16574 1476
rect 5442 1368 5448 1420
rect 5500 1368 5506 1420
rect 5810 1368 5816 1420
rect 5868 1408 5874 1420
rect 6641 1411 6699 1417
rect 6641 1408 6653 1411
rect 5868 1380 6653 1408
rect 5868 1368 5874 1380
rect 5261 1343 5319 1349
rect 5261 1309 5273 1343
rect 5307 1340 5319 1343
rect 5460 1340 5488 1368
rect 6104 1349 6132 1380
rect 6641 1377 6653 1380
rect 6687 1377 6699 1411
rect 6914 1408 6920 1420
rect 6641 1371 6699 1377
rect 6886 1368 6920 1408
rect 6972 1368 6978 1420
rect 8018 1368 8024 1420
rect 8076 1408 8082 1420
rect 9677 1411 9735 1417
rect 8076 1380 8432 1408
rect 8076 1368 8082 1380
rect 5307 1312 5488 1340
rect 5905 1343 5963 1349
rect 5307 1309 5319 1312
rect 5261 1303 5319 1309
rect 5905 1309 5917 1343
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1309 6147 1343
rect 6886 1340 6914 1368
rect 8404 1349 8432 1380
rect 9677 1377 9689 1411
rect 9723 1408 9735 1411
rect 10134 1408 10140 1420
rect 9723 1380 10140 1408
rect 9723 1377 9735 1380
rect 9677 1371 9735 1377
rect 10134 1368 10140 1380
rect 10192 1368 10198 1420
rect 6089 1303 6147 1309
rect 6196 1312 6914 1340
rect 8389 1343 8447 1349
rect 5920 1272 5948 1303
rect 6196 1272 6224 1312
rect 8389 1309 8401 1343
rect 8435 1340 8447 1343
rect 9401 1343 9459 1349
rect 9401 1340 9413 1343
rect 8435 1312 9413 1340
rect 8435 1309 8447 1312
rect 8389 1303 8447 1309
rect 9401 1309 9413 1312
rect 9447 1309 9459 1343
rect 11992 1340 12020 1436
rect 13446 1368 13452 1420
rect 13504 1408 13510 1420
rect 14369 1411 14427 1417
rect 14369 1408 14381 1411
rect 13504 1380 14381 1408
rect 13504 1368 13510 1380
rect 14369 1377 14381 1380
rect 14415 1377 14427 1411
rect 14369 1371 14427 1377
rect 12161 1343 12219 1349
rect 12161 1340 12173 1343
rect 11992 1312 12173 1340
rect 9401 1303 9459 1309
rect 12161 1309 12173 1312
rect 12207 1309 12219 1343
rect 12161 1303 12219 1309
rect 4816 1244 6224 1272
rect 3844 1232 3850 1244
rect 7650 1232 7656 1284
rect 7708 1272 7714 1284
rect 8754 1272 8760 1284
rect 7708 1244 8760 1272
rect 7708 1232 7714 1244
rect 8754 1232 8760 1244
rect 8812 1232 8818 1284
rect 13538 1272 13544 1284
rect 10902 1244 13544 1272
rect 13538 1232 13544 1244
rect 13596 1232 13602 1284
rect 13817 1275 13875 1281
rect 13817 1241 13829 1275
rect 13863 1272 13875 1275
rect 13906 1272 13912 1284
rect 13863 1244 13912 1272
rect 13863 1241 13875 1244
rect 13817 1235 13875 1241
rect 13906 1232 13912 1244
rect 13964 1272 13970 1284
rect 13964 1244 15134 1272
rect 13964 1232 13970 1244
rect 1854 1164 1860 1216
rect 1912 1164 1918 1216
rect 3142 1164 3148 1216
rect 3200 1204 3206 1216
rect 4157 1207 4215 1213
rect 4157 1204 4169 1207
rect 3200 1176 4169 1204
rect 3200 1164 3206 1176
rect 4157 1173 4169 1176
rect 4203 1173 4215 1207
rect 4157 1167 4215 1173
rect 10962 1164 10968 1216
rect 11020 1204 11026 1216
rect 11149 1207 11207 1213
rect 11149 1204 11161 1207
rect 11020 1176 11161 1204
rect 11020 1164 11026 1176
rect 11149 1173 11161 1176
rect 11195 1173 11207 1207
rect 11149 1167 11207 1173
rect 1104 1114 18860 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 18860 1114
rect 1104 1040 18860 1062
rect 1854 960 1860 1012
rect 1912 1000 1918 1012
rect 5626 1000 5632 1012
rect 1912 972 5632 1000
rect 1912 960 1918 972
rect 5626 960 5632 972
rect 5684 960 5690 1012
<< via1 >>
rect 15016 13880 15068 13932
rect 15844 13880 15896 13932
rect 7196 13744 7248 13796
rect 15200 13744 15252 13796
rect 1124 13676 1176 13728
rect 4804 13676 4856 13728
rect 11244 13676 11296 13728
rect 17408 13676 17460 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 10048 13472 10100 13524
rect 7012 13404 7064 13456
rect 11244 13404 11296 13456
rect 1032 13336 1084 13388
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 3884 13336 3936 13388
rect 5080 13268 5132 13320
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 2504 13175 2556 13184
rect 2504 13141 2513 13175
rect 2513 13141 2547 13175
rect 2547 13141 2556 13175
rect 2504 13132 2556 13141
rect 3240 13132 3292 13184
rect 3976 13243 4028 13252
rect 3976 13209 3985 13243
rect 3985 13209 4019 13243
rect 4019 13209 4028 13243
rect 3976 13200 4028 13209
rect 10600 13336 10652 13388
rect 7932 13311 7984 13320
rect 7932 13277 7941 13311
rect 7941 13277 7975 13311
rect 7975 13277 7984 13311
rect 7932 13268 7984 13277
rect 9956 13311 10008 13320
rect 9956 13277 9965 13311
rect 9965 13277 9999 13311
rect 9999 13277 10008 13311
rect 9956 13268 10008 13277
rect 10508 13268 10560 13320
rect 5632 13132 5684 13184
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 6920 13132 6972 13184
rect 8116 13132 8168 13184
rect 8760 13200 8812 13252
rect 9404 13132 9456 13184
rect 10140 13200 10192 13252
rect 12992 13336 13044 13388
rect 13176 13336 13228 13388
rect 10416 13132 10468 13184
rect 11244 13132 11296 13184
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 11980 13132 12032 13184
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 16580 13472 16632 13524
rect 17316 13472 17368 13524
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 15660 13268 15712 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17868 13268 17920 13320
rect 14648 13200 14700 13252
rect 15108 13200 15160 13252
rect 17592 13243 17644 13252
rect 17592 13209 17601 13243
rect 17601 13209 17635 13243
rect 17635 13209 17644 13243
rect 17592 13200 17644 13209
rect 15200 13132 15252 13184
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 16948 13132 17000 13184
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 3056 12903 3108 12912
rect 3056 12869 3065 12903
rect 3065 12869 3099 12903
rect 3099 12869 3108 12903
rect 3056 12860 3108 12869
rect 3976 12860 4028 12912
rect 5632 12860 5684 12912
rect 6460 12928 6512 12980
rect 7012 12928 7064 12980
rect 8760 12928 8812 12980
rect 10140 12928 10192 12980
rect 10600 12928 10652 12980
rect 13728 12928 13780 12980
rect 2688 12724 2740 12776
rect 3884 12792 3936 12844
rect 3240 12724 3292 12776
rect 3792 12724 3844 12776
rect 6184 12792 6236 12844
rect 7932 12860 7984 12912
rect 6552 12792 6604 12844
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 8576 12792 8628 12844
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 5080 12724 5132 12776
rect 10324 12724 10376 12776
rect 11244 12767 11296 12776
rect 11244 12733 11253 12767
rect 11253 12733 11287 12767
rect 11287 12733 11296 12767
rect 11244 12724 11296 12733
rect 12808 12860 12860 12912
rect 13084 12860 13136 12912
rect 13452 12792 13504 12844
rect 14004 12928 14056 12980
rect 15660 12928 15712 12980
rect 15936 12928 15988 12980
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 3332 12588 3384 12640
rect 3884 12588 3936 12640
rect 11612 12656 11664 12708
rect 12900 12656 12952 12708
rect 13636 12656 13688 12708
rect 15108 12860 15160 12912
rect 17408 12903 17460 12912
rect 17408 12869 17417 12903
rect 17417 12869 17451 12903
rect 17451 12869 17460 12903
rect 17408 12860 17460 12869
rect 14740 12792 14792 12844
rect 15568 12792 15620 12844
rect 15844 12792 15896 12844
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 15292 12724 15344 12776
rect 17776 12724 17828 12776
rect 16580 12656 16632 12708
rect 7932 12588 7984 12640
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 9404 12588 9456 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 6552 12384 6604 12436
rect 2596 12316 2648 12368
rect 9680 12384 9732 12436
rect 13544 12384 13596 12436
rect 1584 12248 1636 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3148 12248 3200 12300
rect 3056 12180 3108 12232
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 2504 12112 2556 12164
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 4068 12180 4120 12232
rect 3976 12155 4028 12164
rect 3976 12121 3985 12155
rect 3985 12121 4019 12155
rect 4019 12121 4028 12155
rect 3976 12112 4028 12121
rect 6184 12180 6236 12232
rect 6552 12180 6604 12232
rect 6920 12180 6972 12232
rect 2596 12044 2648 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 6000 12112 6052 12164
rect 6644 12112 6696 12164
rect 6828 12155 6880 12164
rect 6828 12121 6837 12155
rect 6837 12121 6871 12155
rect 6871 12121 6880 12155
rect 6828 12112 6880 12121
rect 8024 12248 8076 12300
rect 9588 12248 9640 12300
rect 13084 12316 13136 12368
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 8116 12180 8168 12232
rect 8576 12155 8628 12164
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 9128 12223 9180 12232
rect 9128 12189 9143 12223
rect 9143 12189 9177 12223
rect 9177 12189 9180 12223
rect 9128 12180 9180 12189
rect 11980 12248 12032 12300
rect 17408 12316 17460 12368
rect 15384 12248 15436 12300
rect 17776 12248 17828 12300
rect 9864 12112 9916 12164
rect 10692 12112 10744 12164
rect 10876 12180 10928 12232
rect 11336 12180 11388 12232
rect 12808 12180 12860 12232
rect 11152 12112 11204 12164
rect 11704 12155 11756 12164
rect 11704 12121 11713 12155
rect 11713 12121 11747 12155
rect 11747 12121 11756 12155
rect 11704 12112 11756 12121
rect 11796 12155 11848 12164
rect 11796 12121 11805 12155
rect 11805 12121 11839 12155
rect 11839 12121 11848 12155
rect 11796 12112 11848 12121
rect 9956 12044 10008 12096
rect 10324 12044 10376 12096
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 10968 12087 11020 12096
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 13084 12044 13136 12096
rect 13360 12044 13412 12096
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 13636 12180 13688 12232
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14740 12180 14792 12232
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 15292 12180 15344 12232
rect 15844 12180 15896 12232
rect 16764 12180 16816 12232
rect 14556 12112 14608 12164
rect 13636 12044 13688 12096
rect 16580 12044 16632 12096
rect 17132 12044 17184 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 1676 11840 1728 11892
rect 3976 11840 4028 11892
rect 6184 11840 6236 11892
rect 7012 11840 7064 11892
rect 8944 11840 8996 11892
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 5724 11704 5776 11756
rect 2964 11568 3016 11620
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 7012 11704 7064 11756
rect 7104 11704 7156 11756
rect 8024 11772 8076 11824
rect 8116 11772 8168 11824
rect 9220 11772 9272 11824
rect 9864 11840 9916 11892
rect 11796 11840 11848 11892
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 6552 11568 6604 11620
rect 7932 11704 7984 11756
rect 6828 11500 6880 11552
rect 7748 11636 7800 11688
rect 9680 11636 9732 11688
rect 10508 11772 10560 11824
rect 10048 11704 10100 11756
rect 11336 11772 11388 11824
rect 11704 11772 11756 11824
rect 12992 11840 13044 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13544 11840 13596 11892
rect 15292 11840 15344 11892
rect 16764 11840 16816 11892
rect 10876 11704 10928 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 10048 11500 10100 11552
rect 13084 11704 13136 11756
rect 13544 11704 13596 11756
rect 13636 11704 13688 11756
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 15016 11772 15068 11824
rect 16580 11772 16632 11824
rect 17592 11772 17644 11824
rect 12624 11636 12676 11688
rect 14372 11568 14424 11620
rect 10508 11500 10560 11552
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 13176 11500 13228 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 13820 11500 13872 11552
rect 14648 11636 14700 11688
rect 15292 11636 15344 11688
rect 15844 11636 15896 11688
rect 16028 11636 16080 11688
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 1860 11296 1912 11348
rect 2412 11296 2464 11348
rect 2872 11296 2924 11348
rect 5540 11296 5592 11348
rect 5724 11296 5776 11348
rect 6460 11296 6512 11348
rect 7656 11296 7708 11348
rect 7932 11296 7984 11348
rect 10416 11296 10468 11348
rect 6736 11228 6788 11280
rect 6828 11228 6880 11280
rect 12624 11228 12676 11280
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2596 11092 2648 11144
rect 3700 11092 3752 11144
rect 4620 11160 4672 11212
rect 4988 11160 5040 11212
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 5540 11092 5592 11101
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 7012 11160 7064 11212
rect 6920 11092 6972 11144
rect 7564 11092 7616 11144
rect 2872 11024 2924 11076
rect 3332 11067 3384 11076
rect 3332 11033 3341 11067
rect 3341 11033 3375 11067
rect 3375 11033 3384 11067
rect 3332 11024 3384 11033
rect 7380 11067 7432 11076
rect 7380 11033 7389 11067
rect 7389 11033 7423 11067
rect 7423 11033 7432 11067
rect 7380 11024 7432 11033
rect 7748 11024 7800 11076
rect 8576 11092 8628 11144
rect 9404 11092 9456 11144
rect 9588 11092 9640 11144
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 10324 11092 10376 11144
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 11060 11024 11112 11076
rect 3424 10956 3476 11008
rect 3976 10956 4028 11008
rect 5356 10956 5408 11008
rect 8116 10956 8168 11008
rect 8760 10956 8812 11008
rect 9956 10956 10008 11008
rect 10876 10956 10928 11008
rect 10968 10956 11020 11008
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 14372 11228 14424 11280
rect 14740 11296 14792 11348
rect 13544 11160 13596 11212
rect 12624 11092 12676 11144
rect 14004 11092 14056 11144
rect 14556 11092 14608 11144
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 14924 11092 14976 11144
rect 16764 11160 16816 11212
rect 16948 11271 17000 11280
rect 16948 11237 16957 11271
rect 16957 11237 16991 11271
rect 16991 11237 17000 11271
rect 16948 11228 17000 11237
rect 17960 11228 18012 11280
rect 14188 11024 14240 11076
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16120 11092 16172 11144
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 17592 11092 17644 11144
rect 14464 10956 14516 11008
rect 15108 10956 15160 11008
rect 18052 11024 18104 11076
rect 18236 10999 18288 11008
rect 18236 10965 18245 10999
rect 18245 10965 18279 10999
rect 18279 10965 18288 10999
rect 18236 10956 18288 10965
rect 18420 10956 18472 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 1492 10752 1544 10804
rect 1952 10616 2004 10668
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2228 10523 2280 10532
rect 2228 10489 2237 10523
rect 2237 10489 2271 10523
rect 2271 10489 2280 10523
rect 2228 10480 2280 10489
rect 3332 10727 3384 10736
rect 3332 10693 3341 10727
rect 3341 10693 3375 10727
rect 3375 10693 3384 10727
rect 3332 10684 3384 10693
rect 4620 10684 4672 10736
rect 3424 10616 3476 10668
rect 5540 10684 5592 10736
rect 3516 10412 3568 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 8668 10752 8720 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 11428 10752 11480 10804
rect 8024 10684 8076 10736
rect 5356 10616 5408 10625
rect 6920 10548 6972 10600
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8576 10616 8628 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 5908 10480 5960 10532
rect 6828 10480 6880 10532
rect 7932 10548 7984 10600
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 8944 10548 8996 10600
rect 9772 10616 9824 10668
rect 10692 10684 10744 10736
rect 10968 10684 11020 10736
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10600 10616 10652 10668
rect 11796 10616 11848 10668
rect 14280 10752 14332 10804
rect 14372 10752 14424 10804
rect 14924 10752 14976 10804
rect 15016 10795 15068 10804
rect 15016 10761 15025 10795
rect 15025 10761 15059 10795
rect 15059 10761 15068 10795
rect 15016 10752 15068 10761
rect 15108 10752 15160 10804
rect 13084 10684 13136 10736
rect 11428 10548 11480 10600
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 13820 10684 13872 10736
rect 12900 10616 12952 10625
rect 7104 10480 7156 10532
rect 9588 10480 9640 10532
rect 9864 10480 9916 10532
rect 7932 10412 7984 10464
rect 9036 10412 9088 10464
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 15200 10616 15252 10668
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 18052 10684 18104 10736
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 16764 10659 16816 10668
rect 16764 10625 16770 10659
rect 16770 10625 16804 10659
rect 16804 10625 16816 10659
rect 16764 10616 16816 10625
rect 18236 10659 18288 10668
rect 18236 10625 18245 10659
rect 18245 10625 18279 10659
rect 18279 10625 18288 10659
rect 18236 10616 18288 10625
rect 11796 10412 11848 10464
rect 13084 10412 13136 10464
rect 13176 10412 13228 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 15476 10412 15528 10464
rect 15660 10412 15712 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 1952 10208 2004 10260
rect 2228 10140 2280 10192
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 7840 10208 7892 10260
rect 8760 10208 8812 10260
rect 9036 10208 9088 10260
rect 9220 10208 9272 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 9956 10208 10008 10260
rect 1308 10072 1360 10124
rect 3516 10115 3568 10124
rect 3516 10081 3525 10115
rect 3525 10081 3559 10115
rect 3559 10081 3568 10115
rect 3516 10072 3568 10081
rect 3976 10004 4028 10056
rect 4068 9868 4120 9920
rect 4712 9868 4764 9920
rect 6184 9979 6236 9988
rect 6184 9945 6193 9979
rect 6193 9945 6227 9979
rect 6227 9945 6236 9979
rect 6184 9936 6236 9945
rect 6276 9979 6328 9988
rect 6276 9945 6285 9979
rect 6285 9945 6319 9979
rect 6319 9945 6328 9979
rect 6276 9936 6328 9945
rect 8944 10140 8996 10192
rect 10232 10115 10284 10124
rect 7012 10004 7064 10056
rect 6736 9936 6788 9988
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 8116 10004 8168 10056
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 9312 10004 9364 10056
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 10508 10072 10560 10124
rect 11796 10140 11848 10192
rect 11888 10140 11940 10192
rect 12624 10140 12676 10192
rect 13452 10208 13504 10260
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 14004 10140 14056 10192
rect 9588 10004 9640 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10416 10004 10468 10056
rect 10968 10047 11020 10056
rect 10968 10013 10970 10047
rect 10970 10013 11004 10047
rect 11004 10013 11020 10047
rect 10968 10004 11020 10013
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 11796 10004 11848 10056
rect 12808 10004 12860 10056
rect 7104 9936 7156 9945
rect 10140 9936 10192 9988
rect 7932 9868 7984 9920
rect 13360 9936 13412 9988
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 15476 10004 15528 10056
rect 15384 9936 15436 9988
rect 16120 10004 16172 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 18328 10072 18380 10124
rect 18052 10004 18104 10056
rect 18236 9936 18288 9988
rect 11980 9868 12032 9920
rect 12624 9868 12676 9920
rect 13176 9868 13228 9920
rect 13912 9868 13964 9920
rect 14464 9868 14516 9920
rect 15568 9868 15620 9920
rect 15752 9868 15804 9920
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 1308 9664 1360 9716
rect 1216 9596 1268 9648
rect 1676 9639 1728 9648
rect 1676 9605 1685 9639
rect 1685 9605 1719 9639
rect 1719 9605 1728 9639
rect 1676 9596 1728 9605
rect 2320 9664 2372 9716
rect 3884 9596 3936 9648
rect 3976 9596 4028 9648
rect 4804 9664 4856 9716
rect 2412 9460 2464 9512
rect 3056 9528 3108 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 4620 9528 4672 9580
rect 6276 9664 6328 9716
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 9128 9664 9180 9716
rect 9312 9664 9364 9716
rect 9588 9664 9640 9716
rect 15660 9664 15712 9716
rect 7012 9596 7064 9648
rect 8024 9596 8076 9648
rect 8944 9639 8996 9648
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 9680 9596 9732 9648
rect 10324 9596 10376 9648
rect 11520 9596 11572 9648
rect 12716 9596 12768 9648
rect 7932 9528 7984 9580
rect 8668 9528 8720 9580
rect 4712 9392 4764 9444
rect 9036 9460 9088 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9772 9460 9824 9512
rect 10416 9460 10468 9512
rect 11336 9528 11388 9580
rect 11980 9528 12032 9580
rect 13268 9528 13320 9580
rect 10876 9460 10928 9512
rect 11060 9460 11112 9512
rect 11612 9460 11664 9512
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2688 9324 2740 9376
rect 3056 9324 3108 9376
rect 3700 9324 3752 9376
rect 7748 9392 7800 9444
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 7288 9324 7340 9376
rect 8852 9392 8904 9444
rect 10048 9392 10100 9444
rect 10600 9392 10652 9444
rect 11888 9392 11940 9444
rect 14280 9460 14332 9512
rect 13268 9392 13320 9444
rect 13728 9392 13780 9444
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 15476 9571 15528 9580
rect 15476 9537 15491 9571
rect 15491 9537 15525 9571
rect 15525 9537 15528 9571
rect 15476 9528 15528 9537
rect 15752 9528 15804 9580
rect 15384 9460 15436 9512
rect 11428 9324 11480 9376
rect 11704 9324 11756 9376
rect 12072 9324 12124 9376
rect 12624 9324 12676 9376
rect 13820 9324 13872 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 14372 9324 14424 9376
rect 15016 9324 15068 9376
rect 16948 9528 17000 9580
rect 16580 9460 16632 9512
rect 17224 9435 17276 9444
rect 17224 9401 17233 9435
rect 17233 9401 17267 9435
rect 17267 9401 17276 9435
rect 17224 9392 17276 9401
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 2136 9120 2188 9172
rect 3884 9120 3936 9172
rect 6184 9120 6236 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 8668 9120 8720 9172
rect 9128 9120 9180 9172
rect 3976 8916 4028 8968
rect 7288 8984 7340 9036
rect 9220 9052 9272 9104
rect 11336 9120 11388 9172
rect 10600 9052 10652 9104
rect 12716 9120 12768 9172
rect 12900 9120 12952 9172
rect 13820 9120 13872 9172
rect 14280 9163 14332 9172
rect 14280 9129 14289 9163
rect 14289 9129 14323 9163
rect 14323 9129 14332 9163
rect 14280 9120 14332 9129
rect 15200 9120 15252 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 18052 9120 18104 9172
rect 2688 8780 2740 8832
rect 4068 8891 4120 8900
rect 4068 8857 4077 8891
rect 4077 8857 4111 8891
rect 4111 8857 4120 8891
rect 4068 8848 4120 8857
rect 4804 8780 4856 8832
rect 5448 8780 5500 8832
rect 6460 8848 6512 8900
rect 7380 8848 7432 8900
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 9404 8984 9456 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 8668 8916 8720 8968
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 8852 8780 8904 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 10784 8780 10836 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 11428 8916 11480 8968
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 11704 8848 11756 8900
rect 12624 8848 12676 8900
rect 13452 8916 13504 8968
rect 13912 8984 13964 9036
rect 17224 8984 17276 9036
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 13820 8916 13872 8968
rect 15292 8916 15344 8968
rect 15476 8916 15528 8968
rect 15660 8916 15712 8968
rect 14740 8891 14792 8900
rect 14740 8857 14749 8891
rect 14749 8857 14783 8891
rect 14783 8857 14792 8891
rect 15936 8916 15988 8968
rect 16580 8916 16632 8968
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 14740 8848 14792 8857
rect 13360 8780 13412 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 2136 8576 2188 8628
rect 4068 8576 4120 8628
rect 4620 8576 4672 8628
rect 6000 8576 6052 8628
rect 1124 8508 1176 8560
rect 1584 8440 1636 8492
rect 2688 8551 2740 8560
rect 2688 8517 2697 8551
rect 2697 8517 2731 8551
rect 2731 8517 2740 8551
rect 2688 8508 2740 8517
rect 3976 8440 4028 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 7288 8576 7340 8628
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 9496 8576 9548 8628
rect 11152 8576 11204 8628
rect 11336 8576 11388 8628
rect 13176 8576 13228 8628
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 5448 8372 5500 8424
rect 4804 8304 4856 8356
rect 9588 8551 9640 8560
rect 9588 8517 9597 8551
rect 9597 8517 9631 8551
rect 9631 8517 9640 8551
rect 9588 8508 9640 8517
rect 7748 8440 7800 8492
rect 8576 8440 8628 8492
rect 9128 8440 9180 8492
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 11888 8440 11940 8492
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 7472 8304 7524 8356
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 8944 8304 8996 8313
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 11980 8304 12032 8356
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13268 8440 13320 8492
rect 12624 8372 12676 8424
rect 16948 8576 17000 8628
rect 18052 8576 18104 8628
rect 18144 8619 18196 8628
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 15844 8508 15896 8560
rect 13452 8304 13504 8356
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 14648 8440 14700 8492
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15292 8440 15344 8492
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 16028 8440 16080 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 14464 8347 14516 8356
rect 14464 8313 14473 8347
rect 14473 8313 14507 8347
rect 14507 8313 14516 8347
rect 14464 8304 14516 8313
rect 15844 8304 15896 8356
rect 13544 8236 13596 8288
rect 15108 8279 15160 8288
rect 15108 8245 15117 8279
rect 15117 8245 15151 8279
rect 15151 8245 15160 8279
rect 15108 8236 15160 8245
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 1676 8032 1728 8084
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 6920 8032 6972 8084
rect 7472 8032 7524 8084
rect 9036 8032 9088 8084
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 13452 8032 13504 8084
rect 3148 8007 3200 8016
rect 3148 7973 3157 8007
rect 3157 7973 3191 8007
rect 3191 7973 3200 8007
rect 3148 7964 3200 7973
rect 4068 7896 4120 7948
rect 7104 7896 7156 7948
rect 8116 7896 8168 7948
rect 8668 7896 8720 7948
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6552 7828 6604 7880
rect 6644 7760 6696 7812
rect 7840 7828 7892 7880
rect 8576 7828 8628 7880
rect 9128 7828 9180 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 11796 7964 11848 8016
rect 11888 7828 11940 7880
rect 15108 8032 15160 8084
rect 15200 8032 15252 8084
rect 18328 8032 18380 8084
rect 14556 7896 14608 7948
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 8024 7803 8076 7812
rect 8024 7769 8033 7803
rect 8033 7769 8067 7803
rect 8067 7769 8076 7803
rect 8024 7760 8076 7769
rect 9588 7803 9640 7812
rect 9588 7769 9597 7803
rect 9597 7769 9631 7803
rect 9631 7769 9640 7803
rect 9588 7760 9640 7769
rect 11980 7760 12032 7812
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 16120 7828 16172 7880
rect 16856 7828 16908 7880
rect 4620 7692 4672 7744
rect 4712 7692 4764 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 11060 7692 11112 7744
rect 11704 7692 11756 7744
rect 14096 7692 14148 7744
rect 15936 7760 15988 7812
rect 16580 7735 16632 7744
rect 16580 7701 16589 7735
rect 16589 7701 16623 7735
rect 16623 7701 16632 7735
rect 16580 7692 16632 7701
rect 17868 7692 17920 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 1492 7420 1544 7472
rect 7012 7488 7064 7540
rect 8024 7488 8076 7540
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 3608 7420 3660 7472
rect 4804 7352 4856 7404
rect 2780 7284 2832 7336
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 5908 7259 5960 7268
rect 5908 7225 5917 7259
rect 5917 7225 5951 7259
rect 5951 7225 5960 7259
rect 5908 7216 5960 7225
rect 6644 7420 6696 7472
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 9404 7420 9456 7472
rect 13728 7488 13780 7540
rect 10876 7420 10928 7472
rect 11704 7420 11756 7472
rect 11888 7420 11940 7472
rect 6920 7284 6972 7336
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10232 7284 10284 7336
rect 8944 7259 8996 7268
rect 8944 7225 8953 7259
rect 8953 7225 8987 7259
rect 8987 7225 8996 7259
rect 8944 7216 8996 7225
rect 12072 7352 12124 7404
rect 13360 7420 13412 7472
rect 14188 7488 14240 7540
rect 14372 7488 14424 7540
rect 14096 7420 14148 7472
rect 12992 7216 13044 7268
rect 4712 7148 4764 7200
rect 5172 7148 5224 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 6920 7148 6972 7200
rect 7012 7148 7064 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 12808 7148 12860 7200
rect 13544 7284 13596 7336
rect 15016 7488 15068 7540
rect 15752 7488 15804 7540
rect 16580 7488 16632 7540
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16856 7463 16908 7472
rect 16856 7429 16865 7463
rect 16865 7429 16899 7463
rect 16899 7429 16908 7463
rect 16856 7420 16908 7429
rect 17960 7488 18012 7540
rect 17040 7352 17092 7404
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 16028 7284 16080 7336
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 17960 7148 18012 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 3148 6944 3200 6996
rect 4804 6944 4856 6996
rect 2596 6851 2648 6860
rect 2596 6817 2605 6851
rect 2605 6817 2639 6851
rect 2639 6817 2648 6851
rect 2596 6808 2648 6817
rect 3792 6808 3844 6860
rect 5264 6944 5316 6996
rect 7012 6944 7064 6996
rect 13544 6944 13596 6996
rect 16028 6944 16080 6996
rect 17592 6944 17644 6996
rect 6552 6876 6604 6928
rect 10048 6876 10100 6928
rect 6368 6808 6420 6860
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 6920 6808 6972 6860
rect 7656 6808 7708 6860
rect 2964 6740 3016 6792
rect 4620 6740 4672 6792
rect 1768 6604 1820 6656
rect 3884 6672 3936 6724
rect 10232 6808 10284 6860
rect 11704 6808 11756 6860
rect 12808 6876 12860 6928
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 10600 6740 10652 6792
rect 10692 6740 10744 6792
rect 4988 6672 5040 6724
rect 2872 6604 2924 6656
rect 3608 6604 3660 6656
rect 7380 6672 7432 6724
rect 9864 6672 9916 6724
rect 12624 6785 12676 6792
rect 12624 6751 12633 6785
rect 12633 6751 12667 6785
rect 12667 6751 12676 6785
rect 12624 6740 12676 6751
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 14648 6808 14700 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 13084 6740 13136 6749
rect 12072 6672 12124 6724
rect 15200 6740 15252 6792
rect 15568 6783 15620 6792
rect 15568 6749 15577 6783
rect 15577 6749 15611 6783
rect 15611 6749 15620 6783
rect 15568 6740 15620 6749
rect 16120 6740 16172 6792
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 17960 6740 18012 6792
rect 7288 6604 7340 6656
rect 8576 6604 8628 6656
rect 9956 6604 10008 6656
rect 10968 6604 11020 6656
rect 15936 6604 15988 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 3608 6443 3660 6452
rect 3608 6409 3617 6443
rect 3617 6409 3651 6443
rect 3651 6409 3660 6443
rect 3608 6400 3660 6409
rect 5172 6400 5224 6452
rect 1768 6375 1820 6384
rect 1768 6341 1777 6375
rect 1777 6341 1811 6375
rect 1811 6341 1820 6375
rect 1768 6332 1820 6341
rect 7288 6400 7340 6452
rect 7380 6400 7432 6452
rect 8576 6400 8628 6452
rect 11796 6400 11848 6452
rect 12072 6400 12124 6452
rect 16948 6400 17000 6452
rect 18052 6400 18104 6452
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 2412 6196 2464 6248
rect 4068 6264 4120 6316
rect 4712 6196 4764 6248
rect 2504 6060 2556 6112
rect 3976 6128 4028 6180
rect 5172 6128 5224 6180
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 7656 6264 7708 6316
rect 7196 6171 7248 6180
rect 7196 6137 7205 6171
rect 7205 6137 7239 6171
rect 7239 6137 7248 6171
rect 7196 6128 7248 6137
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 10416 6307 10468 6316
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 12992 6264 13044 6316
rect 14096 6264 14148 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 11060 6196 11112 6248
rect 11244 6196 11296 6248
rect 13360 6196 13412 6248
rect 10876 6128 10928 6180
rect 15200 6264 15252 6316
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 4804 6060 4856 6112
rect 6368 6060 6420 6112
rect 6460 6060 6512 6112
rect 7932 6060 7984 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 12624 6060 12676 6112
rect 15292 6128 15344 6180
rect 15568 6264 15620 6316
rect 17040 6264 17092 6316
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 16120 6060 16172 6112
rect 16764 6060 16816 6112
rect 17592 6103 17644 6112
rect 17592 6069 17601 6103
rect 17601 6069 17635 6103
rect 17635 6069 17644 6103
rect 17592 6060 17644 6069
rect 17776 6060 17828 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 4068 5856 4120 5908
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 6644 5856 6696 5908
rect 7288 5856 7340 5908
rect 7656 5856 7708 5908
rect 7932 5856 7984 5908
rect 9220 5856 9272 5908
rect 10048 5856 10100 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 2504 5831 2556 5840
rect 2504 5797 2513 5831
rect 2513 5797 2547 5831
rect 2547 5797 2556 5831
rect 2504 5788 2556 5797
rect 2596 5788 2648 5840
rect 1308 5720 1360 5772
rect 3240 5720 3292 5772
rect 3792 5720 3844 5772
rect 3976 5720 4028 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2780 5652 2832 5704
rect 6460 5788 6512 5840
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 4620 5652 4672 5704
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 3424 5516 3476 5568
rect 6368 5627 6420 5636
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 8024 5788 8076 5840
rect 9772 5788 9824 5840
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 5632 5516 5684 5568
rect 7472 5516 7524 5568
rect 7932 5584 7984 5636
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 9956 5652 10008 5704
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 14648 5788 14700 5840
rect 15292 5788 15344 5840
rect 16120 5788 16172 5840
rect 13084 5720 13136 5772
rect 11612 5652 11664 5661
rect 9128 5584 9180 5636
rect 10232 5627 10284 5636
rect 10232 5593 10241 5627
rect 10241 5593 10275 5627
rect 10275 5593 10284 5627
rect 10232 5584 10284 5593
rect 10600 5584 10652 5636
rect 13176 5652 13228 5704
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17592 5856 17644 5908
rect 15384 5584 15436 5636
rect 17592 5652 17644 5704
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 10324 5516 10376 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 1676 5312 1728 5364
rect 2780 5312 2832 5364
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 3240 5312 3292 5364
rect 4620 5312 4672 5364
rect 4896 5312 4948 5364
rect 6368 5312 6420 5364
rect 7380 5312 7432 5364
rect 8576 5312 8628 5364
rect 1124 5176 1176 5228
rect 3424 5244 3476 5296
rect 3884 5244 3936 5296
rect 3608 5176 3660 5228
rect 4804 5176 4856 5228
rect 7656 5287 7708 5296
rect 7656 5253 7665 5287
rect 7665 5253 7699 5287
rect 7699 5253 7708 5287
rect 7656 5244 7708 5253
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 10232 5312 10284 5364
rect 14004 5312 14056 5364
rect 16764 5312 16816 5364
rect 17408 5312 17460 5364
rect 17592 5355 17644 5364
rect 17592 5321 17601 5355
rect 17601 5321 17635 5355
rect 17635 5321 17644 5355
rect 17592 5312 17644 5321
rect 17776 5312 17828 5364
rect 7012 5176 7064 5228
rect 7288 5176 7340 5228
rect 8760 5176 8812 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10600 5176 10652 5228
rect 11612 5209 11664 5228
rect 11612 5176 11622 5209
rect 11622 5176 11656 5209
rect 11656 5176 11664 5209
rect 14096 5244 14148 5296
rect 15384 5287 15436 5296
rect 15384 5253 15393 5287
rect 15393 5253 15427 5287
rect 15427 5253 15436 5287
rect 15384 5244 15436 5253
rect 12716 5176 12768 5228
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 6644 5108 6696 5160
rect 10416 5108 10468 5160
rect 11520 5108 11572 5160
rect 11980 5108 12032 5160
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 14188 5108 14240 5160
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16120 5108 16172 5160
rect 7196 5040 7248 5092
rect 10508 5040 10560 5092
rect 11428 5040 11480 5092
rect 16028 5040 16080 5092
rect 4068 5015 4120 5024
rect 4068 4981 4077 5015
rect 4077 4981 4111 5015
rect 4111 4981 4120 5015
rect 4068 4972 4120 4981
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 7472 4972 7524 5024
rect 9312 4972 9364 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 11888 4972 11940 5024
rect 12072 4972 12124 5024
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 1124 4768 1176 4820
rect 3792 4768 3844 4820
rect 4068 4768 4120 4820
rect 4804 4768 4856 4820
rect 2872 4632 2924 4684
rect 3884 4632 3936 4684
rect 5632 4632 5684 4684
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3608 4564 3660 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 6920 4768 6972 4820
rect 7564 4768 7616 4820
rect 8668 4768 8720 4820
rect 10508 4768 10560 4820
rect 11796 4768 11848 4820
rect 6644 4700 6696 4752
rect 13176 4768 13228 4820
rect 13636 4768 13688 4820
rect 14004 4768 14056 4820
rect 14648 4768 14700 4820
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7288 4632 7340 4684
rect 11060 4632 11112 4684
rect 7196 4564 7248 4616
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 8760 4564 8812 4616
rect 9312 4564 9364 4616
rect 2596 4428 2648 4480
rect 3056 4428 3108 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 13084 4700 13136 4752
rect 14556 4700 14608 4752
rect 11428 4564 11480 4616
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 11888 4496 11940 4548
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 12624 4496 12676 4548
rect 12716 4496 12768 4548
rect 15384 4564 15436 4616
rect 16028 4632 16080 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 16856 4564 16908 4616
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 13176 4428 13228 4480
rect 14648 4428 14700 4480
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 7932 4224 7984 4276
rect 11612 4224 11664 4276
rect 2412 4156 2464 4208
rect 3148 4088 3200 4140
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 3056 4020 3108 4072
rect 3424 3952 3476 4004
rect 5448 4088 5500 4140
rect 5724 4020 5776 4072
rect 5356 3952 5408 4004
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 8116 4088 8168 4140
rect 10232 4156 10284 4208
rect 8576 4088 8628 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 7012 4020 7064 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 11796 4156 11848 4208
rect 10876 4088 10928 4140
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 14188 4224 14240 4276
rect 14556 4224 14608 4276
rect 14648 4224 14700 4276
rect 16856 4224 16908 4276
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11244 4020 11296 4072
rect 11796 4020 11848 4072
rect 13176 4156 13228 4208
rect 12624 4088 12676 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 14924 4156 14976 4208
rect 6736 3952 6788 4004
rect 2504 3884 2556 3936
rect 12808 3952 12860 4004
rect 15292 4020 15344 4072
rect 16120 4020 16172 4072
rect 17316 4020 17368 4072
rect 15568 3995 15620 4004
rect 15568 3961 15577 3995
rect 15577 3961 15611 3995
rect 15611 3961 15620 3995
rect 15568 3952 15620 3961
rect 7104 3884 7156 3936
rect 9772 3884 9824 3936
rect 10508 3884 10560 3936
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 11980 3884 12032 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1768 3680 1820 3732
rect 3148 3680 3200 3732
rect 3240 3680 3292 3732
rect 3976 3680 4028 3732
rect 6828 3680 6880 3732
rect 8116 3680 8168 3732
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 10140 3680 10192 3732
rect 11152 3680 11204 3732
rect 940 3476 992 3528
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 2780 3476 2832 3528
rect 3240 3476 3292 3528
rect 6368 3612 6420 3664
rect 6460 3612 6512 3664
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 2412 3408 2464 3460
rect 3332 3451 3384 3460
rect 3332 3417 3341 3451
rect 3341 3417 3375 3451
rect 3375 3417 3384 3451
rect 3332 3408 3384 3417
rect 4804 3476 4856 3528
rect 4620 3408 4672 3460
rect 7104 3544 7156 3596
rect 6644 3476 6696 3528
rect 8760 3476 8812 3528
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 12808 3680 12860 3732
rect 13084 3680 13136 3732
rect 15568 3680 15620 3732
rect 15660 3680 15712 3732
rect 15936 3680 15988 3732
rect 17868 3680 17920 3732
rect 10692 3544 10744 3596
rect 12624 3612 12676 3664
rect 2872 3340 2924 3392
rect 3516 3340 3568 3392
rect 4896 3340 4948 3392
rect 5540 3340 5592 3392
rect 6736 3340 6788 3392
rect 11520 3476 11572 3528
rect 12716 3544 12768 3596
rect 12072 3408 12124 3460
rect 10968 3340 11020 3392
rect 11244 3340 11296 3392
rect 14004 3476 14056 3528
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14924 3476 14976 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 13176 3383 13228 3392
rect 13176 3349 13185 3383
rect 13185 3349 13219 3383
rect 13219 3349 13228 3383
rect 13176 3340 13228 3349
rect 17592 3340 17644 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 5448 3136 5500 3188
rect 6368 3136 6420 3188
rect 1860 2932 1912 2984
rect 3332 2932 3384 2984
rect 3976 3000 4028 3052
rect 4896 3000 4948 3052
rect 4620 2864 4672 2916
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 7748 3136 7800 3188
rect 8116 3136 8168 3188
rect 7472 3068 7524 3120
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 10784 3136 10836 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 10968 3136 11020 3188
rect 11796 3136 11848 3188
rect 6276 2932 6328 2984
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 7932 3000 7984 3052
rect 8576 3068 8628 3120
rect 9312 3068 9364 3120
rect 10048 3068 10100 3120
rect 13176 3136 13228 3188
rect 14924 3136 14976 3188
rect 15752 3136 15804 3188
rect 13912 3068 13964 3120
rect 14556 3068 14608 3120
rect 10324 3000 10376 3052
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 10692 3000 10744 3052
rect 11704 3000 11756 3052
rect 11060 2932 11112 2984
rect 12072 2932 12124 2984
rect 15292 3043 15344 3052
rect 15292 3009 15301 3043
rect 15301 3009 15335 3043
rect 15335 3009 15344 3043
rect 15292 3000 15344 3009
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 9036 2864 9088 2916
rect 10692 2864 10744 2916
rect 11244 2864 11296 2916
rect 8576 2796 8628 2848
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 12072 2839 12124 2848
rect 12072 2805 12081 2839
rect 12081 2805 12115 2839
rect 12115 2805 12124 2839
rect 12072 2796 12124 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 3884 2592 3936 2644
rect 4620 2592 4672 2644
rect 6736 2592 6788 2644
rect 7012 2592 7064 2644
rect 2412 2456 2464 2508
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 2044 2388 2096 2440
rect 3332 2388 3384 2440
rect 4712 2524 4764 2576
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 5448 2456 5500 2508
rect 5632 2388 5684 2440
rect 7932 2524 7984 2576
rect 9036 2592 9088 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 9220 2456 9272 2508
rect 4804 2320 4856 2372
rect 8668 2388 8720 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10968 2592 11020 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 12072 2592 12124 2644
rect 11796 2567 11848 2576
rect 11796 2533 11805 2567
rect 11805 2533 11839 2567
rect 11839 2533 11848 2567
rect 11796 2524 11848 2533
rect 12808 2456 12860 2508
rect 13452 2456 13504 2508
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 10232 2320 10284 2372
rect 10416 2320 10468 2372
rect 11704 2388 11756 2440
rect 2320 2252 2372 2304
rect 7656 2252 7708 2304
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 11980 2252 12032 2304
rect 12900 2320 12952 2372
rect 14096 2320 14148 2372
rect 14464 2363 14516 2372
rect 14464 2329 14473 2363
rect 14473 2329 14507 2363
rect 14507 2329 14516 2363
rect 14464 2320 14516 2329
rect 16948 2252 17000 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 1860 2048 1912 2100
rect 3424 1980 3476 2032
rect 3148 1887 3200 1896
rect 3148 1853 3157 1887
rect 3157 1853 3191 1887
rect 3191 1853 3200 1887
rect 3148 1844 3200 1853
rect 7012 2048 7064 2100
rect 7932 2048 7984 2100
rect 9680 2048 9732 2100
rect 10048 2048 10100 2100
rect 10232 2048 10284 2100
rect 9312 2023 9364 2032
rect 9312 1989 9321 2023
rect 9321 1989 9355 2023
rect 9355 1989 9364 2023
rect 9312 1980 9364 1989
rect 6920 1955 6972 1964
rect 6920 1921 6929 1955
rect 6929 1921 6963 1955
rect 6963 1921 6972 1955
rect 6920 1912 6972 1921
rect 7012 1955 7064 1964
rect 7012 1921 7021 1955
rect 7021 1921 7055 1955
rect 7055 1921 7064 1955
rect 7012 1912 7064 1921
rect 5448 1844 5500 1896
rect 6368 1844 6420 1896
rect 2780 1708 2832 1760
rect 3332 1708 3384 1760
rect 3792 1751 3844 1760
rect 3792 1717 3801 1751
rect 3801 1717 3835 1751
rect 3835 1717 3844 1751
rect 3792 1708 3844 1717
rect 6644 1776 6696 1828
rect 8024 1844 8076 1896
rect 10416 1980 10468 2032
rect 11704 2091 11756 2100
rect 11704 2057 11713 2091
rect 11713 2057 11747 2091
rect 11747 2057 11756 2091
rect 11704 2048 11756 2057
rect 11796 2048 11848 2100
rect 11060 1980 11112 2032
rect 14464 2048 14516 2100
rect 12900 1980 12952 2032
rect 13912 1980 13964 2032
rect 14924 1980 14976 2032
rect 17592 2023 17644 2032
rect 17592 1989 17601 2023
rect 17601 1989 17635 2023
rect 17635 1989 17644 2023
rect 17592 1980 17644 1989
rect 10968 1912 11020 1964
rect 13452 1955 13504 1964
rect 13452 1921 13461 1955
rect 13461 1921 13495 1955
rect 13495 1921 13504 1955
rect 13452 1912 13504 1921
rect 13544 1912 13596 1964
rect 14096 1912 14148 1964
rect 16120 1912 16172 1964
rect 16948 1912 17000 1964
rect 8760 1776 8812 1828
rect 9680 1819 9732 1828
rect 9680 1785 9689 1819
rect 9689 1785 9723 1819
rect 9723 1785 9732 1819
rect 9680 1776 9732 1785
rect 10140 1751 10192 1760
rect 10140 1717 10149 1751
rect 10149 1717 10183 1751
rect 10183 1717 10192 1751
rect 10140 1708 10192 1717
rect 11796 1776 11848 1828
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2320 1547 2372 1556
rect 2320 1513 2329 1547
rect 2329 1513 2363 1547
rect 2363 1513 2372 1547
rect 2320 1504 2372 1513
rect 3240 1504 3292 1556
rect 6368 1504 6420 1556
rect 2872 1300 2924 1352
rect 3056 1300 3108 1352
rect 3516 1436 3568 1488
rect 3424 1300 3476 1352
rect 3792 1232 3844 1284
rect 7012 1504 7064 1556
rect 7748 1504 7800 1556
rect 9680 1504 9732 1556
rect 11152 1504 11204 1556
rect 11796 1436 11848 1488
rect 11980 1436 12032 1488
rect 16120 1547 16172 1556
rect 16120 1513 16129 1547
rect 16129 1513 16163 1547
rect 16163 1513 16172 1547
rect 16120 1504 16172 1513
rect 16948 1504 17000 1556
rect 5448 1368 5500 1420
rect 5816 1368 5868 1420
rect 6920 1368 6972 1420
rect 8024 1368 8076 1420
rect 10140 1368 10192 1420
rect 13452 1368 13504 1420
rect 7656 1232 7708 1284
rect 8760 1232 8812 1284
rect 13544 1232 13596 1284
rect 13912 1232 13964 1284
rect 1860 1207 1912 1216
rect 1860 1173 1869 1207
rect 1869 1173 1903 1207
rect 1903 1173 1912 1207
rect 1860 1164 1912 1173
rect 3148 1164 3200 1216
rect 10968 1164 11020 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
rect 1860 960 1912 1012
rect 5632 960 5684 1012
<< metal2 >>
rect 1122 14200 1178 15000
rect 2594 14362 2650 15000
rect 2594 14334 2728 14362
rect 2594 14200 2650 14334
rect 1136 13734 1164 14200
rect 1124 13728 1176 13734
rect 1124 13670 1176 13676
rect 1030 13424 1086 13433
rect 1030 13359 1032 13368
rect 1084 13359 1086 13368
rect 1492 13388 1544 13394
rect 1032 13330 1084 13336
rect 1492 13330 1544 13336
rect 1504 10810 1532 13330
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 1582 12744 1638 12753
rect 1582 12679 1638 12688
rect 1596 12306 1624 12679
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1688 12238 1716 12582
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11898 1716 12038
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1872 11354 1900 13126
rect 2516 12170 2544 13126
rect 2700 12782 2728 14334
rect 4066 14200 4122 15000
rect 5538 14200 5594 15000
rect 7010 14200 7066 15000
rect 8482 14362 8538 15000
rect 9954 14362 10010 15000
rect 8482 14334 8892 14362
rect 8482 14200 8538 14334
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 2688 12776 2740 12782
rect 2740 12724 2820 12730
rect 2688 12718 2820 12724
rect 2700 12702 2820 12718
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11801 2544 12106
rect 2608 12102 2636 12310
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2502 11792 2558 11801
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2412 11756 2464 11762
rect 2502 11727 2558 11736
rect 2412 11698 2464 11704
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10985 1716 11086
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1964 10674 1992 11698
rect 2424 11354 2452 11698
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2608 11150 2636 12038
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 1964 10266 1992 10610
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2240 10198 2268 10474
rect 2228 10192 2280 10198
rect 1306 10160 1362 10169
rect 2228 10134 2280 10140
rect 1306 10095 1308 10104
rect 1360 10095 1362 10104
rect 1308 10066 1360 10072
rect 1320 9722 1348 10066
rect 2332 9722 2360 10610
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 1216 9648 1268 9654
rect 1216 9590 1268 9596
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1228 9353 1256 9590
rect 1214 9344 1270 9353
rect 1214 9279 1270 9288
rect 1122 8664 1178 8673
rect 1122 8599 1178 8608
rect 1136 8566 1164 8599
rect 1124 8560 1176 8566
rect 1124 8502 1176 8508
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8090 1624 8434
rect 1688 8090 1716 9590
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2148 9178 2176 9318
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2148 8634 2176 9114
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2424 8090 2452 9454
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 8838 2728 9318
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8566 2728 8774
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2792 8090 2820 12702
rect 3068 12238 3096 12854
rect 3252 12782 3280 13126
rect 3896 12850 3924 13330
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12918 4016 13194
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3792 12776 3844 12782
rect 3844 12724 3924 12730
rect 3792 12718 3924 12724
rect 3804 12702 3924 12718
rect 3896 12646 3924 12702
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11354 2912 12038
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2976 11234 3004 11562
rect 2884 11206 3004 11234
rect 2884 11082 2912 11206
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1504 6254 1532 7414
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 7002 1992 7346
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1780 6390 1808 6598
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1320 5778 1348 6015
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1122 5264 1178 5273
rect 1122 5199 1124 5208
rect 1176 5199 1178 5208
rect 1124 5170 1176 5176
rect 1136 4826 1164 5170
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 952 3534 980 4111
rect 1504 4078 1532 6190
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5370 1716 5646
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 2424 4214 2452 6190
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 5846 2544 6054
rect 2608 5846 2636 6802
rect 2792 6202 2820 7278
rect 2884 6662 2912 11018
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3068 9382 3096 9522
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3160 8022 3188 12242
rect 3344 12238 3372 12582
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11937 3464 12038
rect 3422 11928 3478 11937
rect 3422 11863 3478 11872
rect 3896 11762 3924 12582
rect 4080 12238 4108 14200
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4208 13626 4528 13648
rect 4208 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 4528 13626
rect 4208 12538 4528 13574
rect 4208 12486 4214 12538
rect 4266 12518 4278 12538
rect 4330 12518 4342 12538
rect 4394 12518 4406 12538
rect 4458 12518 4470 12538
rect 4276 12486 4278 12518
rect 4458 12486 4460 12518
rect 4522 12486 4528 12538
rect 4208 12462 4220 12486
rect 4276 12462 4300 12486
rect 4356 12462 4380 12486
rect 4436 12462 4460 12486
rect 4516 12462 4528 12486
rect 4208 12438 4528 12462
rect 4208 12382 4220 12438
rect 4276 12382 4300 12438
rect 4356 12382 4380 12438
rect 4436 12382 4460 12438
rect 4516 12382 4528 12438
rect 4208 12358 4528 12382
rect 4208 12302 4220 12358
rect 4276 12302 4300 12358
rect 4356 12302 4380 12358
rect 4436 12302 4460 12358
rect 4516 12302 4528 12358
rect 4208 12278 4528 12302
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4208 12222 4220 12278
rect 4276 12222 4300 12278
rect 4356 12222 4380 12278
rect 4436 12222 4460 12278
rect 4516 12222 4528 12278
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3988 11898 4016 12106
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4208 11450 4528 12222
rect 4208 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 4528 11450
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 10742 3372 11018
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3436 10674 3464 10950
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3712 10470 3740 11086
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3528 10130 3556 10406
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3422 9616 3478 9625
rect 3422 9551 3424 9560
rect 3476 9551 3478 9560
rect 3424 9522 3476 9528
rect 3712 9382 3740 10406
rect 3988 10062 4016 10950
rect 4208 10362 4528 11398
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10742 4660 11154
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4208 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 4528 10362
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9654 4016 9998
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3976 9648 4028 9654
rect 4080 9625 4108 9862
rect 3976 9590 4028 9596
rect 4066 9616 4122 9625
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3896 9178 3924 9590
rect 4066 9551 4122 9560
rect 4208 9274 4528 10310
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4208 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 4528 9274
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8498 4016 8910
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8634 4108 8842
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4208 8186 4528 9222
rect 4632 8634 4660 9522
rect 4724 9450 4752 9862
rect 4816 9722 4844 13670
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12782 5120 13262
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5092 12442 5120 12718
rect 5080 12436 5132 12442
rect 5552 12434 5580 14200
rect 7024 13462 7052 14200
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 13530 7236 13738
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5644 12918 5672 13126
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5552 12406 5948 12434
rect 5080 12378 5132 12384
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5000 11218 5028 11630
rect 5552 11354 5580 11630
rect 5736 11354 5764 11698
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10674 5396 10950
rect 5552 10742 5580 11086
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5552 10266 5580 10678
rect 5920 10538 5948 12406
rect 6012 12170 6040 13126
rect 6472 12986 6500 13262
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6184 12844 6236 12850
rect 6552 12844 6604 12850
rect 6184 12786 6236 12792
rect 6472 12804 6552 12832
rect 6196 12238 6224 12786
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6472 11354 6500 12804
rect 6552 12786 6604 12792
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6564 12238 6592 12378
rect 6932 12238 6960 13126
rect 7024 12986 7052 13398
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7944 12918 7972 13262
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6644 12164 6696 12170
rect 6828 12164 6880 12170
rect 6696 12124 6828 12152
rect 6644 12106 6696 12112
rect 6828 12106 6880 12112
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7024 11762 7052 11834
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6644 11688 6696 11694
rect 6642 11656 6644 11665
rect 6696 11656 6698 11665
rect 6552 11620 6604 11626
rect 6642 11591 6698 11600
rect 6552 11562 6604 11568
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6564 11150 6592 11562
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11286 6868 11494
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 6748 9994 6776 11222
rect 7024 11218 7052 11698
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10606 6960 11086
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7116 10538 7144 11698
rect 7392 11082 7420 12786
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 11354 7696 12174
rect 7944 11762 7972 12582
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11830 8064 12242
rect 8128 12238 8156 13126
rect 8208 13082 8528 13648
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8208 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 8528 13082
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11830 8156 12174
rect 8208 11994 8528 13030
rect 8772 12986 8800 13194
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8588 12170 8616 12786
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8208 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 8528 11994
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7748 11688 7800 11694
rect 7746 11656 7748 11665
rect 7800 11656 7802 11665
rect 7746 11591 7802 11600
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7576 10810 7604 11086
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7760 10674 7788 11018
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7944 10606 7972 11290
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6840 10305 6868 10474
rect 6826 10296 6882 10305
rect 6826 10231 6882 10240
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 5262 9616 5318 9625
rect 4804 9580 4856 9586
rect 5262 9551 5264 9560
rect 4804 9522 4856 9528
rect 5316 9551 5318 9560
rect 5264 9522 5316 9528
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4816 8838 4844 9522
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4816 8362 4844 8774
rect 5460 8430 5488 8774
rect 6012 8634 6040 9318
rect 6196 9178 6224 9930
rect 6288 9722 6316 9930
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 7024 9654 7052 9998
rect 7116 9994 7144 10474
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6472 8906 6500 9522
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 4208 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 4528 8186
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4080 7721 4108 7890
rect 4066 7712 4122 7721
rect 4066 7647 4122 7656
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3160 7002 3188 7278
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2792 6174 2912 6202
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5370 2820 5646
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2884 5250 2912 6174
rect 2976 5370 3004 6734
rect 3620 6662 3648 7414
rect 4208 7098 4528 8134
rect 5736 7886 5764 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4208 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 4528 7098
rect 3882 6896 3938 6905
rect 3792 6860 3844 6866
rect 3882 6831 3938 6840
rect 3792 6802 3844 6808
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6458 3648 6598
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5778 3280 6054
rect 3804 5778 3832 6802
rect 3896 6730 3924 6831
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5778 4016 6122
rect 4080 5914 4108 6258
rect 4208 6010 4528 7046
rect 4632 6798 4660 7686
rect 4724 7206 4752 7686
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4724 6254 4752 7142
rect 4816 7002 4844 7346
rect 5920 7274 5948 8434
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4208 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 4528 6010
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3252 5370 3280 5714
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3436 5302 3464 5510
rect 3424 5296 3476 5302
rect 2884 5222 3004 5250
rect 3424 5238 3476 5244
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1780 3738 1808 4014
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 2424 3466 2452 4150
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1872 2446 1900 2926
rect 2056 2446 2084 2994
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2516 2802 2544 3878
rect 2608 3534 2636 4422
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2780 3528 2832 3534
rect 2884 3516 2912 4626
rect 2832 3488 2912 3516
rect 2780 3470 2832 3476
rect 2884 3398 2912 3488
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2870 2816 2926 2825
rect 2424 2514 2452 2790
rect 2516 2774 2820 2802
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 1872 2106 1900 2382
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 2332 1562 2360 2246
rect 2792 1766 2820 2774
rect 2870 2751 2926 2760
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 2320 1556 2372 1562
rect 2320 1498 2372 1504
rect 2884 1358 2912 2751
rect 2976 2009 3004 5222
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 4622 3648 5170
rect 3804 4826 3832 5714
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3896 4690 3924 5238
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4208 4922 4528 5958
rect 4816 5778 4844 6054
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5370 4660 5646
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4816 5234 4844 5714
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4908 5370 4936 5646
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4208 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 4528 4922
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3068 4078 3096 4422
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3160 3738 3188 4082
rect 3252 3738 3280 4422
rect 3436 4010 3464 4558
rect 3620 4282 3648 4558
rect 4208 4518 4528 4870
rect 4816 4826 4844 4966
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4208 4462 4220 4518
rect 4276 4462 4300 4518
rect 4356 4462 4380 4518
rect 4436 4462 4460 4518
rect 4516 4462 4528 4518
rect 4208 4438 4528 4462
rect 4208 4382 4220 4438
rect 4276 4382 4300 4438
rect 4356 4382 4380 4438
rect 4436 4382 4460 4438
rect 4516 4382 4528 4438
rect 4208 4358 4528 4382
rect 4208 4302 4220 4358
rect 4276 4302 4300 4358
rect 4356 4302 4380 4358
rect 4436 4302 4460 4358
rect 4516 4302 4528 4358
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 4208 4278 4528 4302
rect 4208 4222 4220 4278
rect 4276 4222 4300 4278
rect 4356 4222 4380 4278
rect 4436 4222 4460 4278
rect 4516 4222 4528 4278
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 4208 3834 4528 4222
rect 4208 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 4528 3834
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3054 3632 3110 3641
rect 3054 3567 3110 3576
rect 2962 2000 3018 2009
rect 2962 1935 3018 1944
rect 3068 1358 3096 3567
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3252 3346 3280 3470
rect 3332 3460 3384 3466
rect 3384 3420 3464 3448
rect 3332 3402 3384 3408
rect 3252 3318 3372 3346
rect 3344 2990 3372 3318
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3344 2446 3372 2926
rect 3436 2514 3464 3420
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3344 1952 3372 2382
rect 3436 2038 3464 2450
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3252 1924 3372 1952
rect 3148 1896 3200 1902
rect 3148 1838 3200 1844
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 3056 1352 3108 1358
rect 3056 1294 3108 1300
rect 3160 1222 3188 1838
rect 3252 1562 3280 1924
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 1860 1216 1912 1222
rect 1860 1158 1912 1164
rect 3148 1216 3200 1222
rect 3344 1193 3372 1702
rect 3528 1494 3556 3334
rect 3988 3058 4016 3674
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3988 2774 4016 2994
rect 3896 2746 4016 2774
rect 4208 2746 4528 3782
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4632 3074 4660 3402
rect 4632 3046 4752 3074
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 3896 2650 3924 2746
rect 4208 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 4528 2746
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3792 1760 3844 1766
rect 3792 1702 3844 1708
rect 3516 1488 3568 1494
rect 3436 1436 3516 1442
rect 3436 1430 3568 1436
rect 3436 1414 3556 1430
rect 3436 1358 3464 1414
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3804 1290 3832 1702
rect 4208 1658 4528 2694
rect 4632 2650 4660 2858
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4724 2582 4752 3046
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 2378 4844 3470
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4208 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 4528 1658
rect 3792 1284 3844 1290
rect 3792 1226 3844 1232
rect 3148 1158 3200 1164
rect 3330 1184 3386 1193
rect 1872 1018 1900 1158
rect 3330 1119 3386 1128
rect 4208 1040 4528 1606
rect 1860 1012 1912 1018
rect 1860 954 1912 960
rect 5000 800 5028 6666
rect 5184 6458 5212 7142
rect 5276 7002 5304 7142
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 6380 6866 6408 7822
rect 6564 6934 6592 7822
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7478 6684 7754
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6656 6866 6684 7414
rect 6932 7342 6960 8026
rect 7116 7954 7144 9930
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9042 7328 9318
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8634 7328 8978
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 8634 7420 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7760 8498 7788 9386
rect 7852 8974 7880 10202
rect 7944 9926 7972 10406
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8036 9654 8064 10678
rect 8128 10062 8156 10950
rect 8208 10906 8528 11942
rect 8576 11144 8628 11150
rect 8628 11104 8708 11132
rect 8576 11086 8628 11092
rect 8208 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 8528 10906
rect 8116 10056 8168 10062
rect 8114 10024 8116 10033
rect 8168 10024 8170 10033
rect 8114 9959 8170 9968
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 9178 7972 9522
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 8090 7512 8298
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7852 7886 7880 8366
rect 8128 7954 8156 9959
rect 8208 9818 8528 10854
rect 8680 10810 8708 11104
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8208 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 8528 9818
rect 8208 8730 8528 9766
rect 8588 9674 8616 10610
rect 8680 10062 8708 10610
rect 8772 10266 8800 10950
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8588 9646 8800 9674
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 9178 8708 9522
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8208 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 8528 8730
rect 8208 8518 8528 8678
rect 8208 8462 8220 8518
rect 8276 8462 8300 8518
rect 8356 8462 8380 8518
rect 8436 8462 8460 8518
rect 8516 8462 8528 8518
rect 8208 8438 8528 8462
rect 8208 8382 8220 8438
rect 8276 8382 8300 8438
rect 8356 8382 8380 8438
rect 8436 8382 8460 8438
rect 8516 8382 8528 8438
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8208 8358 8528 8382
rect 8208 8302 8220 8358
rect 8276 8302 8300 8358
rect 8356 8302 8380 8358
rect 8436 8302 8460 8358
rect 8516 8302 8528 8358
rect 8208 8278 8528 8302
rect 8208 8222 8220 8278
rect 8276 8222 8300 8278
rect 8356 8222 8380 8278
rect 8436 8222 8460 8278
rect 8516 8222 8528 8278
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7546 7052 7686
rect 8036 7546 8064 7754
rect 8208 7642 8528 8222
rect 8588 7886 8616 8434
rect 8680 7954 8708 8910
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8208 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 8528 7642
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6932 6866 6960 7142
rect 7024 7002 7052 7142
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5184 6186 5212 6394
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6380 5914 6408 6054
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6472 5846 6500 6054
rect 6656 5914 6684 6258
rect 7208 6186 7236 7346
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6458 7328 6598
rect 7392 6458 7420 6666
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7300 5914 7328 6394
rect 7668 6322 7696 6802
rect 8208 6554 8528 7590
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8208 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 8528 6554
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 4690 5672 5510
rect 6380 5370 6408 5578
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6656 4758 6684 5102
rect 6932 4826 6960 5646
rect 7392 5370 7420 6258
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5914 7972 6054
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5368 3602 5396 3946
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5460 3194 5488 4082
rect 5736 4078 5764 4558
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5552 3058 5580 3334
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 6288 2990 6316 4558
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6380 3194 6408 3606
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6472 3058 6500 3606
rect 6656 3534 6684 4694
rect 7024 4078 7052 5170
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4622 7236 5034
rect 7300 4690 7328 5170
rect 7484 5030 7512 5510
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7484 4146 7512 4966
rect 7576 4826 7604 5646
rect 7668 5302 7696 5850
rect 8024 5840 8076 5846
rect 7944 5788 8024 5794
rect 7944 5782 8076 5788
rect 7944 5766 8064 5782
rect 7944 5642 7972 5766
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 8128 4622 8156 5510
rect 8208 5466 8528 6502
rect 8588 6458 8616 6598
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8588 6322 8616 6394
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8208 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 8528 5466
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7944 4282 7972 4558
rect 8208 4378 8528 5414
rect 8588 5370 8616 6258
rect 8772 5386 8800 9646
rect 8864 9636 8892 14334
rect 9954 14334 10272 14362
rect 9954 14200 10010 14334
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12646 9444 13126
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8942 11928 8998 11937
rect 8942 11863 8944 11872
rect 8996 11863 8998 11872
rect 8944 11834 8996 11840
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 10198 8984 10542
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10266 9076 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 9140 9722 9168 12174
rect 9232 11830 9260 12582
rect 9680 12436 9732 12442
rect 9968 12424 9996 13262
rect 10060 12594 10088 13466
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 12986 10180 13194
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10060 12566 10180 12594
rect 9732 12396 9996 12424
rect 9680 12378 9732 12384
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9600 12073 9628 12242
rect 10152 12186 10180 12566
rect 9876 12170 10180 12186
rect 9864 12164 10180 12170
rect 9916 12158 10180 12164
rect 9864 12106 9916 12112
rect 9956 12096 10008 12102
rect 9586 12064 9642 12073
rect 9956 12038 10008 12044
rect 9586 11999 9642 12008
rect 9862 11928 9918 11937
rect 9862 11863 9864 11872
rect 9916 11863 9918 11872
rect 9864 11834 9916 11840
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9968 11744 9996 12038
rect 10048 11756 10100 11762
rect 9968 11716 10048 11744
rect 10048 11698 10100 11704
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9232 10266 9260 10610
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9416 10169 9444 11086
rect 9600 10985 9628 11086
rect 9586 10976 9642 10985
rect 9586 10911 9642 10920
rect 9600 10538 9628 10911
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9402 10160 9458 10169
rect 9402 10095 9458 10104
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9722 9352 9998
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8944 9648 8996 9654
rect 8864 9608 8944 9636
rect 8944 9590 8996 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8864 8838 8892 9386
rect 9048 9058 9076 9454
rect 9140 9178 9168 9454
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9220 9104 9272 9110
rect 9048 9052 9220 9058
rect 9048 9046 9272 9052
rect 9048 9030 9260 9046
rect 9416 9042 9444 10095
rect 9588 10056 9640 10062
rect 9586 10024 9588 10033
rect 9640 10024 9642 10033
rect 9586 9959 9642 9968
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9600 9042 9628 9658
rect 9692 9654 9720 11630
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11082 10088 11494
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9784 10062 9812 10610
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9876 10266 9904 10474
rect 9968 10266 9996 10610
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 10152 9994 10180 10610
rect 10244 10130 10272 14334
rect 11426 14200 11482 15000
rect 12898 14200 12954 15000
rect 14370 14200 14426 15000
rect 15842 14200 15898 15000
rect 17314 14200 17370 15000
rect 18786 14200 18842 15000
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13462 11284 13670
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12102 10364 12718
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10428 11354 10456 13126
rect 10520 12186 10548 13262
rect 10612 12986 10640 13330
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 11256 12782 11284 13126
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11440 12434 11468 14200
rect 12208 13626 12528 13648
rect 12208 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 12528 13626
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12850 12020 13126
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11440 12406 11560 12434
rect 10876 12232 10928 12238
rect 10520 12158 10640 12186
rect 10876 12174 10928 12180
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11830 10548 12038
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10336 9654 10364 11086
rect 10520 10130 10548 11494
rect 10612 10674 10640 12158
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11937 10732 12106
rect 10690 11928 10746 11937
rect 10690 11863 10746 11872
rect 10888 11762 10916 12174
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11801 11008 12038
rect 10966 11792 11022 11801
rect 10876 11756 10928 11762
rect 10796 11716 10876 11744
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 10742 10732 11494
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10428 9518 10456 9998
rect 9772 9512 9824 9518
rect 9770 9480 9772 9489
rect 10416 9512 10468 9518
rect 9824 9480 9826 9489
rect 10416 9454 10468 9460
rect 9770 9415 9826 9424
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8956 7274 8984 8298
rect 9048 8090 9076 8366
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9140 7886 9168 8434
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7410 9168 7822
rect 9416 7478 9444 8774
rect 9508 8634 9536 8774
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9600 7818 9628 8502
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 10060 6934 10088 9386
rect 10520 7562 10548 10066
rect 10796 9674 10824 11716
rect 10966 11727 11022 11736
rect 10876 11698 10928 11704
rect 11164 11665 11192 12106
rect 11348 11830 11376 12174
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11150 11656 11206 11665
rect 11150 11591 11206 11600
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10968 11008 11020 11014
rect 11072 10985 11100 11018
rect 10968 10950 11020 10956
rect 11058 10976 11114 10985
rect 10888 10554 10916 10950
rect 10980 10742 11008 10950
rect 11058 10911 11114 10920
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 11348 10690 11376 11766
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10810 11468 11086
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11348 10662 11468 10690
rect 11440 10606 11468 10662
rect 11428 10600 11480 10606
rect 10966 10568 11022 10577
rect 10888 10526 10966 10554
rect 11428 10542 11480 10548
rect 10966 10503 11022 10512
rect 10980 10062 11008 10503
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10796 9646 10916 9674
rect 10888 9518 10916 9646
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 9110 10640 9386
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 7886 10824 8774
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10520 7534 10640 7562
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10244 6866 10272 7278
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9232 5914 9260 6258
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8680 5358 8800 5386
rect 9140 5370 9168 5578
rect 9128 5364 9180 5370
rect 8680 4826 8708 5358
rect 9128 5306 9180 5312
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8772 4622 8800 5170
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4622 9352 4966
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 8208 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 8528 4378
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 1902 5488 2450
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 5460 1426 5488 1838
rect 5448 1420 5500 1426
rect 5448 1362 5500 1368
rect 5644 1018 5672 2382
rect 5828 1426 5856 2518
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6380 1562 6408 1838
rect 6656 1834 6684 3470
rect 6748 3398 6776 3946
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 2650 6776 3334
rect 7024 2650 7052 4014
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 3602 7144 3878
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7484 3126 7512 4082
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7760 3194 7788 4014
rect 8128 3738 8156 4082
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8128 3194 8156 3674
rect 8208 3290 8528 4326
rect 9324 4146 9352 4558
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8208 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 8528 3290
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7024 2106 7052 2586
rect 7944 2582 7972 2994
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 6644 1828 6696 1834
rect 6644 1770 6696 1776
rect 6368 1556 6420 1562
rect 6368 1498 6420 1504
rect 6932 1426 6960 1906
rect 7024 1562 7052 1906
rect 7012 1556 7064 1562
rect 7012 1498 7064 1504
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 7668 1290 7696 2246
rect 7760 1562 7788 2246
rect 7944 2106 7972 2518
rect 8208 2202 8528 3238
rect 8588 3126 8616 4082
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8588 2854 8616 3062
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8680 2446 8708 4082
rect 9324 3738 9352 4082
rect 9784 3942 9812 5782
rect 9876 5710 9904 6666
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 5710 9996 6598
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10060 5914 10088 6054
rect 10152 5914 10180 6054
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10244 5370 10272 5578
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 4214 10272 5170
rect 10232 4208 10284 4214
rect 10152 4168 10232 4196
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 10152 3738 10180 4168
rect 10232 4150 10284 4156
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 3194 8800 3470
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 10048 3120 10100 3126
rect 10152 3108 10180 3674
rect 10100 3080 10180 3108
rect 10048 3062 10100 3068
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9048 2650 9076 2858
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9232 2514 9260 2790
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8208 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 8528 2202
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 8036 1426 8064 1838
rect 8024 1420 8076 1426
rect 8024 1362 8076 1368
rect 7656 1284 7708 1290
rect 7656 1226 7708 1232
rect 8208 1114 8528 2150
rect 9324 2038 9352 3062
rect 10336 3058 10364 5510
rect 10428 5166 10456 6258
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10520 5098 10548 7346
rect 10612 6798 10640 7534
rect 10888 7478 10916 9454
rect 11072 7750 11100 9454
rect 11348 9178 11376 9522
rect 11440 9382 11468 10542
rect 11532 9654 11560 12406
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11624 9518 11652 12650
rect 11992 12306 12020 12786
rect 12208 12538 12528 13574
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12208 12486 12214 12538
rect 12266 12518 12278 12538
rect 12330 12518 12342 12538
rect 12394 12518 12406 12538
rect 12458 12518 12470 12538
rect 12276 12486 12278 12518
rect 12458 12486 12460 12518
rect 12522 12486 12528 12538
rect 12208 12462 12220 12486
rect 12276 12462 12300 12486
rect 12356 12462 12380 12486
rect 12436 12462 12460 12486
rect 12516 12462 12528 12486
rect 12208 12438 12528 12462
rect 12208 12382 12220 12438
rect 12276 12382 12300 12438
rect 12356 12382 12380 12438
rect 12436 12382 12460 12438
rect 12516 12382 12528 12438
rect 12208 12358 12528 12382
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12208 12302 12220 12358
rect 12276 12302 12300 12358
rect 12356 12302 12380 12358
rect 12436 12302 12460 12358
rect 12516 12302 12528 12358
rect 12208 12278 12528 12302
rect 12208 12222 12220 12278
rect 12276 12222 12300 12278
rect 12356 12222 12380 12278
rect 12436 12222 12460 12278
rect 12516 12222 12528 12278
rect 12820 12238 12848 12854
rect 12912 12714 12940 14200
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11716 11830 11744 12106
rect 11808 11898 11836 12106
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10470 11836 10610
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10198 11836 10406
rect 11886 10296 11942 10305
rect 11886 10231 11942 10240
rect 11900 10198 11928 10231
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8634 11192 8774
rect 11348 8634 11376 9114
rect 11440 8974 11468 9318
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11716 8906 11744 9318
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11808 8480 11836 9998
rect 11992 9926 12020 11698
rect 12208 11450 12528 12222
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13004 12050 13032 13330
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12918 13124 13126
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13084 12368 13136 12374
rect 13188 12356 13216 13330
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12434 13492 12786
rect 13556 12442 13584 13126
rect 13740 12986 13768 13262
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13136 12328 13216 12356
rect 13280 12406 13492 12434
rect 13544 12436 13596 12442
rect 13084 12310 13136 12316
rect 13280 12186 13308 12406
rect 13544 12378 13596 12384
rect 13648 12238 13676 12650
rect 13544 12232 13596 12238
rect 13280 12158 13492 12186
rect 13544 12174 13596 12180
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 12728 12022 13032 12050
rect 13084 12096 13136 12102
rect 13360 12096 13412 12102
rect 13084 12038 13136 12044
rect 13280 12056 13360 12084
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12208 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 12528 11450
rect 12208 10362 12528 11398
rect 12636 11286 12664 11630
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12208 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 12528 10362
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11886 9480 11942 9489
rect 11886 9415 11888 9424
rect 11940 9415 11942 9424
rect 11888 9386 11940 9392
rect 11888 8492 11940 8498
rect 11808 8452 11888 8480
rect 11888 8434 11940 8440
rect 11796 8016 11848 8022
rect 11900 8004 11928 8434
rect 11992 8362 12020 9522
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9042 12112 9318
rect 12208 9274 12528 10310
rect 12636 10198 12664 11086
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9382 12664 9862
rect 12728 9654 12756 12022
rect 12990 11928 13046 11937
rect 13096 11898 13124 12038
rect 12990 11863 12992 11872
rect 13044 11863 13046 11872
rect 13084 11892 13136 11898
rect 12992 11834 13044 11840
rect 13084 11834 13136 11840
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13096 10742 13124 11698
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12806 10160 12862 10169
rect 12806 10095 12862 10104
rect 12820 10062 12848 10095
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12208 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 12528 9274
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11848 7976 11928 8004
rect 11796 7958 11848 7964
rect 11900 7886 11928 7976
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 6798 10732 7142
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10874 6216 10930 6225
rect 10874 6151 10876 6160
rect 10928 6151 10930 6160
rect 10876 6122 10928 6128
rect 10980 6118 11008 6598
rect 11072 6254 11100 7686
rect 11716 7478 11744 7686
rect 11900 7478 11928 7822
rect 11992 7818 12020 8298
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12084 7410 12112 8434
rect 12208 8186 12528 9222
rect 12728 9178 12756 9590
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12716 8968 12768 8974
rect 12622 8936 12678 8945
rect 12716 8910 12768 8916
rect 12622 8871 12624 8880
rect 12676 8871 12678 8880
rect 12624 8842 12676 8848
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12208 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 12528 8186
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11060 6248 11112 6254
rect 11244 6248 11296 6254
rect 11060 6190 11112 6196
rect 11164 6208 11244 6236
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10612 5234 10640 5578
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10508 4820 10560 4826
rect 10612 4808 10640 5170
rect 10560 4780 10640 4808
rect 10508 4762 10560 4768
rect 11164 4706 11192 6208
rect 11244 6190 11296 6196
rect 11716 5914 11744 6802
rect 12084 6730 12112 7346
rect 12208 7098 12528 8134
rect 12208 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 12528 7098
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12084 6458 12112 6666
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11808 5914 11836 6394
rect 12208 6010 12528 7046
rect 12636 6798 12664 8366
rect 12728 6866 12756 8910
rect 12820 8090 12848 9998
rect 12912 9178 12940 10610
rect 13188 10606 13216 11494
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13188 10470 13216 10542
rect 13084 10464 13136 10470
rect 13082 10432 13084 10441
rect 13176 10464 13228 10470
rect 13136 10432 13138 10441
rect 13176 10406 13228 10412
rect 13082 10367 13138 10376
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13096 8498 13124 10367
rect 13188 9926 13216 10406
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 8634 13216 9862
rect 13280 9586 13308 12056
rect 13360 12038 13412 12044
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13372 9994 13400 11154
rect 13464 10266 13492 12158
rect 13556 11898 13584 12174
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11937 13676 12038
rect 13634 11928 13690 11937
rect 13544 11892 13596 11898
rect 13634 11863 13690 11872
rect 13544 11834 13596 11840
rect 14016 11762 14044 12922
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13556 11529 13584 11698
rect 13648 11558 13676 11698
rect 13636 11552 13688 11558
rect 13542 11520 13598 11529
rect 13636 11494 13688 11500
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13542 11455 13598 11464
rect 13542 11248 13598 11257
rect 13542 11183 13544 11192
rect 13596 11183 13598 11192
rect 13544 11154 13596 11160
rect 13832 10742 13860 11494
rect 14016 11150 14044 11698
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10554 13768 10610
rect 13740 10526 13860 10554
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13636 10056 13688 10062
rect 13450 10024 13506 10033
rect 13360 9988 13412 9994
rect 13506 10004 13636 10010
rect 13506 9998 13688 10004
rect 13506 9982 13676 9998
rect 13450 9959 13506 9968
rect 13360 9930 13412 9936
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13648 9466 13676 9982
rect 13648 9450 13768 9466
rect 13268 9444 13320 9450
rect 13648 9444 13780 9450
rect 13648 9438 13728 9444
rect 13268 9386 13320 9392
rect 13728 9386 13780 9392
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13280 8498 13308 9386
rect 13832 9382 13860 10526
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9178 13860 9318
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13924 9042 13952 9862
rect 14016 9586 14044 10134
rect 14200 10130 14228 11018
rect 14292 10810 14320 12174
rect 14384 11744 14412 14200
rect 15856 13938 15884 14200
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14568 11801 14596 12106
rect 14554 11792 14610 11801
rect 14384 11716 14504 11744
rect 14554 11727 14610 11736
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 11286 14412 11562
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14384 10810 14412 11222
rect 14476 11014 14504 11716
rect 14660 11694 14688 13194
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14752 12238 14780 12786
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 11552 14608 11558
rect 14554 11520 14556 11529
rect 14608 11520 14610 11529
rect 14554 11455 14610 11464
rect 14752 11354 14780 12174
rect 15028 11830 15056 13874
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15212 13433 15240 13738
rect 15198 13424 15254 13433
rect 15198 13359 15254 13368
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15120 12918 15148 13194
rect 15212 13190 15240 13359
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15120 12238 15148 12854
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 12238 15332 12718
rect 15396 12306 15424 13126
rect 15580 12850 15608 13262
rect 15672 12986 15700 13262
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12986 15976 13126
rect 16208 13082 16528 13648
rect 17328 13530 17356 14200
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 16208 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 16528 13082
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15856 12238 15884 12786
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15304 11898 15332 12174
rect 16208 11994 16528 13030
rect 16592 12714 16620 13466
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16776 12238 16804 12786
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16208 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 16528 11994
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10690 14596 11086
rect 14384 10662 14596 10690
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14384 10010 14412 10662
rect 14462 10568 14518 10577
rect 14844 10554 14872 11086
rect 14936 10810 14964 11086
rect 15028 10810 15056 11766
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 15304 11257 15332 11630
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 14518 10526 14872 10554
rect 14462 10503 14518 10512
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14108 9982 14412 10010
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13084 8492 13136 8498
rect 13004 8452 13084 8480
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 13004 7274 13032 8452
rect 13084 8434 13136 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13372 8090 13400 8774
rect 13464 8362 13492 8910
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13464 8090 13492 8298
rect 13556 8294 13584 8774
rect 13740 8634 13768 8910
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8514 13860 8910
rect 13740 8486 13860 8514
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13740 7546 13768 8486
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6934 12848 7142
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 13004 6882 13032 7210
rect 12716 6860 12768 6866
rect 13004 6854 13216 6882
rect 12716 6802 12768 6808
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 13004 6225 13032 6258
rect 12990 6216 13046 6225
rect 12990 6151 13046 6160
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12208 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 12528 6010
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11624 5234 11652 5646
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11072 4690 11192 4706
rect 11060 4684 11192 4690
rect 11112 4678 11192 4684
rect 11060 4626 11112 4632
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10520 3210 10548 3878
rect 10704 3602 10732 3878
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10520 3182 10732 3210
rect 10796 3194 10824 4014
rect 10888 3194 10916 4082
rect 11164 3738 11192 4678
rect 11440 4622 11468 5034
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4078 11284 4422
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11532 3534 11560 5102
rect 11624 4282 11652 5170
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11808 4826 11836 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11808 4214 11836 4558
rect 11900 4554 11928 4966
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11808 3738 11836 4014
rect 11992 3942 12020 5102
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4146 12112 4966
rect 12208 4922 12528 5958
rect 12636 5522 12664 6054
rect 13096 5778 13124 6734
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12636 5494 12756 5522
rect 12728 5234 12756 5494
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12208 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 12528 4922
rect 12208 4518 12528 4870
rect 12728 4554 12756 5170
rect 13096 4758 13124 5714
rect 13188 5710 13216 6854
rect 13372 6254 13400 7414
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 7002 13584 7278
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 4826 13216 5510
rect 13372 5234 13400 6190
rect 14016 5370 14044 9522
rect 14108 9382 14136 9982
rect 14476 9926 14504 10406
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14292 9178 14320 9454
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14384 8430 14412 9318
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7478 14136 7686
rect 14200 7546 14228 7822
rect 14384 7546 14412 8366
rect 14476 8362 14504 9862
rect 14752 8906 14780 10526
rect 15212 10441 15240 10610
rect 15198 10432 15254 10441
rect 15198 10367 15254 10376
rect 15396 9994 15424 10610
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15488 10062 15516 10406
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15488 9874 15516 9998
rect 15396 9846 15516 9874
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14556 7948 14608 7954
rect 14660 7936 14688 8434
rect 14608 7908 14688 7936
rect 14556 7890 14608 7896
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14108 6322 14136 7414
rect 14660 6866 14688 7908
rect 15028 7546 15056 9318
rect 15212 9178 15240 9522
rect 15396 9518 15424 9846
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15488 9178 15516 9522
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 9058 15608 9862
rect 15672 9722 15700 10406
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15488 9030 15608 9058
rect 15488 8974 15516 9030
rect 15672 8974 15700 9658
rect 15764 9586 15792 9862
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15304 8498 15332 8910
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 8090 15148 8230
rect 15212 8090 15240 8434
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15212 6798 15240 7278
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15212 6322 15240 6734
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13648 4826 13676 5102
rect 14016 4826 14044 5306
rect 14108 5302 14136 6258
rect 14660 5846 14688 6258
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 5846 15332 6122
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15396 5302 15424 5578
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12208 4462 12220 4518
rect 12276 4462 12300 4518
rect 12356 4462 12380 4518
rect 12436 4462 12460 4518
rect 12516 4462 12528 4518
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12208 4438 12528 4462
rect 12208 4382 12220 4438
rect 12276 4382 12300 4438
rect 12356 4382 12380 4438
rect 12436 4382 12460 4438
rect 12516 4382 12528 4438
rect 12208 4358 12528 4382
rect 12208 4302 12220 4358
rect 12276 4302 12300 4358
rect 12356 4302 12380 4358
rect 12436 4302 12460 4358
rect 12516 4302 12528 4358
rect 12208 4278 12528 4302
rect 12208 4222 12220 4278
rect 12276 4222 12300 4278
rect 12356 4222 12380 4278
rect 12436 4222 12460 4278
rect 12516 4222 12528 4278
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 12208 3834 12528 4222
rect 12636 4146 12664 4490
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12208 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 12528 3834
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 10980 3194 11008 3334
rect 10704 3058 10732 3182
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10612 2774 10640 2994
rect 10704 2922 10732 2994
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10428 2746 10640 2774
rect 10428 2650 10456 2746
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 2106 9720 2382
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10060 2106 10088 2246
rect 10244 2106 10272 2314
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10428 2038 10456 2314
rect 9312 2032 9364 2038
rect 9312 1974 9364 1980
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10980 1970 11008 2586
rect 11072 2038 11100 2926
rect 11256 2922 11284 3334
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 2650 11284 2858
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11716 2446 11744 2994
rect 11808 2582 11836 3130
rect 12084 2990 12112 3402
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 2650 12112 2790
rect 12208 2746 12528 3782
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12636 2990 12664 3606
rect 12728 3602 12756 4490
rect 13096 4146 13124 4694
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4214 13216 4422
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12820 3738 12848 3946
rect 13096 3738 13124 4082
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 14016 3534 14044 4762
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 3194 13216 3334
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 12624 2984 12676 2990
rect 12676 2944 12848 2972
rect 12624 2926 12676 2932
rect 12208 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 12528 2746
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 8760 1828 8812 1834
rect 8760 1770 8812 1776
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 8772 1290 8800 1770
rect 9692 1562 9720 1770
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 10152 1426 10180 1702
rect 10140 1420 10192 1426
rect 10140 1362 10192 1368
rect 8760 1284 8812 1290
rect 8760 1226 8812 1232
rect 10980 1222 11008 1906
rect 11164 1562 11192 2382
rect 11716 2106 11744 2382
rect 11808 2106 11836 2518
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11704 2100 11756 2106
rect 11704 2042 11756 2048
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11808 1834 11836 2042
rect 11796 1828 11848 1834
rect 11796 1770 11848 1776
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 11808 1494 11836 1770
rect 11992 1494 12020 2246
rect 12208 1658 12528 2694
rect 12820 2514 12848 2944
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12912 2038 12940 2314
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 13464 1970 13492 2450
rect 13924 2038 13952 3062
rect 14108 2378 14136 5238
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4282 14228 5102
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14384 3534 14412 4558
rect 14568 4282 14596 4694
rect 14660 4486 14688 4762
rect 15396 4622 15424 5238
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14660 4282 14688 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14568 3126 14596 4218
rect 14936 4214 14964 4422
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14936 3534 14964 4150
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14936 3194 14964 3470
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 15304 3058 15332 4014
rect 15488 3641 15516 8910
rect 15764 7546 15792 9522
rect 15856 8673 15884 11630
rect 16040 11150 16068 11630
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16040 10674 16068 11086
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16132 10062 16160 11086
rect 16208 10906 16528 11942
rect 16592 11830 16620 12038
rect 16776 11898 16804 12174
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16960 11286 16988 13126
rect 17144 12102 17172 13262
rect 17420 12918 17448 13670
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17420 12374 17448 12854
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17604 11830 17632 13194
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16208 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 16528 10906
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16208 9818 16528 10854
rect 16776 10674 16804 11154
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16960 10062 16988 11222
rect 17604 11150 17632 11766
rect 17696 11744 17724 12786
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12306 17816 12718
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17776 11756 17828 11762
rect 17696 11716 17776 11744
rect 17776 11698 17828 11704
rect 17788 11665 17816 11698
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17880 11218 17908 13262
rect 18800 12073 18828 14200
rect 18786 12064 18842 12073
rect 18786 11999 18842 12008
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 16208 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 16528 9818
rect 15936 8968 15988 8974
rect 15934 8936 15936 8945
rect 15988 8936 15990 8945
rect 15934 8871 15990 8880
rect 16208 8730 16528 9766
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16592 8974 16620 9454
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16208 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 16528 8730
rect 15842 8664 15898 8673
rect 15842 8599 15898 8608
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 16208 8518 16528 8678
rect 16960 8634 16988 9522
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 9042 17264 9386
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17880 8974 17908 9862
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 15856 8362 15884 8502
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16208 8462 16220 8518
rect 16276 8462 16300 8518
rect 16356 8462 16380 8518
rect 16436 8462 16460 8518
rect 16516 8462 16528 8518
rect 17880 8498 17908 8910
rect 16208 8438 16528 8462
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15580 6322 15608 6734
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15580 3738 15608 3946
rect 15672 3738 15700 4422
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15474 3632 15530 3641
rect 15474 3567 15530 3576
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15764 3194 15792 3470
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 13912 2032 13964 2038
rect 13912 1974 13964 1980
rect 13452 1964 13504 1970
rect 13452 1906 13504 1912
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 12208 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 12528 1658
rect 11796 1488 11848 1494
rect 11796 1430 11848 1436
rect 11980 1488 12032 1494
rect 11980 1430 12032 1436
rect 10968 1216 11020 1222
rect 10968 1158 11020 1164
rect 8208 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 8528 1114
rect 8208 1040 8528 1062
rect 12208 1040 12528 1606
rect 13464 1426 13492 1906
rect 13452 1420 13504 1426
rect 13452 1362 13504 1368
rect 13556 1290 13584 1906
rect 13924 1290 13952 1974
rect 14108 1970 14136 2314
rect 14476 2106 14504 2314
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14924 2032 14976 2038
rect 14924 1974 14976 1980
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 13544 1284 13596 1290
rect 13544 1226 13596 1232
rect 13912 1284 13964 1290
rect 13912 1226 13964 1232
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 14936 800 14964 1974
rect 15856 1193 15884 8298
rect 15948 7818 15976 8434
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7410 15976 7754
rect 16040 7698 16068 8434
rect 16208 8382 16220 8438
rect 16276 8382 16300 8438
rect 16356 8382 16380 8438
rect 16436 8382 16460 8438
rect 16516 8382 16528 8438
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 16208 8358 16528 8382
rect 16208 8302 16220 8358
rect 16276 8302 16300 8358
rect 16356 8302 16380 8358
rect 16436 8302 16460 8358
rect 16516 8302 16528 8358
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16208 8278 16528 8302
rect 16132 7886 16160 8230
rect 16208 8222 16220 8278
rect 16276 8222 16300 8278
rect 16356 8222 16380 8278
rect 16436 8222 16460 8278
rect 16516 8222 16528 8278
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16040 7670 16160 7698
rect 16132 7410 16160 7670
rect 16208 7642 16528 8222
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16208 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 16528 7642
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 7002 16068 7278
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16132 6798 16160 7346
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 5710 15976 6598
rect 16208 6554 16528 7590
rect 16592 7546 16620 7686
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16868 7478 16896 7822
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16208 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 16528 6554
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5846 16160 6054
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 16208 5466 16528 6502
rect 16684 5914 16712 6734
rect 16776 6118 16804 6734
rect 16960 6458 16988 6802
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17052 6322 17080 7346
rect 17604 7002 17632 7890
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16208 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 16528 5466
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15948 3738 15976 5170
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 4690 16068 5034
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16132 4078 16160 5102
rect 16208 4378 16528 5414
rect 16776 5370 16804 6054
rect 17420 5370 17448 6190
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17776 6112 17828 6118
rect 17880 6089 17908 7686
rect 17972 7546 18000 11222
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10742 18092 11018
rect 18236 11008 18288 11014
rect 18420 11008 18472 11014
rect 18236 10950 18288 10956
rect 18418 10976 18420 10985
rect 18472 10976 18474 10985
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18064 10062 18092 10678
rect 18248 10674 18276 10950
rect 18418 10911 18474 10920
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18248 9994 18276 10610
rect 18432 10266 18460 10911
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 9178 18092 9386
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18064 8634 18092 9114
rect 18156 8634 18184 9454
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18248 7410 18276 9930
rect 18340 8090 18368 10066
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6798 18000 7142
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18064 6458 18092 6802
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17776 6054 17828 6060
rect 17866 6080 17922 6089
rect 17604 5914 17632 6054
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5370 17632 5646
rect 17788 5370 17816 6054
rect 17866 6015 17922 6024
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4622 16896 4966
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16208 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 16528 4378
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16208 3290 16528 4326
rect 16868 4282 16896 4558
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 17328 4078 17356 4626
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17880 3738 17908 4558
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 16208 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 16528 3290
rect 16208 2202 16528 3238
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16208 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 16528 2202
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16132 1562 16160 1906
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 15842 1184 15898 1193
rect 15842 1119 15898 1128
rect 16208 1114 16528 2150
rect 16960 1970 16988 2246
rect 17604 2038 17632 3334
rect 17592 2032 17644 2038
rect 17592 1974 17644 1980
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 16960 1562 16988 1906
rect 16948 1556 17000 1562
rect 16948 1498 17000 1504
rect 16208 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 16528 1114
rect 16208 1040 16528 1062
rect 4986 0 5042 800
rect 14922 0 14978 800
<< via2 >>
rect 1030 13388 1086 13424
rect 1030 13368 1032 13388
rect 1032 13368 1084 13388
rect 1084 13368 1086 13388
rect 1582 12688 1638 12744
rect 2502 11736 2558 11792
rect 1674 10920 1730 10976
rect 1306 10124 1362 10160
rect 1306 10104 1308 10124
rect 1308 10104 1360 10124
rect 1360 10104 1362 10124
rect 1214 9288 1270 9344
rect 1122 8608 1178 8664
rect 1306 6024 1362 6080
rect 1122 5228 1178 5264
rect 1122 5208 1124 5228
rect 1124 5208 1176 5228
rect 1176 5208 1178 5228
rect 938 4120 994 4176
rect 3422 11872 3478 11928
rect 4220 12486 4266 12518
rect 4266 12486 4276 12518
rect 4300 12486 4330 12518
rect 4330 12486 4342 12518
rect 4342 12486 4356 12518
rect 4380 12486 4394 12518
rect 4394 12486 4406 12518
rect 4406 12486 4436 12518
rect 4460 12486 4470 12518
rect 4470 12486 4516 12518
rect 4220 12462 4276 12486
rect 4300 12462 4356 12486
rect 4380 12462 4436 12486
rect 4460 12462 4516 12486
rect 4220 12382 4276 12438
rect 4300 12382 4356 12438
rect 4380 12382 4436 12438
rect 4460 12382 4516 12438
rect 4220 12302 4276 12358
rect 4300 12302 4356 12358
rect 4380 12302 4436 12358
rect 4460 12302 4516 12358
rect 4220 12222 4276 12278
rect 4300 12222 4356 12278
rect 4380 12222 4436 12278
rect 4460 12222 4516 12278
rect 3422 9580 3478 9616
rect 3422 9560 3424 9580
rect 3424 9560 3476 9580
rect 3476 9560 3478 9580
rect 4066 9560 4122 9616
rect 6642 11636 6644 11656
rect 6644 11636 6696 11656
rect 6696 11636 6698 11656
rect 6642 11600 6698 11636
rect 7746 11636 7748 11656
rect 7748 11636 7800 11656
rect 7800 11636 7802 11656
rect 7746 11600 7802 11636
rect 6826 10240 6882 10296
rect 5262 9580 5318 9616
rect 5262 9560 5264 9580
rect 5264 9560 5316 9580
rect 5316 9560 5318 9580
rect 4066 7656 4122 7712
rect 3882 6840 3938 6896
rect 2870 2760 2926 2816
rect 4220 4462 4276 4518
rect 4300 4462 4356 4518
rect 4380 4462 4436 4518
rect 4460 4462 4516 4518
rect 4220 4382 4276 4438
rect 4300 4382 4356 4438
rect 4380 4382 4436 4438
rect 4460 4382 4516 4438
rect 4220 4302 4276 4358
rect 4300 4302 4356 4358
rect 4380 4302 4436 4358
rect 4460 4302 4516 4358
rect 4220 4222 4276 4278
rect 4300 4222 4356 4278
rect 4380 4222 4436 4278
rect 4460 4222 4516 4278
rect 3054 3576 3110 3632
rect 2962 1944 3018 2000
rect 3330 1128 3386 1184
rect 8114 10004 8116 10024
rect 8116 10004 8168 10024
rect 8168 10004 8170 10024
rect 8114 9968 8170 10004
rect 8220 8462 8276 8518
rect 8300 8462 8356 8518
rect 8380 8462 8436 8518
rect 8460 8462 8516 8518
rect 8220 8382 8276 8438
rect 8300 8382 8356 8438
rect 8380 8382 8436 8438
rect 8460 8382 8516 8438
rect 8220 8302 8276 8358
rect 8300 8302 8356 8358
rect 8380 8302 8436 8358
rect 8460 8302 8516 8358
rect 8220 8222 8276 8278
rect 8300 8222 8356 8278
rect 8380 8222 8436 8278
rect 8460 8222 8516 8278
rect 8942 11892 8998 11928
rect 8942 11872 8944 11892
rect 8944 11872 8996 11892
rect 8996 11872 8998 11892
rect 9586 12008 9642 12064
rect 9862 11892 9918 11928
rect 9862 11872 9864 11892
rect 9864 11872 9916 11892
rect 9916 11872 9918 11892
rect 9586 10920 9642 10976
rect 9402 10104 9458 10160
rect 9586 10004 9588 10024
rect 9588 10004 9640 10024
rect 9640 10004 9642 10024
rect 9586 9968 9642 10004
rect 10690 11872 10746 11928
rect 9770 9460 9772 9480
rect 9772 9460 9824 9480
rect 9824 9460 9826 9480
rect 9770 9424 9826 9460
rect 10966 11736 11022 11792
rect 11150 11600 11206 11656
rect 11058 10920 11114 10976
rect 10966 10512 11022 10568
rect 12220 12486 12266 12518
rect 12266 12486 12276 12518
rect 12300 12486 12330 12518
rect 12330 12486 12342 12518
rect 12342 12486 12356 12518
rect 12380 12486 12394 12518
rect 12394 12486 12406 12518
rect 12406 12486 12436 12518
rect 12460 12486 12470 12518
rect 12470 12486 12516 12518
rect 12220 12462 12276 12486
rect 12300 12462 12356 12486
rect 12380 12462 12436 12486
rect 12460 12462 12516 12486
rect 12220 12382 12276 12438
rect 12300 12382 12356 12438
rect 12380 12382 12436 12438
rect 12460 12382 12516 12438
rect 12220 12302 12276 12358
rect 12300 12302 12356 12358
rect 12380 12302 12436 12358
rect 12460 12302 12516 12358
rect 12220 12222 12276 12278
rect 12300 12222 12356 12278
rect 12380 12222 12436 12278
rect 12460 12222 12516 12278
rect 11886 10240 11942 10296
rect 11886 9444 11942 9480
rect 11886 9424 11888 9444
rect 11888 9424 11940 9444
rect 11940 9424 11942 9444
rect 12990 11892 13046 11928
rect 12990 11872 12992 11892
rect 12992 11872 13044 11892
rect 13044 11872 13046 11892
rect 12806 10104 12862 10160
rect 10874 6180 10930 6216
rect 10874 6160 10876 6180
rect 10876 6160 10928 6180
rect 10928 6160 10930 6180
rect 12622 8900 12678 8936
rect 12622 8880 12624 8900
rect 12624 8880 12676 8900
rect 12676 8880 12678 8900
rect 13082 10412 13084 10432
rect 13084 10412 13136 10432
rect 13136 10412 13138 10432
rect 13082 10376 13138 10412
rect 13634 11872 13690 11928
rect 13542 11464 13598 11520
rect 13542 11212 13598 11248
rect 13542 11192 13544 11212
rect 13544 11192 13596 11212
rect 13596 11192 13598 11212
rect 13450 9968 13506 10024
rect 14554 11736 14610 11792
rect 14554 11500 14556 11520
rect 14556 11500 14608 11520
rect 14608 11500 14610 11520
rect 14554 11464 14610 11500
rect 15198 13368 15254 13424
rect 14462 10512 14518 10568
rect 15290 11192 15346 11248
rect 12990 6160 13046 6216
rect 15198 10376 15254 10432
rect 12220 4462 12276 4518
rect 12300 4462 12356 4518
rect 12380 4462 12436 4518
rect 12460 4462 12516 4518
rect 12220 4382 12276 4438
rect 12300 4382 12356 4438
rect 12380 4382 12436 4438
rect 12460 4382 12516 4438
rect 12220 4302 12276 4358
rect 12300 4302 12356 4358
rect 12380 4302 12436 4358
rect 12460 4302 12516 4358
rect 12220 4222 12276 4278
rect 12300 4222 12356 4278
rect 12380 4222 12436 4278
rect 12460 4222 12516 4278
rect 17774 11600 17830 11656
rect 18786 12008 18842 12064
rect 15934 8916 15936 8936
rect 15936 8916 15988 8936
rect 15988 8916 15990 8936
rect 15934 8880 15990 8916
rect 15842 8608 15898 8664
rect 16220 8462 16276 8518
rect 16300 8462 16356 8518
rect 16380 8462 16436 8518
rect 16460 8462 16516 8518
rect 15474 3576 15530 3632
rect 16220 8382 16276 8438
rect 16300 8382 16356 8438
rect 16380 8382 16436 8438
rect 16460 8382 16516 8438
rect 16220 8302 16276 8358
rect 16300 8302 16356 8358
rect 16380 8302 16436 8358
rect 16460 8302 16516 8358
rect 16220 8222 16276 8278
rect 16300 8222 16356 8278
rect 16380 8222 16436 8278
rect 16460 8222 16516 8278
rect 18418 10956 18420 10976
rect 18420 10956 18472 10976
rect 18472 10956 18474 10976
rect 18418 10920 18474 10956
rect 17866 6024 17922 6080
rect 15842 1128 15898 1184
<< metal3 >>
rect 0 13426 800 13456
rect 1025 13426 1091 13429
rect 0 13424 1091 13426
rect 0 13368 1030 13424
rect 1086 13368 1091 13424
rect 0 13366 1091 13368
rect 0 13336 800 13366
rect 1025 13363 1091 13366
rect 15193 13426 15259 13429
rect 19200 13426 20000 13456
rect 15193 13424 20000 13426
rect 15193 13368 15198 13424
rect 15254 13368 20000 13424
rect 15193 13366 20000 13368
rect 15193 13363 15259 13366
rect 19200 13336 20000 13366
rect 1577 12746 1643 12749
rect 798 12744 1643 12746
rect 798 12688 1582 12744
rect 1638 12688 1643 12744
rect 798 12686 1643 12688
rect 798 12640 858 12686
rect 1577 12683 1643 12686
rect 0 12550 858 12640
rect 0 12520 800 12550
rect 1056 12518 18908 12530
rect 1056 12462 4220 12518
rect 4276 12462 4300 12518
rect 4356 12462 4380 12518
rect 4436 12462 4460 12518
rect 4516 12462 12220 12518
rect 12276 12462 12300 12518
rect 12356 12462 12380 12518
rect 12436 12462 12460 12518
rect 12516 12462 18908 12518
rect 1056 12438 18908 12462
rect 1056 12382 4220 12438
rect 4276 12382 4300 12438
rect 4356 12382 4380 12438
rect 4436 12382 4460 12438
rect 4516 12382 12220 12438
rect 12276 12382 12300 12438
rect 12356 12382 12380 12438
rect 12436 12382 12460 12438
rect 12516 12382 18908 12438
rect 1056 12358 18908 12382
rect 1056 12302 4220 12358
rect 4276 12302 4300 12358
rect 4356 12302 4380 12358
rect 4436 12302 4460 12358
rect 4516 12302 12220 12358
rect 12276 12302 12300 12358
rect 12356 12302 12380 12358
rect 12436 12302 12460 12358
rect 12516 12302 18908 12358
rect 1056 12278 18908 12302
rect 1056 12222 4220 12278
rect 4276 12222 4300 12278
rect 4356 12222 4380 12278
rect 4436 12222 4460 12278
rect 4516 12222 12220 12278
rect 12276 12222 12300 12278
rect 12356 12222 12380 12278
rect 12436 12222 12460 12278
rect 12516 12222 18908 12278
rect 1056 12210 18908 12222
rect 9581 12066 9647 12069
rect 18781 12066 18847 12069
rect 9581 12064 18847 12066
rect 9581 12008 9586 12064
rect 9642 12008 18786 12064
rect 18842 12008 18847 12064
rect 9581 12006 18847 12008
rect 9581 12003 9647 12006
rect 18781 12003 18847 12006
rect 3417 11930 3483 11933
rect 8937 11930 9003 11933
rect 3417 11928 9003 11930
rect 3417 11872 3422 11928
rect 3478 11872 8942 11928
rect 8998 11872 9003 11928
rect 3417 11870 9003 11872
rect 3417 11867 3483 11870
rect 8937 11867 9003 11870
rect 9857 11930 9923 11933
rect 10685 11930 10751 11933
rect 9857 11928 10751 11930
rect 9857 11872 9862 11928
rect 9918 11872 10690 11928
rect 10746 11872 10751 11928
rect 9857 11870 10751 11872
rect 9857 11867 9923 11870
rect 10685 11867 10751 11870
rect 12985 11930 13051 11933
rect 13629 11930 13695 11933
rect 12985 11928 13695 11930
rect 12985 11872 12990 11928
rect 13046 11872 13634 11928
rect 13690 11872 13695 11928
rect 12985 11870 13695 11872
rect 12985 11867 13051 11870
rect 13629 11867 13695 11870
rect 0 11794 800 11824
rect 2497 11794 2563 11797
rect 0 11792 2563 11794
rect 0 11736 2502 11792
rect 2558 11736 2563 11792
rect 0 11734 2563 11736
rect 0 11704 800 11734
rect 2497 11731 2563 11734
rect 10961 11794 11027 11797
rect 14549 11794 14615 11797
rect 10961 11792 14615 11794
rect 10961 11736 10966 11792
rect 11022 11736 14554 11792
rect 14610 11736 14615 11792
rect 10961 11734 14615 11736
rect 10961 11731 11027 11734
rect 14549 11731 14615 11734
rect 6637 11658 6703 11661
rect 7741 11658 7807 11661
rect 6637 11656 7807 11658
rect 6637 11600 6642 11656
rect 6698 11600 7746 11656
rect 7802 11600 7807 11656
rect 6637 11598 7807 11600
rect 6637 11595 6703 11598
rect 7741 11595 7807 11598
rect 11145 11658 11211 11661
rect 17769 11658 17835 11661
rect 11145 11656 17835 11658
rect 11145 11600 11150 11656
rect 11206 11600 17774 11656
rect 17830 11600 17835 11656
rect 11145 11598 17835 11600
rect 11145 11595 11211 11598
rect 17769 11595 17835 11598
rect 13537 11522 13603 11525
rect 14549 11522 14615 11525
rect 13537 11520 14615 11522
rect 13537 11464 13542 11520
rect 13598 11464 14554 11520
rect 14610 11464 14615 11520
rect 13537 11462 14615 11464
rect 13537 11459 13603 11462
rect 14549 11459 14615 11462
rect 13537 11250 13603 11253
rect 15285 11250 15351 11253
rect 13537 11248 15351 11250
rect 13537 11192 13542 11248
rect 13598 11192 15290 11248
rect 15346 11192 15351 11248
rect 13537 11190 15351 11192
rect 13537 11187 13603 11190
rect 15285 11187 15351 11190
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 9581 10978 9647 10981
rect 11053 10978 11119 10981
rect 9581 10976 11119 10978
rect 9581 10920 9586 10976
rect 9642 10920 11058 10976
rect 11114 10920 11119 10976
rect 9581 10918 11119 10920
rect 9581 10915 9647 10918
rect 11053 10915 11119 10918
rect 18413 10978 18479 10981
rect 19200 10978 20000 11008
rect 18413 10976 20000 10978
rect 18413 10920 18418 10976
rect 18474 10920 20000 10976
rect 18413 10918 20000 10920
rect 18413 10915 18479 10918
rect 19200 10888 20000 10918
rect 10961 10570 11027 10573
rect 14457 10570 14523 10573
rect 10961 10568 14523 10570
rect 10961 10512 10966 10568
rect 11022 10512 14462 10568
rect 14518 10512 14523 10568
rect 10961 10510 14523 10512
rect 10961 10507 11027 10510
rect 14457 10507 14523 10510
rect 13077 10434 13143 10437
rect 15193 10434 15259 10437
rect 13077 10432 15259 10434
rect 13077 10376 13082 10432
rect 13138 10376 15198 10432
rect 15254 10376 15259 10432
rect 13077 10374 15259 10376
rect 13077 10371 13143 10374
rect 15193 10371 15259 10374
rect 6821 10298 6887 10301
rect 11881 10298 11947 10301
rect 6821 10296 11947 10298
rect 6821 10240 6826 10296
rect 6882 10240 11886 10296
rect 11942 10240 11947 10296
rect 6821 10238 11947 10240
rect 6821 10235 6887 10238
rect 11881 10235 11947 10238
rect 0 10162 800 10192
rect 1301 10162 1367 10165
rect 0 10160 1367 10162
rect 0 10104 1306 10160
rect 1362 10104 1367 10160
rect 0 10102 1367 10104
rect 0 10072 800 10102
rect 1301 10099 1367 10102
rect 9397 10162 9463 10165
rect 12801 10162 12867 10165
rect 9397 10160 12867 10162
rect 9397 10104 9402 10160
rect 9458 10104 12806 10160
rect 12862 10104 12867 10160
rect 9397 10102 12867 10104
rect 9397 10099 9463 10102
rect 12801 10099 12867 10102
rect 8109 10026 8175 10029
rect 9581 10026 9647 10029
rect 13445 10026 13511 10029
rect 8109 10024 13511 10026
rect 8109 9968 8114 10024
rect 8170 9968 9586 10024
rect 9642 9968 13450 10024
rect 13506 9968 13511 10024
rect 8109 9966 13511 9968
rect 8109 9963 8175 9966
rect 9581 9963 9647 9966
rect 13445 9963 13511 9966
rect 3417 9618 3483 9621
rect 4061 9618 4127 9621
rect 5257 9618 5323 9621
rect 3417 9616 5323 9618
rect 3417 9560 3422 9616
rect 3478 9560 4066 9616
rect 4122 9560 5262 9616
rect 5318 9560 5323 9616
rect 3417 9558 5323 9560
rect 3417 9555 3483 9558
rect 4061 9555 4127 9558
rect 5257 9555 5323 9558
rect 9765 9482 9831 9485
rect 11881 9482 11947 9485
rect 9765 9480 11947 9482
rect 9765 9424 9770 9480
rect 9826 9424 11886 9480
rect 11942 9424 11947 9480
rect 9765 9422 11947 9424
rect 9765 9419 9831 9422
rect 11881 9419 11947 9422
rect 0 9346 800 9376
rect 1209 9346 1275 9349
rect 0 9344 1275 9346
rect 0 9288 1214 9344
rect 1270 9288 1275 9344
rect 0 9286 1275 9288
rect 0 9256 800 9286
rect 1209 9283 1275 9286
rect 12617 8938 12683 8941
rect 15929 8938 15995 8941
rect 12617 8936 15995 8938
rect 12617 8880 12622 8936
rect 12678 8880 15934 8936
rect 15990 8880 15995 8936
rect 12617 8878 15995 8880
rect 12617 8875 12683 8878
rect 15929 8875 15995 8878
rect 1117 8666 1183 8669
rect 798 8664 1183 8666
rect 798 8608 1122 8664
rect 1178 8608 1183 8664
rect 798 8606 1183 8608
rect 798 8560 858 8606
rect 1117 8603 1183 8606
rect 15837 8666 15903 8669
rect 15837 8664 19074 8666
rect 15837 8608 15842 8664
rect 15898 8608 19074 8664
rect 15837 8606 19074 8608
rect 15837 8603 15903 8606
rect 0 8470 858 8560
rect 19014 8530 19074 8606
rect 19200 8530 20000 8560
rect 1056 8518 18908 8530
rect 0 8440 800 8470
rect 1056 8462 8220 8518
rect 8276 8462 8300 8518
rect 8356 8462 8380 8518
rect 8436 8462 8460 8518
rect 8516 8462 16220 8518
rect 16276 8462 16300 8518
rect 16356 8462 16380 8518
rect 16436 8462 16460 8518
rect 16516 8462 18908 8518
rect 19014 8470 20000 8530
rect 1056 8438 18908 8462
rect 19200 8440 20000 8470
rect 1056 8382 8220 8438
rect 8276 8382 8300 8438
rect 8356 8382 8380 8438
rect 8436 8382 8460 8438
rect 8516 8382 16220 8438
rect 16276 8382 16300 8438
rect 16356 8382 16380 8438
rect 16436 8382 16460 8438
rect 16516 8382 18908 8438
rect 1056 8358 18908 8382
rect 1056 8302 8220 8358
rect 8276 8302 8300 8358
rect 8356 8302 8380 8358
rect 8436 8302 8460 8358
rect 8516 8302 16220 8358
rect 16276 8302 16300 8358
rect 16356 8302 16380 8358
rect 16436 8302 16460 8358
rect 16516 8302 18908 8358
rect 1056 8278 18908 8302
rect 1056 8222 8220 8278
rect 8276 8222 8300 8278
rect 8356 8222 8380 8278
rect 8436 8222 8460 8278
rect 8516 8222 16220 8278
rect 16276 8222 16300 8278
rect 16356 8222 16380 8278
rect 16436 8222 16460 8278
rect 16516 8222 18908 8278
rect 1056 8210 18908 8222
rect 0 7714 800 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 800 7654
rect 4061 7651 4127 7654
rect 0 6898 800 6928
rect 3877 6898 3943 6901
rect 0 6896 3943 6898
rect 0 6840 3882 6896
rect 3938 6840 3943 6896
rect 0 6838 3943 6840
rect 0 6808 800 6838
rect 3877 6835 3943 6838
rect 10869 6218 10935 6221
rect 12985 6218 13051 6221
rect 10869 6216 13051 6218
rect 10869 6160 10874 6216
rect 10930 6160 12990 6216
rect 13046 6160 13051 6216
rect 10869 6158 13051 6160
rect 10869 6155 10935 6158
rect 12985 6155 13051 6158
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 17861 6082 17927 6085
rect 19200 6082 20000 6112
rect 17861 6080 20000 6082
rect 17861 6024 17866 6080
rect 17922 6024 20000 6080
rect 17861 6022 20000 6024
rect 17861 6019 17927 6022
rect 19200 5992 20000 6022
rect 0 5266 800 5296
rect 1117 5266 1183 5269
rect 0 5264 1183 5266
rect 0 5208 1122 5264
rect 1178 5208 1183 5264
rect 0 5206 1183 5208
rect 0 5176 800 5206
rect 1117 5203 1183 5206
rect 1056 4518 18908 4530
rect 0 4450 800 4480
rect 1056 4462 4220 4518
rect 4276 4462 4300 4518
rect 4356 4462 4380 4518
rect 4436 4462 4460 4518
rect 4516 4462 12220 4518
rect 12276 4462 12300 4518
rect 12356 4462 12380 4518
rect 12436 4462 12460 4518
rect 12516 4462 18908 4518
rect 0 4360 858 4450
rect 798 4178 858 4360
rect 1056 4438 18908 4462
rect 1056 4382 4220 4438
rect 4276 4382 4300 4438
rect 4356 4382 4380 4438
rect 4436 4382 4460 4438
rect 4516 4382 12220 4438
rect 12276 4382 12300 4438
rect 12356 4382 12380 4438
rect 12436 4382 12460 4438
rect 12516 4382 18908 4438
rect 1056 4358 18908 4382
rect 1056 4302 4220 4358
rect 4276 4302 4300 4358
rect 4356 4302 4380 4358
rect 4436 4302 4460 4358
rect 4516 4302 12220 4358
rect 12276 4302 12300 4358
rect 12356 4302 12380 4358
rect 12436 4302 12460 4358
rect 12516 4302 18908 4358
rect 1056 4278 18908 4302
rect 1056 4222 4220 4278
rect 4276 4222 4300 4278
rect 4356 4222 4380 4278
rect 4436 4222 4460 4278
rect 4516 4222 12220 4278
rect 12276 4222 12300 4278
rect 12356 4222 12380 4278
rect 12436 4222 12460 4278
rect 12516 4222 18908 4278
rect 1056 4210 18908 4222
rect 933 4178 999 4181
rect 798 4176 999 4178
rect 798 4120 938 4176
rect 994 4120 999 4176
rect 798 4118 999 4120
rect 933 4115 999 4118
rect 0 3634 800 3664
rect 3049 3634 3115 3637
rect 0 3632 3115 3634
rect 0 3576 3054 3632
rect 3110 3576 3115 3632
rect 0 3574 3115 3576
rect 0 3544 800 3574
rect 3049 3571 3115 3574
rect 15469 3634 15535 3637
rect 19200 3634 20000 3664
rect 15469 3632 20000 3634
rect 15469 3576 15474 3632
rect 15530 3576 20000 3632
rect 15469 3574 20000 3576
rect 15469 3571 15535 3574
rect 19200 3544 20000 3574
rect 0 2818 800 2848
rect 2865 2818 2931 2821
rect 0 2816 2931 2818
rect 0 2760 2870 2816
rect 2926 2760 2931 2816
rect 0 2758 2931 2760
rect 0 2728 800 2758
rect 2865 2755 2931 2758
rect 0 2002 800 2032
rect 2957 2002 3023 2005
rect 0 2000 3023 2002
rect 0 1944 2962 2000
rect 3018 1944 3023 2000
rect 0 1942 3023 1944
rect 0 1912 800 1942
rect 2957 1939 3023 1942
rect 0 1186 800 1216
rect 3325 1186 3391 1189
rect 0 1184 3391 1186
rect 0 1128 3330 1184
rect 3386 1128 3391 1184
rect 0 1126 3391 1128
rect 0 1096 800 1126
rect 3325 1123 3391 1126
rect 15837 1186 15903 1189
rect 19200 1186 20000 1216
rect 15837 1184 20000 1186
rect 15837 1128 15842 1184
rect 15898 1128 20000 1184
rect 15837 1126 20000 1128
rect 15837 1123 15903 1126
rect 19200 1096 20000 1126
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count0_reg_0__RESET_B
timestamp 28801
transform 1 0 9568 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count0_reg_1__RESET_B
timestamp 28801
transform 1 0 9016 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count0_reg_2__RESET_B
timestamp 28801
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count0_reg_3__RESET_B
timestamp 28801
transform 1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count0_reg_4__RESET_B
timestamp 28801
transform 1 0 9016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count1_reg_0__RESET_B
timestamp 28801
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count1_reg_1__RESET_B
timestamp 28801
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count1_reg_2__RESET_B
timestamp 28801
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count1_reg_3__RESET_B
timestamp 28801
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_count1_reg_4__RESET_B
timestamp 28801
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_oscbuf_reg_0__D
timestamp 28801
transform -1 0 15916 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_oscbuf_reg_2__RESET_B
timestamp 28801
transform 1 0 13708 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_prep_reg_1__RESET_B
timestamp 28801
transform 1 0 11592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_prep_reg_2__RESET_B
timestamp 28801
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_tval_reg_0__RESET_B
timestamp 28801
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_tval_reg_1__RESET_B
timestamp 28801
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dll_control_tval_reg_2__RESET_B
timestamp 28801
transform 1 0 11592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U118_A1
timestamp 28801
transform -1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U119_B
timestamp 28801
transform -1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U127_A
timestamp 28801
transform -1 0 8280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U128_A
timestamp 28801
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U128_B
timestamp 28801
transform -1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U129_A
timestamp 28801
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U132_A
timestamp 28801
transform -1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U156_A
timestamp 28801
transform -1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U158_A1_N
timestamp 28801
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U158_A2_N
timestamp 28801
transform -1 0 16468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U162_A
timestamp 28801
transform -1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U163_S
timestamp 28801
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U165_A1_N
timestamp 28801
transform 1 0 11592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U165_A2_N
timestamp 28801
transform -1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U167_A
timestamp 28801
transform -1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U170_A
timestamp 28801
transform -1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U174_A
timestamp 28801
transform -1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U215_A
timestamp 28801
transform -1 0 2392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U216_A
timestamp 28801
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U217_A
timestamp 28801
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U219_A
timestamp 28801
transform -1 0 2852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U225_A
timestamp 28801
transform -1 0 4876 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U319_B
timestamp 28801
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U321_B
timestamp 28801
transform -1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U322_A
timestamp 28801
transform -1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U326_B
timestamp 28801
transform -1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U330_B
timestamp 28801
transform -1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U334_A
timestamp 28801
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U334_B
timestamp 28801
transform -1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U336_A
timestamp 28801
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U336_B
timestamp 28801
transform -1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U338_A
timestamp 28801
transform -1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U338_B
timestamp 28801
transform -1 0 2024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U339_A
timestamp 28801
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U339_B
timestamp 28801
transform 1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U340_B
timestamp 28801
transform -1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U343_A2
timestamp 28801
transform -1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U346_A1
timestamp 28801
transform 1 0 16284 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U346_S
timestamp 28801
transform -1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U347_A1
timestamp 28801
transform -1 0 2668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U347_S
timestamp 28801
transform 1 0 2392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U348_A1
timestamp 28801
transform -1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U348_S
timestamp 28801
transform -1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U355_A1
timestamp 28801
transform -1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U356_A
timestamp 28801
transform -1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_U356_B
timestamp 28801
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_count0_reg_0_
timestamp 28801
transform 1 0 7268 0 -1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  dll_control_count0_reg_1_
timestamp 28801
transform -1 0 8464 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  dll_control_count0_reg_2_
timestamp 28801
transform 1 0 6716 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  dll_control_count0_reg_3_
timestamp 28801
transform 1 0 7360 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count0_reg_4_
timestamp 28801
transform 1 0 6624 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count1_reg_0_
timestamp 28801
transform -1 0 3496 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count1_reg_1_
timestamp 28801
transform -1 0 6164 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count1_reg_2_
timestamp 28801
transform 1 0 1472 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count1_reg_3_
timestamp 28801
transform 1 0 1472 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_count1_reg_4_
timestamp 28801
transform 1 0 2852 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_oscbuf_reg_0_
timestamp 28801
transform -1 0 15548 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_oscbuf_reg_1_
timestamp 28801
transform 1 0 14168 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_oscbuf_reg_2_
timestamp 28801
transform 1 0 14352 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_prep_reg_0_
timestamp 28801
transform 1 0 9384 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_prep_reg_1_
timestamp 28801
transform -1 0 13524 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_prep_reg_2_
timestamp 28801
transform -1 0 13892 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  dll_control_tval_reg_0_
timestamp 28801
transform -1 0 11500 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  dll_control_tval_reg_1_
timestamp 28801
transform -1 0 10948 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_tval_reg_2_
timestamp 28801
transform 1 0 12604 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_tval_reg_3_
timestamp 28801
transform 1 0 13340 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_tval_reg_4_
timestamp 28801
transform 1 0 11592 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_tval_reg_5_
timestamp 28801
transform 1 0 13156 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  dll_control_tval_reg_6_
timestamp 28801
transform 1 0 14168 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_4  fanout1
timestamp 28801
transform -1 0 12696 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout2
timestamp 28801
transform 1 0 7820 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3
timestamp 28801
transform 1 0 1380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_10
timestamp 28801
transform 1 0 2024 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15
timestamp 28801
transform 1 0 2484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_19
timestamp 28801
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 28801
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29
timestamp 28801
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_37
timestamp 28801
transform 1 0 4508 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41
timestamp 28801
transform 1 0 4876 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_48
timestamp 28801
transform 1 0 5520 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 28801
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 28801
transform 1 0 6348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_80
timestamp 28801
transform 1 0 8464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 28801
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_88
timestamp 28801
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 28801
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 28801
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_116
timestamp 28801
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_123
timestamp 28801
transform 1 0 12420 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_131
timestamp 28801
transform 1 0 13156 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 28801
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_141
timestamp 28801
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_164
timestamp 28801
transform 1 0 16192 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 28801
transform 1 0 16652 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_177
timestamp 28801
transform 1 0 17388 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_185
timestamp 28801
transform 1 0 18124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 28801
transform 1 0 18492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3
timestamp 28801
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_26
timestamp 28801
transform 1 0 3496 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_31
timestamp 28801
transform 1 0 3956 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 28801
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 28801
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_65
timestamp 28801
transform 1 0 7084 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_90
timestamp 28801
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_94
timestamp 28801
transform 1 0 9752 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_100
timestamp 28801
transform 1 0 10304 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 28801
transform 1 0 11132 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 28801
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_135
timestamp 28801
transform 1 0 13524 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_157
timestamp 28801
transform 1 0 15548 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 28801
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 28801
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 28801
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_183
timestamp 28801
transform 1 0 17940 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 28801
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 28801
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_12
timestamp 28801
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_21
timestamp 28801
transform 1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 28801
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_29
timestamp 28801
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_39
timestamp 28801
transform 1 0 4692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_63
timestamp 28801
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_67
timestamp 28801
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_71
timestamp 28801
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_80
timestamp 28801
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 28801
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_89
timestamp 28801
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_94
timestamp 28801
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_99
timestamp 28801
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_106
timestamp 28801
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_113
timestamp 28801
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_117
timestamp 28801
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 28801
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 28801
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_162
timestamp 28801
transform 1 0 16008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_170
timestamp 28801
transform 1 0 16744 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_178
timestamp 28801
transform 1 0 17480 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_186
timestamp 28801
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 28801
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 28801
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_15
timestamp 28801
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_26
timestamp 28801
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_33
timestamp 28801
transform 1 0 4140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_39
timestamp 28801
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_44
timestamp 28801
transform 1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_49
timestamp 28801
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 28801
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 28801
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_61
timestamp 28801
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 28801
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_69
timestamp 28801
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_81
timestamp 28801
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_85
timestamp 28801
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_91
timestamp 28801
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_95
timestamp 28801
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_99
timestamp 28801
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp 28801
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 28801
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 28801
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_116
timestamp 28801
transform 1 0 11776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_121
timestamp 28801
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_148
timestamp 28801
transform 1 0 14720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_157
timestamp 28801
transform 1 0 15548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 28801
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_169
timestamp 28801
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_177
timestamp 28801
transform 1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_185
timestamp 28801
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 28801
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 28801
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_10
timestamp 28801
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_14
timestamp 28801
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_20
timestamp 28801
transform 1 0 2944 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 28801
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 28801
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_36
timestamp 28801
transform 1 0 4416 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_44
timestamp 28801
transform 1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 28801
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 28801
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 28801
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_91
timestamp 28801
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_113
timestamp 28801
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_118
timestamp 28801
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_126
timestamp 28801
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_132
timestamp 28801
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 28801
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_141
timestamp 28801
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_147
timestamp 28801
transform 1 0 14628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_162
timestamp 28801
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_169
timestamp 28801
transform 1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_174
timestamp 28801
transform 1 0 17112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_182
timestamp 28801
transform 1 0 17848 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 28801
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_24
timestamp 28801
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_43
timestamp 28801
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 28801
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 28801
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 28801
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_63
timestamp 28801
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_74
timestamp 28801
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_86
timestamp 28801
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_90
timestamp 28801
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_98
timestamp 28801
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_106
timestamp 28801
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 28801
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 28801
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_124
timestamp 28801
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_131
timestamp 28801
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_136
timestamp 28801
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_140
timestamp 28801
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_144
timestamp 28801
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_149
timestamp 28801
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_155
timestamp 28801
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_160
timestamp 28801
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 28801
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_173
timestamp 28801
transform 1 0 17020 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_181
timestamp 28801
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 28801
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 28801
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_7
timestamp 28801
transform 1 0 1748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_15
timestamp 28801
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_19
timestamp 28801
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 28801
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 28801
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_37
timestamp 28801
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_45
timestamp 28801
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_52
timestamp 28801
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_57
timestamp 28801
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_61
timestamp 28801
transform 1 0 6716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_69
timestamp 28801
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_73
timestamp 28801
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_77
timestamp 28801
transform 1 0 8188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 28801
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 28801
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_107
timestamp 28801
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_112
timestamp 28801
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_121
timestamp 28801
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_129
timestamp 28801
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 28801
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 28801
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_147
timestamp 28801
transform 1 0 14628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_152
timestamp 28801
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_156
timestamp 28801
transform 1 0 15456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_160
timestamp 28801
transform 1 0 15824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_168
timestamp 28801
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_172
timestamp 28801
transform 1 0 16928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_180
timestamp 28801
transform 1 0 17664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_185
timestamp 28801
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_189
timestamp 28801
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 28801
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_10
timestamp 28801
transform 1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_14
timestamp 28801
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_18
timestamp 28801
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_22
timestamp 28801
transform 1 0 3128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_30
timestamp 28801
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_34
timestamp 28801
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_38
timestamp 28801
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_42
timestamp 28801
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_49
timestamp 28801
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 28801
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 28801
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_66
timestamp 28801
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_89
timestamp 28801
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_95
timestamp 28801
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_101
timestamp 28801
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_105
timestamp 28801
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 28801
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 28801
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_118
timestamp 28801
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_122
timestamp 28801
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_126
timestamp 28801
transform 1 0 12696 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_132
timestamp 28801
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_156
timestamp 28801
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 28801
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 28801
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_173
timestamp 28801
transform 1 0 17020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_180
timestamp 28801
transform 1 0 17664 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_188
timestamp 28801
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_3
timestamp 28801
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_9
timestamp 28801
transform 1 0 1932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 28801
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 28801
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_35
timestamp 28801
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_46
timestamp 28801
transform 1 0 5336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_54
timestamp 28801
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_61
timestamp 28801
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_66
timestamp 28801
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_74
timestamp 28801
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 28801
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 28801
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 28801
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_89
timestamp 28801
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_96
timestamp 28801
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_102
timestamp 28801
transform 1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_110
timestamp 28801
transform 1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_118
timestamp 28801
transform 1 0 11960 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_124
timestamp 28801
transform 1 0 12512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_128
timestamp 28801
transform 1 0 12880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 28801
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 28801
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp 28801
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_149
timestamp 28801
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_153
timestamp 28801
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_157
timestamp 28801
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_164
timestamp 28801
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_171
timestamp 28801
transform 1 0 16836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_179
timestamp 28801
transform 1 0 17572 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_187
timestamp 28801
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 28801
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_24
timestamp 28801
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_28
timestamp 28801
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_46
timestamp 28801
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 28801
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 28801
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_61
timestamp 28801
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 28801
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_70
timestamp 28801
transform 1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 28801
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_91
timestamp 28801
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_95
timestamp 28801
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_102
timestamp 28801
transform 1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 28801
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 28801
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 28801
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_145
timestamp 28801
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_150
timestamp 28801
transform 1 0 14904 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_157
timestamp 28801
transform 1 0 15548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 28801
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 28801
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_181
timestamp 28801
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_186
timestamp 28801
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 28801
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 28801
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_12
timestamp 28801
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 28801
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 28801
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_34
timestamp 28801
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_39
timestamp 28801
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_44
timestamp 28801
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_48
timestamp 28801
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_52
timestamp 28801
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_57
timestamp 28801
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 28801
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 28801
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_88
timestamp 28801
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_95
timestamp 28801
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_103
timestamp 28801
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_108
timestamp 28801
transform 1 0 11040 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_119
timestamp 28801
transform 1 0 12052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_128
timestamp 28801
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 28801
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_141
timestamp 28801
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_147
timestamp 28801
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_153
timestamp 28801
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_158
timestamp 28801
transform 1 0 15640 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_166
timestamp 28801
transform 1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_173
timestamp 28801
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_188
timestamp 28801
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 28801
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_17
timestamp 28801
transform 1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_39
timestamp 28801
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_43
timestamp 28801
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_47
timestamp 28801
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_51
timestamp 28801
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 28801
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 28801
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_62
timestamp 28801
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_69
timestamp 28801
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_89
timestamp 28801
transform 1 0 9292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_97
timestamp 28801
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_101
timestamp 28801
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 28801
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 28801
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_117
timestamp 28801
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_121
timestamp 28801
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_128
timestamp 28801
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_154
timestamp 28801
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_159
timestamp 28801
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_164
timestamp 28801
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 28801
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_173
timestamp 28801
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_180
timestamp 28801
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_187
timestamp 28801
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 28801
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_7
timestamp 28801
transform 1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_11
timestamp 28801
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_15
timestamp 28801
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_19
timestamp 28801
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 28801
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 28801
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 28801
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_36
timestamp 28801
transform 1 0 4416 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_55
timestamp 28801
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_62
timestamp 28801
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_73
timestamp 28801
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 28801
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_85
timestamp 28801
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_89
timestamp 28801
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_93
timestamp 28801
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp 28801
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 28801
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_106
timestamp 28801
transform 1 0 10856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_117
timestamp 28801
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_124
timestamp 28801
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_129
timestamp 28801
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 28801
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 28801
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_165
timestamp 28801
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_170
timestamp 28801
transform 1 0 16744 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_174
timestamp 28801
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_183
timestamp 28801
transform 1 0 17940 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_188
timestamp 28801
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 28801
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_10
timestamp 28801
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_19
timestamp 28801
transform 1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_24
timestamp 28801
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_34
timestamp 28801
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_40
timestamp 28801
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_48
timestamp 28801
transform 1 0 5520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 28801
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 28801
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 28801
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_71
timestamp 28801
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_76
timestamp 28801
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_87
timestamp 28801
transform 1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 28801
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 28801
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 28801
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_116
timestamp 28801
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_122
timestamp 28801
transform 1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_126
timestamp 28801
transform 1 0 12696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_132
timestamp 28801
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_139
timestamp 28801
transform 1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_149
timestamp 28801
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_154
timestamp 28801
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_158
timestamp 28801
transform 1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 28801
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 28801
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_183
timestamp 28801
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_188
timestamp 28801
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 28801
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 28801
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 28801
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_41
timestamp 28801
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_62
timestamp 28801
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_67
timestamp 28801
transform 1 0 7268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_76
timestamp 28801
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 28801
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 28801
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_95
timestamp 28801
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_101
timestamp 28801
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_105
timestamp 28801
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_112
timestamp 28801
transform 1 0 11408 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_116
timestamp 28801
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_124
timestamp 28801
transform 1 0 12512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_129
timestamp 28801
transform 1 0 12972 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 28801
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 28801
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_145
timestamp 28801
transform 1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_150
timestamp 28801
transform 1 0 14904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_154
timestamp 28801
transform 1 0 15272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_158
timestamp 28801
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_163
timestamp 28801
transform 1 0 16100 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_184
timestamp 28801
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_189
timestamp 28801
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 28801
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_13
timestamp 28801
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_18
timestamp 28801
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_26
timestamp 28801
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_36
timestamp 28801
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_41
timestamp 28801
transform 1 0 4876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_46
timestamp 28801
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_50
timestamp 28801
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 28801
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 28801
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_69
timestamp 28801
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_78
timestamp 28801
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_89
timestamp 28801
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_93
timestamp 28801
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_98
timestamp 28801
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 28801
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 28801
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_116
timestamp 28801
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_127
timestamp 28801
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_136
timestamp 28801
transform 1 0 13616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_149
timestamp 28801
transform 1 0 14812 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_154
timestamp 28801
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_159
timestamp 28801
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 28801
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 28801
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_177
timestamp 28801
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_186
timestamp 28801
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 28801
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_7
timestamp 28801
transform 1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 28801
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 28801
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_41
timestamp 28801
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_45
timestamp 28801
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_50
timestamp 28801
transform 1 0 5704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_54
timestamp 28801
transform 1 0 6072 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_62
timestamp 28801
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_66
timestamp 28801
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_71
timestamp 28801
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_78
timestamp 28801
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 28801
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 28801
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_91
timestamp 28801
transform 1 0 9476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_97
timestamp 28801
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_101
timestamp 28801
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_108
timestamp 28801
transform 1 0 11040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_113
timestamp 28801
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_120
timestamp 28801
transform 1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_126
timestamp 28801
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_130
timestamp 28801
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_134
timestamp 28801
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 28801
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 28801
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_146
timestamp 28801
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_152
timestamp 28801
transform 1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_163
timestamp 28801
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_176
timestamp 28801
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_180
timestamp 28801
transform 1 0 17664 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_185
timestamp 28801
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_189
timestamp 28801
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_3
timestamp 28801
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_7
timestamp 28801
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_14
timestamp 28801
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_25
timestamp 28801
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_29
timestamp 28801
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_36
timestamp 28801
transform 1 0 4416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_42
timestamp 28801
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 28801
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 28801
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_65
timestamp 28801
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_69
timestamp 28801
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_74
timestamp 28801
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_78
timestamp 28801
transform 1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_86
timestamp 28801
transform 1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_91
timestamp 28801
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_99
timestamp 28801
transform 1 0 10212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_107
timestamp 28801
transform 1 0 10948 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 28801
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 28801
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_122
timestamp 28801
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_133
timestamp 28801
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_138
timestamp 28801
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_142
timestamp 28801
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_148
timestamp 28801
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_152
timestamp 28801
transform 1 0 15088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_158
timestamp 28801
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_163
timestamp 28801
transform 1 0 16100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 28801
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 28801
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_188
timestamp 28801
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 28801
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_9
timestamp 28801
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_20
timestamp 28801
transform 1 0 2944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 28801
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 28801
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_33
timestamp 28801
transform 1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_53
timestamp 28801
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_57
timestamp 28801
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_62
timestamp 28801
transform 1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_69
timestamp 28801
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_76
timestamp 28801
transform 1 0 8096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 28801
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 28801
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_92
timestamp 28801
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_99
timestamp 28801
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 28801
transform 1 0 10856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 28801
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_120
timestamp 28801
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_125
timestamp 28801
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_129
timestamp 28801
transform 1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 28801
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 28801
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_150
timestamp 28801
transform 1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_159
timestamp 28801
transform 1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_165
timestamp 28801
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_174
timestamp 28801
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_183
timestamp 28801
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 28801
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 28801
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_12
timestamp 28801
transform 1 0 2208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_32
timestamp 28801
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_37
timestamp 28801
transform 1 0 4508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_41
timestamp 28801
transform 1 0 4876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_49
timestamp 28801
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 28801
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 28801
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_62
timestamp 28801
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_66
timestamp 28801
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_71
timestamp 28801
transform 1 0 7636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_80
timestamp 28801
transform 1 0 8464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_87
timestamp 28801
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_92
timestamp 28801
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_101
timestamp 28801
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_106
timestamp 28801
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 28801
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 28801
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_123
timestamp 28801
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_127
timestamp 28801
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_132
timestamp 28801
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_138
timestamp 28801
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_143
timestamp 28801
transform 1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_148
timestamp 28801
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_161
timestamp 28801
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 28801
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 28801
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 28801
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 28801
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_9
timestamp 28801
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_13
timestamp 28801
transform 1 0 2300 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_16
timestamp 28801
transform 1 0 2576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_21
timestamp 28801
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 28801
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 28801
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_34
timestamp 28801
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_45
timestamp 28801
transform 1 0 5244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_59
timestamp 28801
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_68
timestamp 28801
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 28801
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 28801
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_90
timestamp 28801
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_103
timestamp 28801
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_108
timestamp 28801
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_117
timestamp 28801
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_127
timestamp 28801
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 28801
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 28801
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_145
timestamp 28801
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_154
timestamp 28801
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_158
timestamp 28801
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_177
timestamp 28801
transform 1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_186
timestamp 28801
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 28801
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_7
timestamp 28801
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 28801
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_16
timestamp 28801
transform 1 0 2576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_29
timestamp 28801
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_35
timestamp 28801
transform 1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 28801
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 28801
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_61
timestamp 28801
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_66
timestamp 28801
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_86
timestamp 28801
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_91
timestamp 28801
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 28801
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 28801
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_116
timestamp 28801
transform 1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_129
timestamp 28801
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_141
timestamp 28801
transform 1 0 14076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_156
timestamp 28801
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 28801
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 28801
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_181
timestamp 28801
transform 1 0 17756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_187
timestamp 28801
transform 1 0 18308 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 28801
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_6
timestamp 28801
transform 1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_10
timestamp 28801
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_14
timestamp 28801
transform 1 0 2392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_17
timestamp 28801
transform 1 0 2668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_21
timestamp 28801
transform 1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 28801
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 28801
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_37
timestamp 28801
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_41
timestamp 28801
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_49
timestamp 28801
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_54
timestamp 28801
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_57
timestamp 28801
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_61
timestamp 28801
transform 1 0 6716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_67
timestamp 28801
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_72
timestamp 28801
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 28801
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 28801
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_92
timestamp 28801
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_102
timestamp 28801
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_106
timestamp 28801
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_111
timestamp 28801
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_113
timestamp 28801
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_121
timestamp 28801
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_128
timestamp 28801
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_133
timestamp 28801
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 28801
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_141
timestamp 28801
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_147
timestamp 28801
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_153
timestamp 28801
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_158
timestamp 28801
transform 1 0 15640 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_163
timestamp 28801
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_167
timestamp 28801
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_169
timestamp 28801
transform 1 0 16652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_172
timestamp 28801
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_181
timestamp 28801
transform 1 0 17756 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_186
timestamp 28801
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 28801
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 28801
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 28801
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 28801
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 28801
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 28801
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 28801
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 28801
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 28801
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 28801
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 28801
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 28801
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 28801
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 28801
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 28801
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 28801
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 28801
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 28801
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 28801
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 28801
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 28801
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 28801
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 28801
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 28801
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 28801
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 28801
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 28801
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 28801
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 28801
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 28801
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 28801
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 28801
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 28801
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 28801
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 28801
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 28801
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 28801
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 28801
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 28801
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 28801
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 28801
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 28801
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 28801
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 28801
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 28801
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 28801
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_0__id_delaybuf0
timestamp 28801
transform -1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_0__id_delaybuf1
timestamp 28801
transform 1 0 6992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_0__id_delayen0
timestamp 28801
transform -1 0 7084 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_0__id_delayen1
timestamp 28801
transform -1 0 6808 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_0__id_delayenb0
timestamp 28801
transform -1 0 6808 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_0__id_delayenb1
timestamp 28801
transform -1 0 7452 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_0__id_delayint0
timestamp 28801
transform -1 0 6164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_1__id_delaybuf0
timestamp 28801
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_1__id_delaybuf1
timestamp 28801
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_1__id_delayen0
timestamp 28801
transform 1 0 2208 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_1__id_delayen1
timestamp 28801
transform 1 0 3588 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_1__id_delayenb0
timestamp 28801
transform 1 0 1748 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_1__id_delayenb1
timestamp 28801
transform -1 0 4876 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_1__id_delayint0
timestamp 28801
transform -1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_2__id_delaybuf0
timestamp 28801
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_2__id_delaybuf1
timestamp 28801
transform 1 0 5060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_2__id_delayen0
timestamp 28801
transform 1 0 2760 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_2__id_delayen1
timestamp 28801
transform 1 0 3772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_2__id_delayenb0
timestamp 28801
transform 1 0 1932 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_2__id_delayenb1
timestamp 28801
transform -1 0 4876 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_2__id_delayint0
timestamp 28801
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_3__id_delaybuf0
timestamp 28801
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_3__id_delaybuf1
timestamp 28801
transform -1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_3__id_delayen0
timestamp 28801
transform 1 0 4968 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_3__id_delayen1
timestamp 28801
transform -1 0 7084 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_3__id_delayenb0
timestamp 28801
transform 1 0 4324 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_3__id_delayenb1
timestamp 28801
transform -1 0 6164 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_3__id_delayint0
timestamp 28801
transform -1 0 4140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_4__id_delaybuf0
timestamp 28801
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_4__id_delaybuf1
timestamp 28801
transform -1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_4__id_delayen0
timestamp 28801
transform 1 0 4968 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_4__id_delayen1
timestamp 28801
transform -1 0 7360 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_4__id_delayenb0
timestamp 28801
transform 1 0 4508 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_4__id_delayenb1
timestamp 28801
transform -1 0 6532 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_4__id_delayint0
timestamp 28801
transform -1 0 6072 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_5__id_delaybuf0
timestamp 28801
transform -1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_5__id_delaybuf1
timestamp 28801
transform -1 0 3496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_5__id_delayen0
timestamp 28801
transform 1 0 2300 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_5__id_delayen1
timestamp 28801
transform -1 0 4508 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_5__id_delayenb0
timestamp 28801
transform 1 0 2392 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_5__id_delayenb1
timestamp 28801
transform -1 0 3772 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_5__id_delayint0
timestamp 28801
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_6__id_delaybuf0
timestamp 28801
transform 1 0 3864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_6__id_delaybuf1
timestamp 28801
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_6__id_delayen0
timestamp 28801
transform 1 0 7912 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_6__id_delayen1
timestamp 28801
transform 1 0 7820 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_6__id_delayenb0
timestamp 28801
transform 1 0 7360 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_6__id_delayenb1
timestamp 28801
transform 1 0 7636 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_6__id_delayint0
timestamp 28801
transform -1 0 7728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_7__id_delaybuf0
timestamp 28801
transform 1 0 9200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_7__id_delaybuf1
timestamp 28801
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_7__id_delayen0
timestamp 28801
transform 1 0 11592 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_7__id_delayen1
timestamp 28801
transform 1 0 12144 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_7__id_delayenb0
timestamp 28801
transform 1 0 9660 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_7__id_delayenb1
timestamp 28801
transform 1 0 11960 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_7__id_delayint0
timestamp 28801
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_8__id_delaybuf0
timestamp 28801
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_8__id_delaybuf1
timestamp 28801
transform 1 0 15364 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_8__id_delayen0
timestamp 28801
transform 1 0 15640 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_8__id_delayen1
timestamp 28801
transform 1 0 14628 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_8__id_delayenb0
timestamp 28801
transform 1 0 15732 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_8__id_delayenb1
timestamp 28801
transform 1 0 14444 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_8__id_delayint0
timestamp 28801
transform 1 0 15824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_9__id_delaybuf0
timestamp 28801
transform 1 0 17940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_9__id_delaybuf1
timestamp 28801
transform -1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_9__id_delayen0
timestamp 28801
transform 1 0 17112 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_9__id_delayen1
timestamp 28801
transform -1 0 18216 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_9__id_delayenb0
timestamp 28801
transform 1 0 16836 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_9__id_delayenb1
timestamp 28801
transform 1 0 16744 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_9__id_delayint0
timestamp 28801
transform -1 0 11316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_10__id_delaybuf0
timestamp 28801
transform -1 0 18492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_10__id_delaybuf1
timestamp 28801
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_10__id_delayen0
timestamp 28801
transform 1 0 17296 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_10__id_delayen1
timestamp 28801
transform 1 0 16468 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_10__id_delayenb0
timestamp 28801
transform 1 0 16744 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_10__id_delayenb1
timestamp 28801
transform 1 0 16284 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_10__id_delayint0
timestamp 28801
transform 1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc_dstage_11__id_delaybuf0
timestamp 28801
transform -1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_dstage_11__id_delaybuf1
timestamp 28801
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_11__id_delayen0
timestamp 28801
transform 1 0 16744 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_dstage_11__id_delayen1
timestamp 28801
transform 1 0 17572 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_dstage_11__id_delayenb0
timestamp 28801
transform 1 0 16376 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_dstage_11__id_delayenb1
timestamp 28801
transform 1 0 16928 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_dstage_11__id_delayint0
timestamp 28801
transform 1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc_ibufp00
timestamp 28801
transform -1 0 5980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc_ibufp01
timestamp 28801
transform -1 0 6164 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc_ibufp10
timestamp 28801
transform -1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc_ibufp11
timestamp 28801
transform 1 0 1472 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc_iss_const1
timestamp 28801
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc_iss_ctrlen0
timestamp 28801
transform -1 0 8464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc_iss_delaybuf0
timestamp 28801
transform 1 0 11132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc_iss_delayen0
timestamp 28801
transform 1 0 8464 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc_iss_delayen1
timestamp 28801
transform 1 0 10580 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc_iss_delayenb0
timestamp 28801
transform 1 0 7636 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc_iss_delayenb1
timestamp 28801
transform -1 0 10396 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc_iss_delayint0
timestamp 28801
transform -1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc_iss_reseten0
timestamp 28801
transform -1 0 6808 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 28801
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 28801
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 28801
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 28801
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 28801
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 28801
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 28801
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 28801
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 28801
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 28801
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 28801
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 28801
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 28801
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 28801
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 28801
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 28801
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 28801
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 28801
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 28801
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 28801
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 28801
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 28801
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 28801
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 28801
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 28801
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 28801
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 28801
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 28801
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 28801
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 28801
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 28801
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 28801
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 28801
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 28801
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 28801
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 28801
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 28801
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 28801
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 28801
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 28801
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 28801
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 28801
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 28801
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 28801
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 28801
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 28801
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 28801
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 28801
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 28801
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 28801
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 28801
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 28801
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 28801
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 28801
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 28801
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 28801
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 28801
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 28801
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 28801
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 28801
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 28801
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 28801
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 28801
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 28801
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 28801
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 28801
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 28801
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 28801
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 28801
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 28801
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 28801
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 28801
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 28801
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 28801
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 28801
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  U104
timestamp 28801
transform 1 0 6992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  U105
timestamp 28801
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  U106
timestamp 28801
transform 1 0 6992 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  U107
timestamp 28801
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  U108
timestamp 28801
transform -1 0 8096 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  U109
timestamp 28801
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  U110
timestamp 28801
transform 1 0 9752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  U111
timestamp 28801
transform -1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U112
timestamp 28801
transform -1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  U113
timestamp 28801
transform -1 0 13616 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  U114
timestamp 28801
transform -1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  U115
timestamp 28801
transform 1 0 11592 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  U116
timestamp 28801
transform 1 0 11960 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  U117
timestamp 28801
transform 1 0 9016 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  U118
timestamp 28801
transform 1 0 8464 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  U119
timestamp 28801
transform -1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U120
timestamp 28801
transform 1 0 15824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  U121
timestamp 28801
transform 1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  U122
timestamp 28801
transform -1 0 9016 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  U123
timestamp 28801
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U124
timestamp 28801
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  U125
timestamp 28801
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U126
timestamp 28801
transform -1 0 9108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U127
timestamp 28801
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U128
timestamp 28801
transform -1 0 7636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U129
timestamp 28801
transform 1 0 7360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U130
timestamp 28801
transform -1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U131
timestamp 28801
transform -1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U132
timestamp 28801
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U133
timestamp 28801
transform -1 0 8648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U134
timestamp 28801
transform -1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U135
timestamp 28801
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U136
timestamp 28801
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  U137
timestamp 28801
transform 1 0 9752 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  U138
timestamp 28801
transform 1 0 10672 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  U139
timestamp 28801
transform -1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  U140
timestamp 28801
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U141
timestamp 28801
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  U142
timestamp 28801
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  U143
timestamp 28801
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  U144
timestamp 28801
transform 1 0 16744 0 -1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  U145
timestamp 28801
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U146
timestamp 28801
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U147
timestamp 28801
transform -1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  U148
timestamp 28801
transform -1 0 14812 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  U149
timestamp 28801
transform -1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U150
timestamp 28801
transform -1 0 15640 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U151
timestamp 28801
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  U152
timestamp 28801
transform -1 0 12512 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  U153
timestamp 28801
transform -1 0 13248 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  U154
timestamp 28801
transform 1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U155
timestamp 28801
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U156
timestamp 28801
transform -1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U157
timestamp 28801
transform 1 0 13616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  U158
timestamp 28801
transform 1 0 14168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  U159
timestamp 28801
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U160
timestamp 28801
transform -1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U161
timestamp 28801
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U162
timestamp 28801
transform 1 0 14168 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  U163
timestamp 28801
transform 1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  U164
timestamp 28801
transform -1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  U165
timestamp 28801
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  U166
timestamp 28801
transform -1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U167
timestamp 28801
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U168
timestamp 28801
transform -1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  U169
timestamp 28801
transform -1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U170
timestamp 28801
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U171
timestamp 28801
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  U172
timestamp 28801
transform 1 0 11684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U173
timestamp 28801
transform -1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U174
timestamp 28801
transform 1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U175
timestamp 28801
transform 1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U176
timestamp 28801
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U177
timestamp 28801
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U178
timestamp 28801
transform -1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  U179
timestamp 28801
transform -1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U180
timestamp 28801
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U181
timestamp 28801
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U182
timestamp 28801
transform -1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U183
timestamp 28801
transform -1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U184
timestamp 28801
transform 1 0 10028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U185
timestamp 28801
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U186
timestamp 28801
transform 1 0 12144 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U187
timestamp 28801
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U188
timestamp 28801
transform 1 0 11132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U189
timestamp 28801
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U190
timestamp 28801
transform -1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  U191
timestamp 28801
transform 1 0 7728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  U192
timestamp 28801
transform 1 0 7820 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  U193
timestamp 28801
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  U194
timestamp 28801
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  U195
timestamp 28801
transform 1 0 6808 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  U196
timestamp 28801
transform -1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U197
timestamp 28801
transform -1 0 6164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  U198
timestamp 28801
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  U199
timestamp 28801
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U200
timestamp 28801
transform -1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U201
timestamp 28801
transform -1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U202
timestamp 28801
transform -1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U203
timestamp 28801
transform -1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U204
timestamp 28801
transform -1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U205
timestamp 28801
transform -1 0 2944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U206
timestamp 28801
transform -1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U207
timestamp 28801
transform -1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U208
timestamp 28801
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U209
timestamp 28801
transform 1 0 5244 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U210
timestamp 28801
transform -1 0 6164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U211
timestamp 28801
transform -1 0 7084 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U212
timestamp 28801
transform 1 0 3680 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U213
timestamp 28801
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U214
timestamp 28801
transform -1 0 4508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U215
timestamp 28801
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U216
timestamp 28801
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U217
timestamp 28801
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  U218
timestamp 28801
transform 1 0 3864 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  U219
timestamp 28801
transform -1 0 2484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  U220
timestamp 28801
transform 1 0 1840 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  U221
timestamp 28801
transform 1 0 2392 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  U222
timestamp 28801
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U223
timestamp 28801
transform -1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  U224
timestamp 28801
transform 1 0 1748 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  U225
timestamp 28801
transform 1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  U226
timestamp 28801
transform 1 0 4048 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U227
timestamp 28801
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U228
timestamp 28801
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fa_1  U229
timestamp 28801
transform -1 0 6900 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  U230
timestamp 28801
transform 1 0 3588 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__xor2_1  U231
timestamp 28801
transform -1 0 5980 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  U232
timestamp 28801
transform -1 0 6900 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  U233
timestamp 28801
transform -1 0 5612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U234
timestamp 28801
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U235
timestamp 28801
transform -1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fa_1  U236
timestamp 28801
transform -1 0 3588 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  U237
timestamp 28801
transform -1 0 5336 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__xor2_1  U238
timestamp 28801
transform 1 0 4692 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  U239
timestamp 28801
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  U240
timestamp 28801
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_2  U241
timestamp 28801
transform 1 0 5520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  U242
timestamp 28801
transform -1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  U243
timestamp 28801
transform -1 0 10856 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U244
timestamp 28801
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U245
timestamp 28801
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U246
timestamp 28801
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  U247
timestamp 28801
transform -1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  U248
timestamp 28801
transform -1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U249
timestamp 28801
transform -1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U250
timestamp 28801
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U251
timestamp 28801
transform -1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U252
timestamp 28801
transform -1 0 6716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U253
timestamp 28801
transform 1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  U254
timestamp 28801
transform 1 0 9016 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  U255
timestamp 28801
transform -1 0 10488 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  U256
timestamp 28801
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  U257
timestamp 28801
transform -1 0 10856 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  U258
timestamp 28801
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  U259
timestamp 28801
transform -1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U260
timestamp 28801
transform -1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U261
timestamp 28801
transform 1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U262
timestamp 28801
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U263
timestamp 28801
transform -1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U264
timestamp 28801
transform -1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U265
timestamp 28801
transform -1 0 15088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U266
timestamp 28801
transform 1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U267
timestamp 28801
transform -1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U268
timestamp 28801
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  U269
timestamp 28801
transform 1 0 11868 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U270
timestamp 28801
transform 1 0 16744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U271
timestamp 28801
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U272
timestamp 28801
transform 1 0 16744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  U273
timestamp 28801
transform 1 0 15732 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U274
timestamp 28801
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U275
timestamp 28801
transform -1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  U276
timestamp 28801
transform -1 0 18400 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U277
timestamp 28801
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U278
timestamp 28801
transform 1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U279
timestamp 28801
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U280
timestamp 28801
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U281
timestamp 28801
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U282
timestamp 28801
transform -1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U283
timestamp 28801
transform -1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  U284
timestamp 28801
transform 1 0 11592 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U285
timestamp 28801
transform -1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U286
timestamp 28801
transform 1 0 11592 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U287
timestamp 28801
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U288
timestamp 28801
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U289
timestamp 28801
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U290
timestamp 28801
transform 1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  U291
timestamp 28801
transform -1 0 16008 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U292
timestamp 28801
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U293
timestamp 28801
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U294
timestamp 28801
transform -1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U295
timestamp 28801
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U296
timestamp 28801
transform 1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  U297
timestamp 28801
transform -1 0 18308 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U298
timestamp 28801
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U299
timestamp 28801
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  U300
timestamp 28801
transform -1 0 16192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U301
timestamp 28801
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U302
timestamp 28801
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U303
timestamp 28801
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U304
timestamp 28801
transform -1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U305
timestamp 28801
transform 1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  U306
timestamp 28801
transform 1 0 15916 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  U307
timestamp 28801
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  U308
timestamp 28801
transform -1 0 17940 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U309
timestamp 28801
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U310
timestamp 28801
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U311
timestamp 28801
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U312
timestamp 28801
transform -1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U313
timestamp 28801
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  U314
timestamp 28801
transform -1 0 17664 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  U315
timestamp 28801
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U316
timestamp 28801
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  U317
timestamp 28801
transform 1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  U318
timestamp 28801
transform -1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U319
timestamp 28801
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U320
timestamp 28801
transform -1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U321
timestamp 28801
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U322
timestamp 28801
transform -1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U323
timestamp 28801
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  U324
timestamp 28801
transform 1 0 10120 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  U325
timestamp 28801
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U326
timestamp 28801
transform -1 0 12604 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U327
timestamp 28801
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U328
timestamp 28801
transform 1 0 14168 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U329
timestamp 28801
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U330
timestamp 28801
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  U331
timestamp 28801
transform -1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  U332
timestamp 28801
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  U333
timestamp 28801
transform -1 0 8280 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  U334
timestamp 28801
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U335
timestamp 28801
transform -1 0 13248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U336
timestamp 28801
transform -1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  U337
timestamp 28801
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U338
timestamp 28801
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U339
timestamp 28801
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U340
timestamp 28801
transform -1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U341
timestamp 28801
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  U342
timestamp 28801
transform 1 0 10488 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  U343
timestamp 28801
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  U344
timestamp 28801
transform -1 0 13892 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  U345
timestamp 28801
transform 1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  U346
timestamp 28801
transform 1 0 13248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  U347
timestamp 28801
transform -1 0 5244 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  U348
timestamp 28801
transform -1 0 2300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  U349
timestamp 28801
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U350
timestamp 28801
transform -1 0 13800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  U351
timestamp 28801
transform -1 0 12512 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  U352
timestamp 28801
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  U353
timestamp 28801
transform 1 0 15272 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  U354
timestamp 28801
transform 1 0 11224 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  U355
timestamp 28801
transform -1 0 15916 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  U356
timestamp 28801
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U357
timestamp 28801
transform 1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  U358
timestamp 28801
transform -1 0 2208 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  U359
timestamp 28801
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  U360
timestamp 28801
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  U361
timestamp 28801
transform 1 0 11684 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  U362
timestamp 28801
transform -1 0 2392 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  U363
timestamp 28801
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
<< labels >>
flabel metal2 s 8208 1040 8528 13648 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 16208 1040 16528 13648 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 1056 8210 18908 8530 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 4208 1040 4528 13648 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 12208 1040 12528 13648 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 1056 4210 18908 4530 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 1056 12210 18908 12530 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 5538 14200 5594 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 7010 14200 7066 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 8482 14200 8538 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 9954 14200 10010 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 11426 14200 11482 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 12898 14200 12954 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 15842 14200 15898 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 17314 14200 17370 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 18786 14200 18842 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 19200 13336 20000 13456 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 19200 8440 20000 8560 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 19200 5992 20000 6112 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 19200 3544 20000 3664 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 19200 1096 20000 1216 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 1122 14200 1178 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 2594 14200 2650 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 4066 14200 4122 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
rlabel metal1 9982 13056 9982 13056 0 VGND
rlabel metal1 9982 13600 9982 13600 0 VPWR
rlabel metal1 3404 1870 3404 1870 0 clockp[0]
rlabel metal3 1832 1972 1832 1972 0 clockp[1]
rlabel metal1 6900 7378 6900 7378 0 creset
rlabel metal1 5612 7922 5612 7922 0 dco
rlabel metal1 2806 1326 2806 1326 0 div[0]
rlabel metal1 1794 1292 1794 1292 0 div[1]
rlabel metal1 1380 3502 1380 3502 0 div[2]
rlabel metal1 1472 5202 1472 5202 0 div[3]
rlabel metal1 1702 5712 1702 5712 0 div[4]
rlabel metal1 2990 2414 2990 2414 0 dll_control_count0[0]
rlabel metal1 6118 1360 6118 1360 0 dll_control_count0[1]
rlabel metal1 4048 3978 4048 3978 0 dll_control_count0[2]
rlabel metal2 2530 5950 2530 5950 0 dll_control_count0[3]
rlabel metal1 5382 7344 5382 7344 0 dll_control_count0[4]
rlabel metal1 2714 2074 2714 2074 0 dll_control_count1[0]
rlabel metal1 5382 1326 5382 1326 0 dll_control_count1[1]
rlabel metal1 3581 4046 3581 4046 0 dll_control_count1[2]
rlabel metal2 3266 5916 3266 5916 0 dll_control_count1[3]
rlabel metal1 4692 7174 4692 7174 0 dll_control_count1[4]
rlabel metal1 14122 2074 14122 2074 0 dll_control_oscbuf[0]
rlabel metal2 16974 2108 16974 2108 0 dll_control_oscbuf[1]
rlabel metal2 16146 1734 16146 1734 0 dll_control_oscbuf[2]
rlabel metal1 10948 1938 10948 1938 0 dll_control_prep[0]
rlabel metal1 11040 2346 11040 2346 0 dll_control_prep[1]
rlabel metal1 11354 2278 11354 2278 0 dll_control_prep[2]
rlabel metal1 14490 10064 14490 10064 0 dll_control_tint[0]
rlabel metal2 13110 9452 13110 9452 0 dll_control_tint[1]
rlabel metal1 13018 8500 13018 8500 0 dll_control_tint[2]
rlabel metal1 11868 10030 11868 10030 0 dll_control_tint[3]
rlabel metal1 16100 7786 16100 7786 0 dll_control_tint[4]
rlabel metal1 10028 5202 10028 5202 0 dll_control_tval[0]
rlabel metal1 11270 5202 11270 5202 0 dll_control_tval[1]
rlabel metal1 4232 6698 4232 6698 0 enable
rlabel metal1 1472 8466 1472 8466 0 ext_trim[0]
rlabel metal1 12696 11118 12696 11118 0 ext_trim[10]
rlabel metal1 6486 12852 6486 12852 0 ext_trim[11]
rlabel metal2 8701 14348 8701 14348 0 ext_trim[12]
rlabel metal2 10127 14348 10127 14348 0 ext_trim[13]
rlabel metal2 11454 13377 11454 13377 0 ext_trim[14]
rlabel metal2 12926 13508 12926 13508 0 ext_trim[15]
rlabel metal1 14766 10982 14766 10982 0 ext_trim[16]
rlabel metal2 15042 12342 15042 12342 0 ext_trim[17]
rlabel metal1 16882 13498 16882 13498 0 ext_trim[18]
rlabel metal1 7590 11764 7590 11764 0 ext_trim[19]
rlabel metal1 1472 9622 1472 9622 0 ext_trim[1]
rlabel metal1 14582 13226 14582 13226 0 ext_trim[20]
rlabel metal2 18446 10591 18446 10591 0 ext_trim[21]
rlabel metal1 15640 11662 15640 11662 0 ext_trim[22]
rlabel metal1 18124 7854 18124 7854 0 ext_trim[23]
rlabel metal1 15456 8942 15456 8942 0 ext_trim[24]
rlabel metal3 17626 1156 17626 1156 0 ext_trim[25]
rlabel metal1 1472 10098 1472 10098 0 ext_trim[2]
rlabel metal1 1702 11152 1702 11152 0 ext_trim[3]
rlabel metal2 2530 12461 2530 12461 0 ext_trim[4]
rlabel metal1 1886 12240 1886 12240 0 ext_trim[5]
rlabel metal1 1288 13362 1288 13362 0 ext_trim[6]
rlabel metal1 6670 9554 6670 9554 0 ext_trim[7]
rlabel metal1 2530 12784 2530 12784 0 ext_trim[8]
rlabel metal1 2714 12614 2714 12614 0 ext_trim[9]
rlabel metal1 6670 7854 6670 7854 0 ireset
rlabel metal1 6762 8976 6762 8976 0 itrim[0]
rlabel metal1 17158 11118 17158 11118 0 itrim[10]
rlabel metal1 16192 8942 16192 8942 0 itrim[11]
rlabel metal1 8142 8466 8142 8466 0 itrim[12]
rlabel metal1 7406 9588 7406 9588 0 itrim[13]
rlabel metal1 5290 8942 5290 8942 0 itrim[14]
rlabel metal1 4830 9962 4830 9962 0 itrim[15]
rlabel metal2 13386 10574 13386 10574 0 itrim[16]
rlabel metal1 7314 12308 7314 12308 0 itrim[17]
rlabel metal1 5658 13362 5658 13362 0 itrim[18]
rlabel metal1 1978 8942 1978 8942 0 itrim[1]
rlabel metal1 12328 13158 12328 13158 0 itrim[20]
rlabel metal1 14628 12818 14628 12818 0 itrim[21]
rlabel metal1 16330 11866 16330 11866 0 itrim[22]
rlabel metal1 16238 10030 16238 10030 0 itrim[23]
rlabel metal1 17066 9554 17066 9554 0 itrim[24]
rlabel metal1 10626 8330 10626 8330 0 itrim[25]
rlabel metal1 2116 10030 2116 10030 0 itrim[2]
rlabel metal1 4370 11152 4370 11152 0 itrim[3]
rlabel metal1 4554 12784 4554 12784 0 itrim[4]
rlabel metal1 2438 11764 2438 11764 0 itrim[5]
rlabel metal1 7682 12818 7682 12818 0 itrim[6]
rlabel metal1 10764 13226 10764 13226 0 itrim[7]
rlabel metal1 15502 12750 15502 12750 0 itrim[8]
rlabel metal1 16744 11730 16744 11730 0 itrim[9]
rlabel metal1 10534 7854 10534 7854 0 n100
rlabel metal1 8510 10030 8510 10030 0 n101
rlabel metal1 9982 11050 9982 11050 0 n102
rlabel metal1 10074 2006 10074 2006 0 n103
rlabel metal1 11776 2482 11776 2482 0 n104
rlabel metal1 11730 1530 11730 1530 0 n105
rlabel metal1 8786 2482 8786 2482 0 n106
rlabel metal1 9108 2618 9108 2618 0 n107
rlabel metal1 7820 3162 7820 3162 0 n108
rlabel metal1 6702 4590 6702 4590 0 n109
rlabel metal1 7452 4794 7452 4794 0 n110
rlabel metal1 8786 3026 8786 3026 0 n111
rlabel metal1 7590 4590 7590 4590 0 n112
rlabel metal1 6716 5270 6716 5270 0 n113
rlabel metal2 7222 6766 7222 6766 0 n114
rlabel metal1 4416 6834 4416 6834 0 n115
rlabel metal1 4416 6766 4416 6766 0 n116
rlabel metal2 2622 6324 2622 6324 0 n117
rlabel metal2 2990 6052 2990 6052 0 n118
rlabel metal1 3082 3570 3082 3570 0 n119
rlabel metal2 2622 3978 2622 3978 0 n120
rlabel metal1 6578 1870 6578 1870 0 n121
rlabel metal1 6141 1462 6141 1462 0 n122
rlabel metal1 3818 1394 3818 1394 0 n123
rlabel metal1 4462 1292 4462 1292 0 n124
rlabel metal2 2438 2652 2438 2652 0 n125
rlabel metal1 3450 3094 3450 3094 0 n126
rlabel metal1 2162 2414 2162 2414 0 n127
rlabel metal1 4278 2482 4278 2482 0 n128
rlabel metal1 4370 2414 4370 2414 0 n129
rlabel metal1 5014 2958 5014 2958 0 n130
rlabel metal1 4830 3060 4830 3060 0 n131
rlabel metal2 1886 1088 1886 1088 0 n132
rlabel metal1 3174 3672 3174 3672 0 n133
rlabel metal1 6808 2618 6808 2618 0 n134
rlabel metal1 6348 3570 6348 3570 0 n135
rlabel metal1 6026 4114 6026 4114 0 n136
rlabel metal1 5290 3162 5290 3162 0 n137
rlabel metal1 3864 4590 3864 4590 0 n138
rlabel metal1 4186 5236 4186 5236 0 n139
rlabel metal1 4830 4658 4830 4658 0 n140
rlabel metal1 5658 3978 5658 3978 0 n141
rlabel metal2 2806 5508 2806 5508 0 n142
rlabel metal2 4094 6086 4094 6086 0 n143
rlabel metal1 4830 5678 4830 5678 0 n144
rlabel metal2 4830 5916 4830 5916 0 n145
rlabel metal1 5980 5338 5980 5338 0 n146
rlabel metal1 5612 4522 5612 4522 0 n147
rlabel metal1 6164 6222 6164 6222 0 n148
rlabel metal1 10442 5066 10442 5066 0 n149
rlabel metal1 10764 6766 10764 6766 0 n150
rlabel metal1 10626 10030 10626 10030 0 n151
rlabel metal1 10074 5678 10074 5678 0 n152
rlabel metal1 4600 2618 4600 2618 0 n153
rlabel metal1 3404 2618 3404 2618 0 n154
rlabel metal1 5474 3570 5474 3570 0 n155
rlabel metal1 5382 2958 5382 2958 0 n156
rlabel metal1 5888 2958 5888 2958 0 n157
rlabel metal1 5842 4658 5842 4658 0 n158
rlabel metal1 6670 5712 6670 5712 0 n159
rlabel metal1 6624 4794 6624 4794 0 n160
rlabel metal1 6854 5882 6854 5882 0 n161
rlabel metal1 6072 6290 6072 6290 0 n162
rlabel metal1 9062 5712 9062 5712 0 n163
rlabel metal1 9200 5882 9200 5882 0 n164
rlabel metal1 9062 6324 9062 6324 0 n165
rlabel metal1 9706 6290 9706 6290 0 n166
rlabel metal2 10166 5984 10166 5984 0 n167
rlabel metal1 11362 7718 11362 7718 0 n168
rlabel metal1 9706 5712 9706 5712 0 n169
rlabel metal2 9890 6188 9890 6188 0 n170
rlabel metal2 10442 2689 10442 2689 0 n171
rlabel metal1 10902 2992 10902 2992 0 n172
rlabel metal1 15548 6970 15548 6970 0 n173
rlabel metal1 16514 4046 16514 4046 0 n174
rlabel metal1 16192 3706 16192 3706 0 n175
rlabel metal1 17756 6426 17756 6426 0 n176
rlabel metal1 18078 6766 18078 6766 0 n177
rlabel metal1 14582 6834 14582 6834 0 n178
rlabel metal1 13938 6834 13938 6834 0 n179
rlabel metal1 12834 6834 12834 6834 0 n180
rlabel metal1 10488 3162 10488 3162 0 n181
rlabel metal1 10856 4114 10856 4114 0 n182
rlabel metal2 12098 4556 12098 4556 0 n183
rlabel metal1 12466 4114 12466 4114 0 n184
rlabel metal1 13386 4080 13386 4080 0 n185
rlabel metal1 13340 4182 13340 4182 0 n186
rlabel metal2 11822 4386 11822 4386 0 n187
rlabel metal1 12650 4590 12650 4590 0 n188
rlabel metal2 12006 4522 12006 4522 0 n189
rlabel metal1 11408 4998 11408 4998 0 n190
rlabel metal1 15686 3026 15686 3026 0 n191
rlabel metal1 14168 4114 14168 4114 0 n192
rlabel metal1 15640 3162 15640 3162 0 n193
rlabel metal1 14582 3536 14582 3536 0 n194
rlabel metal1 13846 3570 13846 3570 0 n195
rlabel metal1 13386 3502 13386 3502 0 n196
rlabel metal1 17710 5202 17710 5202 0 n197
rlabel metal2 17618 5508 17618 5508 0 n198
rlabel metal1 12834 5780 12834 5780 0 n199
rlabel metal1 12328 5746 12328 5746 0 n200
rlabel metal1 16330 7854 16330 7854 0 n201
rlabel metal1 12696 5202 12696 5202 0 n202
rlabel metal1 16790 7412 16790 7412 0 n203
rlabel metal1 16974 7446 16974 7446 0 n204
rlabel metal1 16146 5746 16146 5746 0 n205
rlabel metal1 15732 6630 15732 6630 0 n206
rlabel metal1 16606 5644 16606 5644 0 n207
rlabel metal1 16146 6324 16146 6324 0 n208
rlabel metal1 16514 6222 16514 6222 0 n209
rlabel metal1 16652 6426 16652 6426 0 n210
rlabel metal2 16790 6052 16790 6052 0 n211
rlabel metal2 16698 6324 16698 6324 0 n212
rlabel metal1 17250 6970 17250 6970 0 n213
rlabel metal2 16882 7650 16882 7650 0 n214
rlabel metal1 16330 8058 16330 8058 0 n215
rlabel viali 13570 7926 13570 7926 0 n216
rlabel metal2 14858 10829 14858 10829 0 n217
rlabel metal1 16606 3570 16606 3570 0 n218
rlabel metal1 16928 4114 16928 4114 0 n219
rlabel metal1 17434 3706 17434 3706 0 n220
rlabel metal1 15778 4080 15778 4080 0 n221
rlabel metal1 14904 3978 14904 3978 0 n222
rlabel metal1 15226 4114 15226 4114 0 n223
rlabel metal1 16514 3978 16514 3978 0 n224
rlabel metal1 17434 4624 17434 4624 0 n225
rlabel metal1 14582 4556 14582 4556 0 n226
rlabel metal1 14030 4658 14030 4658 0 n227
rlabel metal1 13294 4794 13294 4794 0 n228
rlabel metal1 14398 6732 14398 6732 0 n229
rlabel metal1 11132 6834 11132 6834 0 n230
rlabel metal1 8740 11118 8740 11118 0 n231
rlabel metal1 8878 10608 8878 10608 0 n232
rlabel metal1 12374 11152 12374 11152 0 n233
rlabel metal1 12880 9146 12880 9146 0 n234
rlabel metal2 13754 8007 13754 8007 0 n235
rlabel metal2 14306 9316 14306 9316 0 n236
rlabel metal1 10442 9962 10442 9962 0 n237
rlabel metal1 9890 10676 9890 10676 0 n238
rlabel metal1 12834 10676 12834 10676 0 n239
rlabel metal1 15640 8942 15640 8942 0 n240
rlabel metal1 9016 2346 9016 2346 0 n241
rlabel metal1 13110 3400 13110 3400 0 n242
rlabel metal1 8004 3026 8004 3026 0 n243
rlabel metal2 5934 7854 5934 7854 0 n244
rlabel metal1 9292 8466 9292 8466 0 n245
rlabel metal1 15916 9554 15916 9554 0 n246
rlabel via1 13662 10013 13662 10013 0 n247
rlabel metal1 15226 11628 15226 11628 0 n248
rlabel metal1 2530 12070 2530 12070 0 n249
rlabel metal1 8878 9078 8878 9078 0 n250
rlabel metal2 13754 8772 13754 8772 0 n251
rlabel metal1 13570 8976 13570 8976 0 n252
rlabel via1 15505 9554 15505 9554 0 n253
rlabel metal1 11822 8874 11822 8874 0 n254
rlabel metal1 18308 8058 18308 8058 0 n255
rlabel metal1 12098 11084 12098 11084 0 n256
rlabel metal1 11316 10778 11316 10778 0 n257
rlabel metal1 11730 11866 11730 11866 0 n258
rlabel metal1 10442 11798 10442 11798 0 n259
rlabel metal1 11270 10064 11270 10064 0 n260
rlabel metal1 13248 13294 13248 13294 0 n261
rlabel metal1 10856 11730 10856 11730 0 n262
rlabel metal2 9844 12410 9844 12410 0 n263
rlabel metal2 10442 12240 10442 12240 0 n264
rlabel metal1 7452 11118 7452 11118 0 n265
rlabel metal1 13570 12818 13570 12818 0 n266
rlabel metal1 9844 9622 9844 9622 0 n267
rlabel metal1 1702 11798 1702 11798 0 n268
rlabel metal1 2162 11628 2162 11628 0 n269
rlabel via2 14582 11509 14582 11509 0 n270
rlabel metal1 13800 11866 13800 11866 0 n271
rlabel metal1 13570 9588 13570 9588 0 n272
rlabel metal2 13110 11968 13110 11968 0 n273
rlabel metal2 12650 9622 12650 9622 0 n274
rlabel metal1 10902 11798 10902 11798 0 n275
rlabel metal1 13478 11220 13478 11220 0 n276
rlabel metal1 14812 10778 14812 10778 0 n277
rlabel metal1 2714 11016 2714 11016 0 n278
rlabel metal1 9246 10506 9246 10506 0 n279
rlabel metal1 12489 10778 12489 10778 0 n280
rlabel metal2 14490 9384 14490 9384 0 n281
rlabel metal1 2484 9690 2484 9690 0 n282
rlabel metal1 10580 8942 10580 8942 0 n283
rlabel metal1 12972 9622 12972 9622 0 n284
rlabel metal1 12742 10030 12742 10030 0 n285
rlabel metal1 9292 10234 9292 10234 0 n286
rlabel metal1 9430 10608 9430 10608 0 n287
rlabel metal1 2024 10642 2024 10642 0 n288
rlabel metal2 13754 10591 13754 10591 0 n289
rlabel metal1 8878 9146 8878 9146 0 n290
rlabel metal1 7866 9554 7866 9554 0 n291
rlabel metal1 7774 6290 7774 6290 0 n292
rlabel metal1 12144 1870 12144 1870 0 n54
rlabel metal1 7636 7854 7636 7854 0 n55
rlabel metal1 9936 1394 9936 1394 0 n56
rlabel metal1 3588 6970 3588 6970 0 n57
rlabel metal1 2208 6630 2208 6630 0 n58
rlabel metal2 1794 3876 1794 3876 0 n59
rlabel metal1 3680 1190 3680 1190 0 n60
rlabel metal1 7774 5882 7774 5882 0 n61
rlabel metal1 7084 3570 7084 3570 0 n62
rlabel metal1 7964 1530 7964 1530 0 n63
rlabel metal1 6985 6970 6985 6970 0 n65
rlabel metal1 13432 6970 13432 6970 0 n66
rlabel metal2 11822 6154 11822 6154 0 n67
rlabel metal1 13570 4794 13570 4794 0 n68
rlabel metal1 12926 3128 12926 3128 0 n69
rlabel metal1 11233 4794 11233 4794 0 n70
rlabel metal1 10948 3570 10948 3570 0 n71
rlabel metal1 14030 7786 14030 7786 0 n72
rlabel metal1 6302 2006 6302 2006 0 n73
rlabel metal1 13570 2312 13570 2312 0 n74
rlabel metal1 7820 11662 7820 11662 0 n76
rlabel metal1 4140 11866 4140 11866 0 n77
rlabel metal1 6808 11118 6808 11118 0 n78
rlabel metal1 7498 12614 7498 12614 0 n79
rlabel metal1 7176 11322 7176 11322 0 n80
rlabel metal1 6578 11662 6578 11662 0 n81
rlabel metal1 7774 10574 7774 10574 0 n82
rlabel metal1 3174 10608 3174 10608 0 n83
rlabel metal1 8602 4794 8602 4794 0 n84
rlabel metal1 9062 11662 9062 11662 0 n85
rlabel metal1 15594 9078 15594 9078 0 n86
rlabel metal1 15272 7378 15272 7378 0 n87
rlabel metal2 8142 5066 8142 5066 0 n88
rlabel metal1 7682 4658 7682 4658 0 n89
rlabel metal1 15088 10574 15088 10574 0 n90
rlabel metal1 6394 12716 6394 12716 0 n91
rlabel via2 9890 11883 9890 11883 0 n92
rlabel metal2 12742 7888 12742 7888 0 n93
rlabel metal1 13662 10778 13662 10778 0 n94
rlabel metal1 1886 8364 1886 8364 0 n95
rlabel metal1 6578 12648 6578 12648 0 n96
rlabel metal1 12742 7820 12742 7820 0 n97
rlabel metal1 12282 10030 12282 10030 0 n98
rlabel metal1 10994 11662 10994 11662 0 n99
rlabel metal1 5934 1292 5934 1292 0 net1
rlabel metal2 2438 5202 2438 5202 0 net2
rlabel metal1 15088 2006 15088 2006 0 osc
rlabel viali 5106 6767 5106 6767 0 resetb
rlabel metal2 5750 8058 5750 8058 0 ringosc_c[0]
rlabel metal2 1978 7174 1978 7174 0 ringosc_c[1]
rlabel metal2 8970 7786 8970 7786 0 ringosc_d[0]
rlabel metal1 18032 11798 18032 11798 0 ringosc_d[10]
rlabel metal1 18216 10710 18216 10710 0 ringosc_d[11]
rlabel metal1 11086 8942 11086 8942 0 ringosc_d[12]
rlabel metal1 4646 8432 4646 8432 0 ringosc_d[1]
rlabel metal2 2714 8670 2714 8670 0 ringosc_d[2]
rlabel metal1 4508 10098 4508 10098 0 ringosc_d[3]
rlabel metal1 5704 11730 5704 11730 0 ringosc_d[4]
rlabel metal1 5474 13192 5474 13192 0 ringosc_d[5]
rlabel metal1 2162 6732 2162 6732 0 ringosc_d[6]
rlabel metal1 8878 13226 8878 13226 0 ringosc_d[7]
rlabel metal1 14950 13362 14950 13362 0 ringosc_d[8]
rlabel metal1 18078 12784 18078 12784 0 ringosc_d[9]
rlabel metal1 6624 9146 6624 9146 0 ringosc_dstage_0__id_d0
rlabel metal1 6210 9690 6210 9690 0 ringosc_dstage_0__id_d1
rlabel metal1 6256 8534 6256 8534 0 ringosc_dstage_0__id_d2
rlabel metal1 7314 8942 7314 8942 0 ringosc_dstage_0__id_ts
rlabel metal1 18032 7514 18032 7514 0 ringosc_dstage_10__id_d0
rlabel metal1 17480 13158 17480 13158 0 ringosc_dstage_10__id_d1
rlabel metal1 17986 13294 17986 13294 0 ringosc_dstage_10__id_d2
rlabel metal2 18262 9010 18262 9010 0 ringosc_dstage_10__id_ts
rlabel metal2 18170 9044 18170 9044 0 ringosc_dstage_11__id_d0
rlabel metal1 18170 8942 18170 8942 0 ringosc_dstage_11__id_d1
rlabel metal1 18630 9146 18630 9146 0 ringosc_dstage_11__id_d2
rlabel metal2 17894 9418 17894 9418 0 ringosc_dstage_11__id_ts
rlabel viali 4646 9675 4646 9675 0 ringosc_dstage_1__id_d0
rlabel metal1 4094 8534 4094 8534 0 ringosc_dstage_1__id_d1
rlabel metal1 2944 8466 2944 8466 0 ringosc_dstage_1__id_d2
rlabel metal1 4646 8330 4646 8330 0 ringosc_dstage_1__id_ts
rlabel metal1 4738 9486 4738 9486 0 ringosc_dstage_2__id_d0
rlabel metal1 4048 10030 4048 10030 0 ringosc_dstage_2__id_d1
rlabel metal2 3358 10880 3358 10880 0 ringosc_dstage_2__id_d2
rlabel metal1 3910 9928 3910 9928 0 ringosc_dstage_2__id_ts
rlabel metal1 5704 10574 5704 10574 0 ringosc_dstage_3__id_d0
rlabel metal2 5382 10812 5382 10812 0 ringosc_dstage_3__id_d1
rlabel metal1 4784 11322 4784 11322 0 ringosc_dstage_3__id_d2
rlabel metal1 5382 10710 5382 10710 0 ringosc_dstage_3__id_ts
rlabel viali 6762 12207 6762 12207 0 ringosc_dstage_4__id_d0
rlabel metal1 5934 12138 5934 12138 0 ringosc_dstage_4__id_d1
rlabel metal1 5704 13226 5704 13226 0 ringosc_dstage_4__id_d2
rlabel metal1 6118 12818 6118 12818 0 ringosc_dstage_4__id_ts
rlabel metal1 3910 13192 3910 13192 0 ringosc_dstage_5__id_d0
rlabel metal1 3542 12886 3542 12886 0 ringosc_dstage_5__id_d1
rlabel metal1 2898 11254 2898 11254 0 ringosc_dstage_5__id_d2
rlabel metal1 4002 12614 4002 12614 0 ringosc_dstage_5__id_ts
rlabel metal1 8832 11798 8832 11798 0 ringosc_dstage_6__id_d0
rlabel metal1 7912 13158 7912 13158 0 ringosc_dstage_6__id_d1
rlabel metal1 8050 13362 8050 13362 0 ringosc_dstage_6__id_d2
rlabel metal1 9154 12818 9154 12818 0 ringosc_dstage_6__id_ts
rlabel metal1 12972 12274 12972 12274 0 ringosc_dstage_7__id_d0
rlabel metal1 12926 12886 12926 12886 0 ringosc_dstage_7__id_d1
rlabel metal1 12696 13226 12696 13226 0 ringosc_dstage_7__id_d2
rlabel metal1 12926 12784 12926 12784 0 ringosc_dstage_7__id_ts
rlabel metal1 15318 12274 15318 12274 0 ringosc_dstage_8__id_d0
rlabel metal1 15180 12886 15180 12886 0 ringosc_dstage_8__id_d1
rlabel metal1 16100 12886 16100 12886 0 ringosc_dstage_8__id_d2
rlabel metal1 15640 12818 15640 12818 0 ringosc_dstage_8__id_ts
rlabel metal1 16100 12138 16100 12138 0 ringosc_dstage_9__id_d0
rlabel metal2 17434 13294 17434 13294 0 ringosc_dstage_9__id_d1
rlabel metal1 16468 13362 16468 13362 0 ringosc_dstage_9__id_d2
rlabel metal2 17802 11679 17802 11679 0 ringosc_dstage_9__id_ts
rlabel metal1 7866 7378 7866 7378 0 ringosc_iss_ctrl0
rlabel metal1 11178 8534 11178 8534 0 ringosc_iss_d0
rlabel metal1 10350 8534 10350 8534 0 ringosc_iss_d1
rlabel metal1 9292 8058 9292 8058 0 ringosc_iss_d2
rlabel metal1 6348 6834 6348 6834 0 ringosc_iss_one
<< properties >>
string FIXED_BBOX 0 0 20000 15000
<< end >>
