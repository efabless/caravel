VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_logo
  CLASS BLOCK ;
  FOREIGN caravan_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 25.000 ;
END caravan_logo
END LIBRARY

