magic
tech sky130A
timestamp 1605459841
<< psubdiff >>
rect 145 1334 199 260000
rect 299 1334 355 260000
rect 145 1197 355 1334
rect 145 1037 531 1197
rect 145 998 652 1037
rect 253 900 652 998
rect 355 797 792 900
rect 453 795 792 797
rect 453 690 900 795
rect 565 652 900 690
rect 565 582 1049 652
rect 663 523 1049 582
rect 663 480 1197 523
rect 775 366 1197 480
rect 862 355 1197 366
rect 862 299 180000 355
rect 862 270 1511 299
rect 985 199 1511 270
rect 985 145 180000 199
<< psubdiffcont >>
rect 199 1334 299 260000
rect 1511 199 180000 299
<< locali >>
rect 199 1214 299 1334
rect 100 100 500 500
rect 1437 199 1511 299
<< metal1 >>
rect 275 325 325 420
rect 180 275 420 325
rect 275 180 325 275
<< end >>
