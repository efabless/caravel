magic
tech sky130A
magscale 1 2
timestamp 1665667071
<< viali >>
rect 3525 13481 3559 13515
rect 7849 13481 7883 13515
rect 9229 13481 9263 13515
rect 9597 13481 9631 13515
rect 2697 13413 2731 13447
rect 7297 13413 7331 13447
rect 3341 13345 3375 13379
rect 5181 13345 5215 13379
rect 6469 13345 6503 13379
rect 7757 13345 7791 13379
rect 10977 13345 11011 13379
rect 12725 13345 12759 13379
rect 10149 13311 10183 13345
rect 2053 13277 2087 13311
rect 2789 13277 2823 13311
rect 3801 13277 3835 13311
rect 3893 13277 3927 13311
rect 4077 13277 4111 13311
rect 4629 13277 4663 13311
rect 5273 13277 5307 13311
rect 6101 13277 6135 13311
rect 6745 13277 6779 13311
rect 7118 13277 7152 13311
rect 8217 13277 8251 13311
rect 8677 13277 8711 13311
rect 9413 13277 9447 13311
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 12081 13277 12115 13311
rect 12173 13277 12207 13311
rect 12817 13277 12851 13311
rect 1501 13209 1535 13243
rect 1593 13209 1627 13243
rect 2145 13209 2179 13243
rect 3249 13209 3283 13243
rect 4261 13209 4295 13243
rect 5089 13209 5123 13243
rect 5733 13209 5767 13243
rect 5825 13209 5859 13243
rect 6377 13209 6411 13243
rect 6929 13209 6963 13243
rect 7021 13209 7055 13243
rect 7573 13209 7607 13243
rect 8769 13209 8803 13243
rect 9965 13209 9999 13243
rect 10425 13209 10459 13243
rect 11069 13209 11103 13243
rect 11529 13209 11563 13243
rect 11621 13209 11655 13243
rect 12633 13209 12667 13243
rect 13277 13209 13311 13243
rect 13369 13209 13403 13243
rect 2237 13141 2271 13175
rect 2513 13141 2547 13175
rect 4445 13141 4479 13175
rect 5917 13141 5951 13175
rect 8033 13141 8067 13175
rect 8953 13141 8987 13175
rect 9689 13141 9723 13175
rect 10517 13141 10551 13175
rect 10609 13141 10643 13175
rect 11345 13141 11379 13175
rect 13461 13141 13495 13175
rect 1409 12937 1443 12971
rect 1777 12937 1811 12971
rect 7849 12937 7883 12971
rect 6193 12869 6227 12903
rect 7941 12869 7975 12903
rect 13093 12869 13127 12903
rect 13369 12869 13403 12903
rect 1593 12801 1627 12835
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 2145 12801 2179 12835
rect 2329 12801 2363 12835
rect 3249 12801 3283 12835
rect 4077 12801 4111 12835
rect 4629 12801 4663 12835
rect 6101 12801 6135 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 6837 12801 6871 12835
rect 6981 12801 7015 12835
rect 7481 12801 7515 12835
rect 7737 12801 7771 12835
rect 8125 12801 8159 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 9137 12801 9171 12835
rect 9321 12801 9355 12835
rect 10241 12801 10275 12835
rect 11069 12801 11103 12835
rect 11529 12801 11563 12835
rect 12449 12801 12483 12835
rect 4353 12733 4387 12767
rect 6377 12733 6411 12767
rect 7297 12733 7331 12767
rect 8033 12733 8067 12767
rect 11253 12733 11287 12767
rect 3801 12665 3835 12699
rect 10609 12665 10643 12699
rect 13185 12665 13219 12699
rect 4445 12597 4479 12631
rect 7113 12597 7147 12631
rect 4721 12393 4755 12427
rect 6285 12393 6319 12427
rect 7205 12393 7239 12427
rect 7757 12393 7791 12427
rect 8953 12393 8987 12427
rect 9321 12393 9355 12427
rect 10425 12393 10459 12427
rect 2881 12325 2915 12359
rect 3433 12325 3467 12359
rect 3985 12325 4019 12359
rect 8217 12325 8251 12359
rect 9505 12325 9539 12359
rect 10057 12325 10091 12359
rect 13277 12325 13311 12359
rect 3525 12257 3559 12291
rect 7389 12257 7423 12291
rect 9597 12257 9631 12291
rect 10149 12257 10183 12291
rect 1409 12189 1443 12223
rect 2145 12189 2179 12223
rect 2973 12189 3007 12223
rect 4123 12189 4157 12223
rect 4353 12189 4387 12223
rect 4537 12189 4571 12223
rect 5089 12189 5123 12223
rect 5733 12189 5767 12223
rect 6653 12189 6687 12223
rect 6929 12189 6963 12223
rect 7073 12189 7107 12223
rect 8396 12189 8430 12223
rect 8493 12189 8527 12223
rect 8748 12189 8782 12223
rect 9137 12189 9171 12223
rect 10977 12189 11011 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 12909 12189 12943 12223
rect 2329 12121 2363 12155
rect 2697 12121 2731 12155
rect 4261 12121 4295 12155
rect 4905 12121 4939 12155
rect 6009 12121 6043 12155
rect 6377 12121 6411 12155
rect 6561 12121 6595 12155
rect 6837 12121 6871 12155
rect 7573 12121 7607 12155
rect 8585 12121 8619 12155
rect 10241 12121 10275 12155
rect 10793 12121 10827 12155
rect 2513 12053 2547 12087
rect 4629 12053 4663 12087
rect 7757 12053 7791 12087
rect 7941 12053 7975 12087
rect 10425 12053 10459 12087
rect 10609 12053 10643 12087
rect 6929 11849 6963 11883
rect 9229 11849 9263 11883
rect 11621 11849 11655 11883
rect 2237 11781 2271 11815
rect 2329 11781 2363 11815
rect 3525 11781 3559 11815
rect 4537 11781 4571 11815
rect 5457 11781 5491 11815
rect 6561 11781 6595 11815
rect 7757 11781 7791 11815
rect 10149 11781 10183 11815
rect 10333 11781 10367 11815
rect 10977 11781 11011 11815
rect 13001 11781 13035 11815
rect 13277 11781 13311 11815
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 3709 11713 3743 11747
rect 3801 11713 3835 11747
rect 4905 11713 4939 11747
rect 5273 11713 5307 11747
rect 5549 11713 5583 11747
rect 5824 11713 5858 11747
rect 5916 11735 5950 11769
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 6377 11713 6411 11747
rect 7113 11713 7147 11747
rect 7205 11713 7239 11747
rect 7941 11713 7975 11747
rect 8125 11713 8159 11747
rect 8217 11713 8251 11747
rect 8585 11713 8619 11747
rect 8677 11713 8711 11747
rect 9321 11713 9355 11747
rect 9689 11713 9723 11747
rect 9781 11713 9815 11747
rect 10701 11713 10735 11747
rect 10839 11713 10873 11747
rect 11074 11713 11108 11747
rect 11529 11713 11563 11747
rect 11737 11713 11771 11747
rect 12081 11713 12115 11747
rect 12909 11713 12943 11747
rect 1685 11645 1719 11679
rect 4353 11645 4387 11679
rect 7481 11645 7515 11679
rect 8309 11645 8343 11679
rect 9413 11645 9447 11679
rect 11821 11645 11855 11679
rect 12449 11645 12483 11679
rect 2145 11577 2179 11611
rect 4261 11577 4295 11611
rect 4721 11577 4755 11611
rect 8401 11577 8435 11611
rect 1593 11509 1627 11543
rect 5089 11509 5123 11543
rect 6653 11509 6687 11543
rect 7389 11509 7423 11543
rect 8861 11509 8895 11543
rect 9505 11509 9539 11543
rect 9965 11509 9999 11543
rect 10333 11509 10367 11543
rect 10517 11509 10551 11543
rect 11253 11509 11287 11543
rect 12081 11509 12115 11543
rect 13369 11509 13403 11543
rect 5733 11305 5767 11339
rect 8125 11305 8159 11339
rect 9137 11305 9171 11339
rect 10425 11305 10459 11339
rect 10793 11305 10827 11339
rect 12173 11305 12207 11339
rect 2697 11237 2731 11271
rect 5089 11237 5123 11271
rect 8309 11237 8343 11271
rect 3525 11169 3559 11203
rect 6193 11169 6227 11203
rect 6285 11169 6319 11203
rect 8033 11169 8067 11203
rect 9965 11169 9999 11203
rect 10333 11169 10367 11203
rect 11529 11169 11563 11203
rect 1409 11101 1443 11135
rect 2329 11101 2363 11135
rect 3065 11101 3099 11135
rect 3341 11101 3375 11135
rect 3801 11101 3835 11135
rect 4721 11101 4755 11135
rect 5963 11101 5997 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 6871 11101 6905 11135
rect 7205 11101 7239 11135
rect 7390 11101 7424 11135
rect 7481 11101 7515 11135
rect 7607 11101 7641 11135
rect 7941 11101 7975 11135
rect 9413 11101 9447 11135
rect 9597 11101 9631 11135
rect 9780 11101 9814 11135
rect 9873 11101 9907 11135
rect 10149 11101 10183 11135
rect 10425 11101 10459 11135
rect 10609 11101 10643 11135
rect 10977 11101 11011 11135
rect 11161 11101 11195 11135
rect 11437 11101 11471 11135
rect 11645 11101 11679 11135
rect 11759 11101 11793 11135
rect 11989 11101 12023 11135
rect 12357 11101 12391 11135
rect 13001 11101 13035 11135
rect 5733 11033 5767 11067
rect 7113 11033 7147 11067
rect 7849 11033 7883 11067
rect 8953 11033 8987 11067
rect 9137 11033 9171 11067
rect 13277 11033 13311 11067
rect 3157 10965 3191 10999
rect 6101 10965 6135 10999
rect 8585 10965 8619 10999
rect 8677 10965 8711 10999
rect 11253 10965 11287 10999
rect 13369 10965 13403 10999
rect 13461 10965 13495 10999
rect 3065 10761 3099 10795
rect 3617 10761 3651 10795
rect 4077 10761 4111 10795
rect 6193 10761 6227 10795
rect 10885 10761 10919 10795
rect 2605 10693 2639 10727
rect 3341 10693 3375 10727
rect 4261 10693 4295 10727
rect 5273 10693 5307 10727
rect 7021 10693 7055 10727
rect 7205 10693 7239 10727
rect 8217 10693 8251 10727
rect 8401 10693 8435 10727
rect 8585 10693 8619 10727
rect 8769 10693 8803 10727
rect 9137 10693 9171 10727
rect 9781 10693 9815 10727
rect 10241 10693 10275 10727
rect 11805 10693 11839 10727
rect 12725 10693 12759 10727
rect 13461 10693 13495 10727
rect 1633 10625 1667 10659
rect 1777 10625 1811 10659
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 3433 10625 3467 10659
rect 4169 10625 4203 10659
rect 4537 10625 4571 10659
rect 5181 10625 5215 10659
rect 7389 10625 7423 10659
rect 7665 10625 7699 10659
rect 7849 10625 7883 10659
rect 8033 10625 8067 10659
rect 8953 10625 8987 10659
rect 9689 10625 9723 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 10701 10625 10735 10659
rect 11161 10625 11195 10659
rect 11345 10625 11379 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11949 10625 11983 10659
rect 2145 10557 2179 10591
rect 2697 10557 2731 10591
rect 5365 10557 5399 10591
rect 5825 10557 5859 10591
rect 6929 10557 6963 10591
rect 9597 10557 9631 10591
rect 12265 10557 12299 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 1501 10489 1535 10523
rect 6469 10489 6503 10523
rect 6653 10489 6687 10523
rect 7665 10489 7699 10523
rect 10609 10489 10643 10523
rect 13369 10489 13403 10523
rect 2973 10421 3007 10455
rect 3801 10421 3835 10455
rect 6009 10421 6043 10455
rect 9321 10421 9355 10455
rect 9505 10421 9539 10455
rect 11069 10421 11103 10455
rect 12081 10421 12115 10455
rect 1501 10217 1535 10251
rect 3341 10217 3375 10251
rect 3617 10217 3651 10251
rect 3985 10217 4019 10251
rect 5641 10217 5675 10251
rect 6469 10217 6503 10251
rect 7389 10217 7423 10251
rect 8401 10217 8435 10251
rect 8585 10217 8619 10251
rect 11161 10217 11195 10251
rect 11805 10217 11839 10251
rect 2881 10149 2915 10183
rect 6837 10149 6871 10183
rect 7205 10149 7239 10183
rect 13277 10149 13311 10183
rect 4629 10081 4663 10115
rect 9045 10081 9079 10115
rect 10224 10081 10258 10115
rect 10517 10081 10551 10115
rect 1593 10013 1627 10047
rect 3065 10013 3099 10047
rect 4077 10013 4111 10047
rect 4905 10013 4939 10047
rect 5273 10013 5307 10047
rect 5917 10013 5951 10047
rect 6290 10013 6324 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 7021 10013 7055 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 7942 10013 7976 10047
rect 8677 10013 8711 10047
rect 8769 10013 8803 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9505 10013 9539 10047
rect 9597 10013 9631 10047
rect 10609 10013 10643 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11253 10013 11287 10047
rect 11529 10013 11563 10047
rect 11989 10013 12023 10047
rect 13369 10013 13403 10047
rect 4537 9945 4571 9979
rect 5089 9945 5123 9979
rect 5825 9945 5859 9979
rect 6101 9945 6135 9979
rect 6193 9945 6227 9979
rect 8217 9945 8251 9979
rect 9781 9945 9815 9979
rect 9965 9945 9999 9979
rect 11713 9945 11747 9979
rect 3249 9877 3283 9911
rect 4721 9877 4755 9911
rect 5457 9877 5491 9911
rect 5641 9877 5675 9911
rect 10333 9877 10367 9911
rect 10425 9877 10459 9911
rect 10885 9877 10919 9911
rect 1501 9673 1535 9707
rect 10885 9673 10919 9707
rect 13185 9673 13219 9707
rect 2973 9605 3007 9639
rect 6837 9605 6871 9639
rect 8125 9605 8159 9639
rect 9781 9605 9815 9639
rect 10517 9605 10551 9639
rect 10701 9605 10735 9639
rect 2145 9537 2179 9571
rect 2237 9537 2271 9571
rect 3157 9537 3191 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 5549 9537 5583 9571
rect 6193 9537 6227 9571
rect 6601 9537 6635 9571
rect 6745 9537 6779 9571
rect 7021 9537 7055 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 7936 9537 7970 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 8769 9537 8803 9571
rect 8953 9537 8987 9571
rect 9137 9537 9171 9571
rect 9413 9537 9447 9571
rect 9873 9537 9907 9571
rect 10057 9537 10091 9571
rect 10333 9537 10367 9571
rect 11161 9537 11195 9571
rect 11253 9537 11287 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 12081 9537 12115 9571
rect 12173 9537 12207 9571
rect 12817 9537 12851 9571
rect 13093 9537 13127 9571
rect 13369 9537 13403 9571
rect 3249 9469 3283 9503
rect 9229 9469 9263 9503
rect 1685 9401 1719 9435
rect 4905 9401 4939 9435
rect 7757 9401 7791 9435
rect 8493 9401 8527 9435
rect 11253 9401 11287 9435
rect 11713 9401 11747 9435
rect 2145 9333 2179 9367
rect 6469 9333 6503 9367
rect 8769 9333 8803 9367
rect 9413 9333 9447 9367
rect 9597 9333 9631 9367
rect 13553 9333 13587 9367
rect 1409 9129 1443 9163
rect 3341 9129 3375 9163
rect 4905 9129 4939 9163
rect 6101 9129 6135 9163
rect 9321 9129 9355 9163
rect 9873 9129 9907 9163
rect 11897 9129 11931 9163
rect 2881 9061 2915 9095
rect 4261 9061 4295 9095
rect 5549 9061 5583 9095
rect 5733 9061 5767 9095
rect 7481 9061 7515 9095
rect 8217 9061 8251 9095
rect 9597 9061 9631 9095
rect 10517 9061 10551 9095
rect 11621 9061 11655 9095
rect 2421 8993 2455 9027
rect 5089 8993 5123 9027
rect 5641 8993 5675 9027
rect 8493 8993 8527 9027
rect 12449 8993 12483 9027
rect 3249 8925 3283 8959
rect 4077 8925 4111 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 7665 8925 7699 8959
rect 8033 8925 8067 8959
rect 8309 8925 8343 8959
rect 8401 8925 8435 8959
rect 8953 8925 8987 8959
rect 9413 8925 9447 8959
rect 9689 8925 9723 8959
rect 9965 8925 9999 8959
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 11069 8925 11103 8959
rect 11345 8925 11379 8959
rect 11489 8925 11523 8959
rect 12081 8925 12115 8959
rect 13277 8925 13311 8959
rect 2973 8857 3007 8891
rect 3617 8857 3651 8891
rect 3801 8857 3835 8891
rect 6837 8857 6871 8891
rect 7849 8857 7883 8891
rect 10057 8857 10091 8891
rect 10701 8857 10735 8891
rect 10885 8857 10919 8891
rect 11253 8857 11287 8891
rect 12265 8857 12299 8891
rect 12357 8857 12391 8891
rect 12909 8857 12943 8891
rect 13001 8857 13035 8891
rect 13461 8857 13495 8891
rect 3065 8789 3099 8823
rect 3893 8789 3927 8823
rect 4537 8789 4571 8823
rect 7297 8789 7331 8823
rect 9045 8789 9079 8823
rect 5365 8585 5399 8619
rect 7389 8585 7423 8619
rect 10057 8585 10091 8619
rect 11529 8585 11563 8619
rect 11713 8585 11747 8619
rect 12265 8585 12299 8619
rect 6009 8517 6043 8551
rect 10977 8517 11011 8551
rect 13001 8517 13035 8551
rect 13369 8517 13403 8551
rect 1501 8449 1535 8483
rect 3525 8449 3559 8483
rect 4721 8449 4755 8483
rect 5273 8449 5307 8483
rect 5825 8449 5859 8483
rect 6837 8449 6871 8483
rect 7205 8449 7239 8483
rect 7573 8449 7607 8483
rect 7941 8449 7975 8483
rect 8585 8449 8619 8483
rect 9137 8449 9171 8483
rect 9413 8449 9447 8483
rect 9873 8449 9907 8483
rect 10057 8449 10091 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 11161 8449 11195 8483
rect 12081 8449 12115 8483
rect 12357 8449 12391 8483
rect 13277 8449 13311 8483
rect 7021 8381 7055 8415
rect 9781 8381 9815 8415
rect 10425 8381 10459 8415
rect 10517 8381 10551 8415
rect 3341 8313 3375 8347
rect 4813 8313 4847 8347
rect 5733 8313 5767 8347
rect 6377 8313 6411 8347
rect 6929 8313 6963 8347
rect 11345 8313 11379 8347
rect 11989 8313 12023 8347
rect 13461 8313 13495 8347
rect 6101 8245 6135 8279
rect 1501 8041 1535 8075
rect 3617 8041 3651 8075
rect 11345 8041 11379 8075
rect 4537 7973 4571 8007
rect 13185 7973 13219 8007
rect 4077 7905 4111 7939
rect 4629 7905 4663 7939
rect 6837 7905 6871 7939
rect 9597 7905 9631 7939
rect 2145 7837 2179 7871
rect 2789 7837 2823 7871
rect 3157 7837 3191 7871
rect 3341 7837 3375 7871
rect 4721 7837 4755 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 6193 7837 6227 7871
rect 6377 7837 6411 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 8309 7837 8343 7871
rect 8493 7837 8527 7871
rect 9393 7837 9427 7871
rect 9689 7837 9723 7871
rect 10149 7837 10183 7871
rect 10425 7837 10459 7871
rect 11437 7837 11471 7871
rect 11805 7837 11839 7871
rect 11897 7837 11931 7871
rect 12909 7837 12943 7871
rect 2605 7769 2639 7803
rect 2973 7769 3007 7803
rect 3065 7769 3099 7803
rect 8953 7769 8987 7803
rect 9137 7769 9171 7803
rect 11621 7769 11655 7803
rect 3893 7701 3927 7735
rect 8217 7701 8251 7735
rect 8677 7701 8711 7735
rect 9505 7701 9539 7735
rect 10977 7701 11011 7735
rect 2237 7497 2271 7531
rect 2421 7497 2455 7531
rect 2973 7497 3007 7531
rect 7941 7497 7975 7531
rect 9045 7497 9079 7531
rect 5365 7429 5399 7463
rect 5641 7429 5675 7463
rect 10333 7429 10367 7463
rect 12357 7429 12391 7463
rect 1961 7361 1995 7395
rect 2145 7361 2179 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4169 7361 4203 7395
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5825 7361 5859 7395
rect 6193 7361 6227 7395
rect 6837 7361 6871 7395
rect 6929 7361 6963 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 7829 7361 7863 7395
rect 8033 7361 8067 7395
rect 8493 7361 8527 7395
rect 9195 7361 9229 7395
rect 9602 7361 9636 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10058 7361 10092 7395
rect 3065 7293 3099 7327
rect 3249 7293 3283 7327
rect 3433 7293 3467 7327
rect 4353 7293 4387 7327
rect 5457 7293 5491 7327
rect 7113 7293 7147 7327
rect 7205 7293 7239 7327
rect 8125 7293 8159 7327
rect 8677 7293 8711 7327
rect 9485 7293 9519 7327
rect 11805 7293 11839 7327
rect 12449 7293 12483 7327
rect 12817 7293 12851 7327
rect 12909 7293 12943 7327
rect 6009 7225 6043 7259
rect 12265 7225 12299 7259
rect 1777 7157 1811 7191
rect 2605 7157 2639 7191
rect 4721 7157 4755 7191
rect 6653 7157 6687 7191
rect 8309 7157 8343 7191
rect 12817 7157 12851 7191
rect 2040 6953 2074 6987
rect 3525 6953 3559 6987
rect 6088 6953 6122 6987
rect 13277 6885 13311 6919
rect 1777 6817 1811 6851
rect 3801 6817 3835 6851
rect 5825 6817 5859 6851
rect 7573 6817 7607 6851
rect 8033 6817 8067 6851
rect 9229 6817 9263 6851
rect 11621 6817 11655 6851
rect 8217 6749 8251 6783
rect 8585 6749 8619 6783
rect 9413 6749 9447 6783
rect 9873 6749 9907 6783
rect 11989 6749 12023 6783
rect 13461 6749 13495 6783
rect 4077 6681 4111 6715
rect 10149 6681 10183 6715
rect 1409 6613 1443 6647
rect 1685 6613 1719 6647
rect 5549 6613 5583 6647
rect 8493 6613 8527 6647
rect 9321 6613 9355 6647
rect 9781 6613 9815 6647
rect 4077 6409 4111 6443
rect 4537 6409 4571 6443
rect 6653 6409 6687 6443
rect 7297 6409 7331 6443
rect 11345 6409 11379 6443
rect 3985 6341 4019 6375
rect 5181 6341 5215 6375
rect 9045 6341 9079 6375
rect 11989 6341 12023 6375
rect 12449 6341 12483 6375
rect 13093 6341 13127 6375
rect 1835 6273 1869 6307
rect 1961 6273 1995 6307
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 3249 6273 3283 6307
rect 3801 6273 3835 6307
rect 4445 6273 4479 6307
rect 5733 6273 5767 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 7113 6273 7147 6307
rect 7389 6273 7423 6307
rect 7481 6273 7515 6307
rect 7757 6273 7791 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 9505 6273 9539 6307
rect 9781 6273 9815 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 10701 6273 10735 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12173 6273 12207 6307
rect 12265 6273 12299 6307
rect 12633 6273 12667 6307
rect 2605 6205 2639 6239
rect 4721 6205 4755 6239
rect 9137 6205 9171 6239
rect 13185 6205 13219 6239
rect 1593 6137 1627 6171
rect 2421 6137 2455 6171
rect 3617 6137 3651 6171
rect 10517 6137 10551 6171
rect 11621 6137 11655 6171
rect 1409 6069 1443 6103
rect 2789 6069 2823 6103
rect 4905 6069 4939 6103
rect 6377 6069 6411 6103
rect 10885 6069 10919 6103
rect 1685 5865 1719 5899
rect 6561 5865 6595 5899
rect 9229 5865 9263 5899
rect 9505 5865 9539 5899
rect 12081 5865 12115 5899
rect 13277 5865 13311 5899
rect 2237 5797 2271 5831
rect 3341 5797 3375 5831
rect 10057 5797 10091 5831
rect 4813 5729 4847 5763
rect 8217 5729 8251 5763
rect 8309 5729 8343 5763
rect 10333 5729 10367 5763
rect 10609 5729 10643 5763
rect 1869 5661 1903 5695
rect 1961 5661 1995 5695
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 4445 5661 4479 5695
rect 7021 5661 7055 5695
rect 7481 5661 7515 5695
rect 9045 5661 9079 5695
rect 9321 5661 9355 5695
rect 9687 5661 9721 5695
rect 10149 5661 10183 5695
rect 3801 5593 3835 5627
rect 3985 5593 4019 5627
rect 4353 5593 4387 5627
rect 5089 5593 5123 5627
rect 8401 5593 8435 5627
rect 1501 5525 1535 5559
rect 2697 5525 2731 5559
rect 4077 5525 4111 5559
rect 4169 5525 4203 5559
rect 4537 5525 4571 5559
rect 7849 5525 7883 5559
rect 8769 5525 8803 5559
rect 9689 5525 9723 5559
rect 13185 5525 13219 5559
rect 2697 5321 2731 5355
rect 4905 5321 4939 5355
rect 5457 5321 5491 5355
rect 12274 5321 12308 5355
rect 1961 5253 1995 5287
rect 2789 5253 2823 5287
rect 3985 5253 4019 5287
rect 4261 5253 4295 5287
rect 8861 5253 8895 5287
rect 9781 5253 9815 5287
rect 11529 5253 11563 5287
rect 11713 5253 11747 5287
rect 11897 5253 11931 5287
rect 13277 5253 13311 5287
rect 1777 5185 1811 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 3617 5185 3651 5219
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 4169 5185 4203 5219
rect 4445 5185 4479 5219
rect 5089 5185 5123 5219
rect 5181 5185 5215 5219
rect 5917 5185 5951 5219
rect 6561 5185 6595 5219
rect 6929 5185 6963 5219
rect 9045 5185 9079 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 12633 5185 12667 5219
rect 13553 5185 13587 5219
rect 2588 5117 2622 5151
rect 2881 5117 2915 5151
rect 5641 5117 5675 5151
rect 6377 5117 6411 5151
rect 7205 5117 7239 5151
rect 1593 5049 1627 5083
rect 3249 5049 3283 5083
rect 5825 5049 5859 5083
rect 6745 5049 6779 5083
rect 11253 5049 11287 5083
rect 2145 4981 2179 5015
rect 4629 4981 4663 5015
rect 8677 4981 8711 5015
rect 12265 4981 12299 5015
rect 12449 4981 12483 5015
rect 7297 4777 7331 4811
rect 8493 4777 8527 4811
rect 9229 4777 9263 4811
rect 12081 4777 12115 4811
rect 2881 4709 2915 4743
rect 2969 4709 3003 4743
rect 3249 4709 3283 4743
rect 6745 4709 6779 4743
rect 13185 4709 13219 4743
rect 1869 4641 1903 4675
rect 3801 4641 3835 4675
rect 6837 4641 6871 4675
rect 7757 4641 7791 4675
rect 7941 4641 7975 4675
rect 10333 4641 10367 4675
rect 10609 4641 10643 4675
rect 1777 4573 1811 4607
rect 2053 4573 2087 4607
rect 2421 4573 2455 4607
rect 2605 4573 2639 4607
rect 2789 4573 2823 4607
rect 3065 4573 3099 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6010 4551 6044 4585
rect 6135 4573 6169 4607
rect 6561 4573 6595 4607
rect 7665 4573 7699 4607
rect 8585 4573 8619 4607
rect 9229 4573 9263 4607
rect 9597 4573 9631 4607
rect 9689 4573 9723 4607
rect 10057 4573 10091 4607
rect 10241 4573 10275 4607
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 13553 4573 13587 4607
rect 4077 4505 4111 4539
rect 6377 4505 6411 4539
rect 8769 4505 8803 4539
rect 9873 4505 9907 4539
rect 12265 4505 12299 4539
rect 13277 4505 13311 4539
rect 1409 4437 1443 4471
rect 2605 4437 2639 4471
rect 3525 4437 3559 4471
rect 5549 4437 5583 4471
rect 8125 4437 8159 4471
rect 9045 4437 9079 4471
rect 13369 4437 13403 4471
rect 1501 4233 1535 4267
rect 4537 4233 4571 4267
rect 4997 4233 5031 4267
rect 5733 4233 5767 4267
rect 6469 4233 6503 4267
rect 8585 4233 8619 4267
rect 9229 4233 9263 4267
rect 11621 4233 11655 4267
rect 12909 4233 12943 4267
rect 13093 4233 13127 4267
rect 13277 4233 13311 4267
rect 4077 4165 4111 4199
rect 4445 4165 4479 4199
rect 11989 4165 12023 4199
rect 12541 4165 12575 4199
rect 1593 4097 1627 4131
rect 1777 4097 1811 4131
rect 2145 4097 2179 4131
rect 2329 4097 2363 4131
rect 2513 4097 2547 4131
rect 3433 4097 3467 4131
rect 4261 4097 4295 4131
rect 4905 4097 4939 4131
rect 5549 4097 5583 4131
rect 5641 4097 5675 4131
rect 5917 4097 5951 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 8585 4097 8619 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 11621 4097 11655 4131
rect 11897 4097 11931 4131
rect 12081 4097 12115 4131
rect 12265 4097 12299 4131
rect 12725 4097 12759 4131
rect 13001 4097 13035 4131
rect 2789 4029 2823 4063
rect 3341 4029 3375 4063
rect 5181 4029 5215 4063
rect 6101 4029 6135 4063
rect 7941 4029 7975 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 9413 3961 9447 3995
rect 1777 3893 1811 3927
rect 1961 3893 1995 3927
rect 8861 3893 8895 3927
rect 11253 3893 11287 3927
rect 13553 3893 13587 3927
rect 2237 3689 2271 3723
rect 2697 3689 2731 3723
rect 4077 3689 4111 3723
rect 9137 3689 9171 3723
rect 9321 3689 9355 3723
rect 9689 3689 9723 3723
rect 10333 3689 10367 3723
rect 12817 3689 12851 3723
rect 13001 3689 13035 3723
rect 1685 3621 1719 3655
rect 2881 3621 2915 3655
rect 3341 3621 3375 3655
rect 6285 3621 6319 3655
rect 10057 3621 10091 3655
rect 2027 3553 2061 3587
rect 2605 3553 2639 3587
rect 5457 3553 5491 3587
rect 6837 3553 6871 3587
rect 8769 3553 8803 3587
rect 10425 3553 10459 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1869 3485 1903 3519
rect 2237 3485 2271 3519
rect 2513 3485 2547 3519
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 4261 3485 4295 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6193 3485 6227 3519
rect 6377 3485 6411 3519
rect 6469 3485 6503 3519
rect 6653 3485 6687 3519
rect 9873 3485 9907 3519
rect 10149 3485 10183 3519
rect 12449 3485 12483 3519
rect 12725 3485 12759 3519
rect 3065 3417 3099 3451
rect 4997 3417 5031 3451
rect 8493 3417 8527 3451
rect 9505 3417 9539 3451
rect 10701 3417 10735 3451
rect 12357 3417 12391 3451
rect 7021 3349 7055 3383
rect 9321 3349 9355 3383
rect 12173 3349 12207 3383
rect 2329 3145 2363 3179
rect 5181 3145 5215 3179
rect 6101 3145 6135 3179
rect 7481 3145 7515 3179
rect 7941 3145 7975 3179
rect 10057 3145 10091 3179
rect 10609 3145 10643 3179
rect 11069 3145 11103 3179
rect 11345 3145 11379 3179
rect 2881 3077 2915 3111
rect 2973 3077 3007 3111
rect 3249 3077 3283 3111
rect 3709 3077 3743 3111
rect 4905 3077 4939 3111
rect 5733 3077 5767 3111
rect 5917 3077 5951 3111
rect 1501 3009 1535 3043
rect 1777 3009 1811 3043
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 3433 3009 3467 3043
rect 3617 3009 3651 3043
rect 4169 3009 4203 3043
rect 4537 3009 4571 3043
rect 5365 3009 5399 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 10701 3009 10735 3043
rect 11621 3009 11655 3043
rect 11897 3009 11931 3043
rect 12633 3009 12667 3043
rect 1593 2941 1627 2975
rect 2697 2941 2731 2975
rect 5549 2941 5583 2975
rect 7021 2941 7055 2975
rect 7573 2941 7607 2975
rect 8585 2941 8619 2975
rect 10517 2941 10551 2975
rect 11989 2941 12023 2975
rect 12725 2941 12759 2975
rect 6837 2873 6871 2907
rect 11621 2873 11655 2907
rect 2053 2805 2087 2839
rect 5917 2805 5951 2839
rect 1501 2601 1535 2635
rect 2421 2601 2455 2635
rect 4169 2601 4203 2635
rect 8401 2601 8435 2635
rect 8953 2601 8987 2635
rect 10333 2601 10367 2635
rect 2237 2465 2271 2499
rect 3249 2465 3283 2499
rect 3433 2465 3467 2499
rect 5549 2465 5583 2499
rect 8677 2465 8711 2499
rect 9597 2465 9631 2499
rect 9781 2465 9815 2499
rect 10701 2465 10735 2499
rect 12173 2465 12207 2499
rect 13185 2465 13219 2499
rect 1777 2397 1811 2431
rect 1961 2397 1995 2431
rect 2053 2397 2087 2431
rect 2329 2397 2363 2431
rect 2513 2397 2547 2431
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 5365 2397 5399 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 8033 2397 8067 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 10425 2397 10459 2431
rect 1593 2329 1627 2363
rect 4629 2329 4663 2363
rect 5825 2329 5859 2363
rect 8125 2329 8159 2363
rect 8309 2329 8343 2363
rect 12357 2329 12391 2363
rect 2789 2261 2823 2295
rect 3157 2261 3191 2295
rect 7297 2261 7331 2295
rect 7941 2261 7975 2295
rect 9413 2261 9447 2295
rect 3525 2057 3559 2091
rect 3617 2057 3651 2091
rect 5549 2057 5583 2091
rect 6101 2057 6135 2091
rect 6469 2057 6503 2091
rect 10241 2057 10275 2091
rect 10977 2057 11011 2091
rect 13277 2057 13311 2091
rect 8125 1989 8159 2023
rect 3341 1921 3375 1955
rect 3801 1921 3835 1955
rect 5917 1921 5951 1955
rect 6009 1921 6043 1955
rect 10517 1921 10551 1955
rect 10701 1921 10735 1955
rect 10977 1921 11011 1955
rect 11161 1921 11195 1955
rect 11529 1921 11563 1955
rect 2697 1853 2731 1887
rect 4077 1853 4111 1887
rect 8401 1853 8435 1887
rect 8493 1853 8527 1887
rect 8769 1853 8803 1887
rect 10425 1853 10459 1887
rect 11805 1853 11839 1887
rect 6653 1717 6687 1751
rect 3893 1513 3927 1547
rect 4721 1513 4755 1547
rect 5641 1513 5675 1547
rect 8493 1513 8527 1547
rect 9768 1513 9802 1547
rect 11253 1513 11287 1547
rect 12541 1513 12575 1547
rect 12725 1513 12759 1547
rect 13093 1513 13127 1547
rect 3525 1445 3559 1479
rect 8953 1445 8987 1479
rect 2053 1377 2087 1411
rect 5365 1377 5399 1411
rect 7205 1377 7239 1411
rect 7665 1377 7699 1411
rect 7941 1377 7975 1411
rect 9505 1377 9539 1411
rect 1501 1309 1535 1343
rect 1777 1309 1811 1343
rect 3801 1309 3835 1343
rect 3985 1309 4019 1343
rect 4261 1309 4295 1343
rect 4445 1309 4479 1343
rect 4629 1309 4663 1343
rect 5089 1309 5123 1343
rect 5549 1309 5583 1343
rect 5917 1309 5951 1343
rect 6193 1309 6227 1343
rect 7113 1309 7147 1343
rect 8125 1309 8159 1343
rect 8309 1309 8343 1343
rect 8401 1309 8435 1343
rect 8677 1309 8711 1343
rect 9137 1309 9171 1343
rect 11621 1309 11655 1343
rect 11805 1309 11839 1343
rect 11989 1309 12023 1343
rect 12173 1309 12207 1343
rect 12357 1309 12391 1343
rect 5181 1241 5215 1275
rect 9321 1241 9355 1275
rect 6469 1173 6503 1207
rect 12173 1173 12207 1207
rect 12909 1173 12943 1207
<< metal1 >>
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 12066 13852 12072 13864
rect 9456 13824 12072 13852
rect 9456 13812 9462 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 9950 13784 9956 13796
rect 2096 13756 9956 13784
rect 2096 13744 2102 13756
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 7098 13716 7104 13728
rect 1728 13688 7104 13716
rect 1728 13676 1734 13688
rect 7098 13676 7104 13688
rect 7156 13716 7162 13728
rect 7374 13716 7380 13728
rect 7156 13688 7380 13716
rect 7156 13676 7162 13688
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 11790 13716 11796 13728
rect 7524 13688 11796 13716
rect 7524 13676 7530 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 566 13472 572 13524
rect 624 13512 630 13524
rect 3513 13515 3571 13521
rect 3513 13512 3525 13515
rect 624 13484 3525 13512
rect 624 13472 630 13484
rect 3513 13481 3525 13484
rect 3559 13512 3571 13515
rect 3559 13484 6868 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13444 2743 13447
rect 4062 13444 4068 13456
rect 2731 13416 4068 13444
rect 2731 13413 2743 13416
rect 2685 13407 2743 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 6638 13444 6644 13456
rect 4908 13416 6644 13444
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 4706 13376 4712 13388
rect 3375 13348 4712 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2372 13280 2789 13308
rect 2372 13268 2378 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 3786 13308 3792 13320
rect 3747 13280 3792 13308
rect 2777 13271 2835 13277
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 3970 13308 3976 13320
rect 3927 13280 3976 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4614 13308 4620 13320
rect 4111 13280 4522 13308
rect 4575 13280 4620 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 1452 13212 1501 13240
rect 1452 13200 1458 13212
rect 1489 13209 1501 13212
rect 1535 13209 1547 13243
rect 1489 13203 1547 13209
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13240 1639 13243
rect 2130 13240 2136 13252
rect 1627 13212 2136 13240
rect 1627 13209 1639 13212
rect 1581 13203 1639 13209
rect 2130 13200 2136 13212
rect 2188 13200 2194 13252
rect 3234 13240 3240 13252
rect 3195 13212 3240 13240
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 4212 13212 4261 13240
rect 4212 13200 4218 13212
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 4494 13240 4522 13280
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 4908 13240 4936 13416
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13376 5227 13379
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 5215 13348 6469 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 5258 13308 5264 13320
rect 5219 13280 5264 13308
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 6086 13308 6092 13320
rect 5736 13280 5948 13308
rect 6047 13280 6092 13308
rect 5736 13252 5764 13280
rect 5074 13240 5080 13252
rect 4494 13212 4936 13240
rect 5035 13212 5080 13240
rect 4249 13203 4307 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5718 13240 5724 13252
rect 5679 13212 5724 13240
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 5813 13243 5871 13249
rect 5813 13209 5825 13243
rect 5859 13209 5871 13243
rect 5920 13240 5948 13280
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6730 13308 6736 13320
rect 6691 13280 6736 13308
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 6840 13308 6868 13484
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7432 13484 7849 13512
rect 7432 13472 7438 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 7837 13475 7895 13481
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 9398 13512 9404 13524
rect 9263 13484 9404 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9585 13515 9643 13521
rect 9585 13481 9597 13515
rect 9631 13512 9643 13515
rect 11330 13512 11336 13524
rect 9631 13484 11336 13512
rect 9631 13481 9643 13484
rect 9585 13475 9643 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 7285 13447 7343 13453
rect 7285 13413 7297 13447
rect 7331 13444 7343 13447
rect 9306 13444 9312 13456
rect 7331 13416 9312 13444
rect 7331 13413 7343 13416
rect 7285 13407 7343 13413
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 9548 13416 10364 13444
rect 9548 13404 9554 13416
rect 7745 13379 7803 13385
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 9030 13376 9036 13388
rect 7791 13348 9036 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 9030 13336 9036 13348
rect 9088 13336 9094 13388
rect 10137 13345 10195 13351
rect 7106 13311 7164 13317
rect 7106 13308 7118 13311
rect 6840 13280 7118 13308
rect 7106 13277 7118 13280
rect 7152 13277 7164 13311
rect 7106 13271 7164 13277
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 8168 13280 8217 13308
rect 8168 13268 8174 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8846 13308 8852 13320
rect 8711 13280 8852 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8846 13268 8852 13280
rect 8904 13308 8910 13320
rect 9401 13311 9459 13317
rect 8904 13280 9352 13308
rect 8904 13268 8910 13280
rect 6365 13243 6423 13249
rect 6365 13240 6377 13243
rect 5920 13212 6377 13240
rect 5813 13203 5871 13209
rect 6365 13209 6377 13212
rect 6411 13209 6423 13243
rect 6914 13240 6920 13252
rect 6875 13212 6920 13240
rect 6365 13203 6423 13209
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 2501 13175 2559 13181
rect 2280 13144 2325 13172
rect 2280 13132 2286 13144
rect 2501 13141 2513 13175
rect 2547 13172 2559 13175
rect 2774 13172 2780 13184
rect 2547 13144 2780 13172
rect 2547 13141 2559 13144
rect 2501 13135 2559 13141
rect 2774 13132 2780 13144
rect 2832 13132 2838 13184
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 4430 13172 4436 13184
rect 2924 13144 4436 13172
rect 2924 13132 2930 13144
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 5828 13172 5856 13203
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13209 7067 13243
rect 7558 13240 7564 13252
rect 7519 13212 7564 13240
rect 7009 13203 7067 13209
rect 5905 13175 5963 13181
rect 5905 13172 5917 13175
rect 5828 13144 5917 13172
rect 5905 13141 5917 13144
rect 5951 13141 5963 13175
rect 5905 13135 5963 13141
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7024 13172 7052 13203
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 9324 13240 9352 13280
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 10137 13311 10149 13345
rect 10183 13311 10195 13345
rect 10137 13308 10195 13311
rect 10226 13308 10232 13320
rect 9447 13280 10088 13308
rect 10137 13305 10232 13308
rect 10152 13280 10232 13305
rect 9447 13277 9459 13280
rect 9401 13271 9459 13277
rect 9950 13240 9956 13252
rect 8812 13212 8857 13240
rect 9324 13212 9812 13240
rect 9911 13212 9956 13240
rect 8812 13200 8818 13212
rect 7374 13172 7380 13184
rect 6880 13144 7380 13172
rect 6880 13132 6886 13144
rect 7374 13132 7380 13144
rect 7432 13172 7438 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 7432 13144 8033 13172
rect 7432 13132 7438 13144
rect 8021 13141 8033 13144
rect 8067 13172 8079 13175
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 8067 13144 8953 13172
rect 8067 13141 8079 13144
rect 8021 13135 8079 13141
rect 8941 13141 8953 13144
rect 8987 13172 8999 13175
rect 9490 13172 9496 13184
rect 8987 13144 9496 13172
rect 8987 13141 8999 13144
rect 8941 13135 8999 13141
rect 9490 13132 9496 13144
rect 9548 13172 9554 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 9548 13144 9689 13172
rect 9548 13132 9554 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9784 13172 9812 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10060 13240 10088 13280
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10336 13317 10364 13416
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 11011 13348 12725 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 11146 13308 11152 13320
rect 11107 13280 11152 13308
rect 10321 13271 10379 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 12066 13308 12072 13320
rect 11440 13280 11652 13308
rect 12027 13280 12072 13308
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 10060 13212 10425 13240
rect 10413 13209 10425 13212
rect 10459 13240 10471 13243
rect 10870 13240 10876 13252
rect 10459 13212 10876 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 11057 13243 11115 13249
rect 11057 13209 11069 13243
rect 11103 13240 11115 13243
rect 11440 13240 11468 13280
rect 11624 13252 11652 13280
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12216 13280 12261 13308
rect 12406 13280 12817 13308
rect 12216 13268 12222 13280
rect 11103 13212 11468 13240
rect 11517 13243 11575 13249
rect 11103 13209 11115 13212
rect 11057 13203 11115 13209
rect 11517 13209 11529 13243
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 10505 13175 10563 13181
rect 10505 13172 10517 13175
rect 9784 13144 10517 13172
rect 9677 13135 9735 13141
rect 10505 13141 10517 13144
rect 10551 13141 10563 13175
rect 10505 13135 10563 13141
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 11333 13175 11391 13181
rect 10652 13144 10697 13172
rect 10652 13132 10658 13144
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11532 13172 11560 13203
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 11664 13212 11709 13240
rect 11664 13200 11670 13212
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12406 13240 12434 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12618 13240 12624 13252
rect 11848 13212 12434 13240
rect 12579 13212 12624 13240
rect 11848 13200 11854 13212
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 13262 13240 13268 13252
rect 13223 13212 13268 13240
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13412 13212 13457 13240
rect 13412 13200 13418 13212
rect 11379 13144 11560 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 13449 13175 13507 13181
rect 13449 13172 13461 13175
rect 13228 13144 13461 13172
rect 13228 13132 13234 13144
rect 13449 13141 13461 13144
rect 13495 13141 13507 13175
rect 13449 13135 13507 13141
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 1394 12968 1400 12980
rect 1355 12940 1400 12968
rect 1394 12928 1400 12940
rect 1452 12928 1458 12980
rect 1765 12971 1823 12977
rect 1765 12937 1777 12971
rect 1811 12968 1823 12971
rect 2774 12968 2780 12980
rect 1811 12940 2780 12968
rect 1811 12937 1823 12940
rect 1765 12931 1823 12937
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 7006 12968 7012 12980
rect 4488 12940 7012 12968
rect 4488 12928 4494 12940
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7340 12940 7849 12968
rect 7340 12928 7346 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 7837 12931 7895 12937
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9088 12940 10272 12968
rect 9088 12928 9094 12940
rect 1964 12872 5028 12900
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 1964 12841 1992 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2314 12832 2320 12844
rect 2179 12804 2320 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 1394 12724 1400 12776
rect 1452 12764 1458 12776
rect 1688 12764 1716 12795
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 2924 12804 3249 12832
rect 2924 12792 2930 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 3237 12795 3295 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4614 12832 4620 12844
rect 4575 12804 4620 12832
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5000 12832 5028 12872
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 6181 12903 6239 12909
rect 6181 12900 6193 12903
rect 5132 12872 6193 12900
rect 5132 12860 5138 12872
rect 6181 12869 6193 12872
rect 6227 12900 6239 12903
rect 7558 12900 7564 12912
rect 6227 12872 7564 12900
rect 6227 12869 6239 12872
rect 6181 12863 6239 12869
rect 7558 12860 7564 12872
rect 7616 12860 7622 12912
rect 7929 12903 7987 12909
rect 7668 12872 7880 12900
rect 5534 12832 5540 12844
rect 5000 12804 5540 12832
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 6086 12832 6092 12844
rect 5684 12804 6092 12832
rect 5684 12792 5690 12804
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 1452 12736 1716 12764
rect 1452 12724 1458 12736
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4028 12736 4353 12764
rect 4028 12724 4034 12736
rect 4341 12733 4353 12736
rect 4387 12764 4399 12767
rect 6365 12767 6423 12773
rect 6365 12764 6377 12767
rect 4387 12736 6377 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 6365 12733 6377 12736
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 3789 12699 3847 12705
rect 3789 12696 3801 12699
rect 3292 12668 3801 12696
rect 3292 12656 3298 12668
rect 3789 12665 3801 12668
rect 3835 12696 3847 12699
rect 4798 12696 4804 12708
rect 3835 12668 4804 12696
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12628 4491 12631
rect 4982 12628 4988 12640
rect 4479 12600 4988 12628
rect 4479 12597 4491 12600
rect 4433 12591 4491 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6380 12628 6408 12727
rect 6564 12696 6592 12795
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6696 12804 6745 12832
rect 6696 12792 6702 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6748 12764 6776 12795
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7006 12841 7012 12844
rect 6969 12835 7012 12841
rect 6880 12804 6925 12832
rect 6880 12792 6886 12804
rect 6969 12801 6981 12835
rect 6969 12795 7012 12801
rect 7006 12792 7012 12795
rect 7064 12792 7070 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7432 12804 7481 12832
rect 7432 12792 7438 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7285 12767 7343 12773
rect 6748 12736 7253 12764
rect 6914 12696 6920 12708
rect 6564 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7225 12696 7253 12736
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7668 12764 7696 12872
rect 7725 12835 7783 12841
rect 7725 12801 7737 12835
rect 7771 12832 7783 12835
rect 7852 12832 7880 12872
rect 7929 12869 7941 12903
rect 7975 12900 7987 12903
rect 8938 12900 8944 12912
rect 7975 12872 8944 12900
rect 7975 12869 7987 12872
rect 7929 12863 7987 12869
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9674 12900 9680 12912
rect 9232 12872 9680 12900
rect 8110 12832 8116 12844
rect 7771 12801 7788 12832
rect 7852 12804 8116 12832
rect 7725 12795 7788 12801
rect 7331 12736 7696 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7374 12696 7380 12708
rect 7225 12668 7380 12696
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 6822 12628 6828 12640
rect 6380 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7466 12628 7472 12640
rect 7147 12600 7472 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7760 12628 7788 12795
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9030 12832 9036 12844
rect 8991 12804 9036 12832
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9232 12832 9260 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 9309 12835 9367 12841
rect 9180 12804 9273 12832
rect 9180 12792 9186 12804
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 9398 12832 9404 12844
rect 9355 12804 9404 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 10244 12841 10272 12940
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10962 12968 10968 12980
rect 10376 12940 10968 12968
rect 10376 12928 10382 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12676 12872 13093 12900
rect 12676 12860 12682 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 13127 12872 13369 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 13357 12863 13415 12869
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10520 12804 10824 12832
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 10520 12764 10548 12804
rect 8067 12736 10548 12764
rect 10796 12764 10824 12804
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10928 12804 11069 12832
rect 10928 12792 10934 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11514 12832 11520 12844
rect 11475 12804 11520 12832
rect 11057 12795 11115 12801
rect 11514 12792 11520 12804
rect 11572 12832 11578 12844
rect 12158 12832 12164 12844
rect 11572 12804 12164 12832
rect 11572 12792 11578 12804
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 10796 12736 11100 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 11072 12708 11100 12736
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11204 12736 11253 12764
rect 11204 12724 11210 12736
rect 11241 12733 11253 12736
rect 11287 12764 11299 12767
rect 11882 12764 11888 12776
rect 11287 12736 11888 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11882 12724 11888 12736
rect 11940 12764 11946 12776
rect 12452 12764 12480 12795
rect 11940 12736 12480 12764
rect 11940 12724 11946 12736
rect 8478 12656 8484 12708
rect 8536 12696 8542 12708
rect 8846 12696 8852 12708
rect 8536 12668 8852 12696
rect 8536 12656 8542 12668
rect 8846 12656 8852 12668
rect 8904 12696 8910 12708
rect 8904 12668 9674 12696
rect 8904 12656 8910 12668
rect 9646 12640 9674 12668
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10100 12668 10609 12696
rect 10100 12656 10106 12668
rect 10597 12665 10609 12668
rect 10643 12696 10655 12699
rect 10870 12696 10876 12708
rect 10643 12668 10876 12696
rect 10643 12665 10655 12668
rect 10597 12659 10655 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 11054 12656 11060 12708
rect 11112 12656 11118 12708
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 13173 12699 13231 12705
rect 13173 12696 13185 12699
rect 12952 12668 13185 12696
rect 12952 12656 12958 12668
rect 13173 12665 13185 12668
rect 13219 12665 13231 12699
rect 13173 12659 13231 12665
rect 9122 12628 9128 12640
rect 7760 12600 9128 12628
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9582 12588 9588 12640
rect 9640 12628 9674 12640
rect 10410 12628 10416 12640
rect 9640 12600 10416 12628
rect 9640 12588 9646 12600
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 4706 12424 4712 12436
rect 4667 12396 4712 12424
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 6273 12427 6331 12433
rect 6273 12393 6285 12427
rect 6319 12424 6331 12427
rect 6730 12424 6736 12436
rect 6319 12396 6736 12424
rect 6319 12393 6331 12396
rect 6273 12387 6331 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7745 12427 7803 12433
rect 7745 12393 7757 12427
rect 7791 12424 7803 12427
rect 8478 12424 8484 12436
rect 7791 12396 8484 12424
rect 7791 12393 7803 12396
rect 7745 12387 7803 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8812 12396 8953 12424
rect 8812 12384 8818 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 9180 12396 9321 12424
rect 9180 12384 9186 12396
rect 9309 12393 9321 12396
rect 9355 12424 9367 12427
rect 10410 12424 10416 12436
rect 9355 12396 10180 12424
rect 10371 12396 10416 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 2866 12356 2872 12368
rect 2827 12328 2872 12356
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 3421 12359 3479 12365
rect 3421 12325 3433 12359
rect 3467 12356 3479 12359
rect 3602 12356 3608 12368
rect 3467 12328 3608 12356
rect 3467 12325 3479 12328
rect 3421 12319 3479 12325
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 3973 12359 4031 12365
rect 3973 12325 3985 12359
rect 4019 12356 4031 12359
rect 4614 12356 4620 12368
rect 4019 12328 4620 12356
rect 4019 12325 4031 12328
rect 3973 12319 4031 12325
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 5258 12356 5264 12368
rect 5092 12328 5264 12356
rect 2038 12288 2044 12300
rect 1412 12260 2044 12288
rect 1412 12229 1440 12260
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 3510 12288 3516 12300
rect 3471 12260 3516 12288
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 4540 12260 5028 12288
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 1397 12183 1455 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2958 12220 2964 12232
rect 2919 12192 2964 12220
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3344 12192 3648 12220
rect 1578 12112 1584 12164
rect 1636 12152 1642 12164
rect 2314 12152 2320 12164
rect 1636 12124 2320 12152
rect 1636 12112 1642 12124
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 2682 12152 2688 12164
rect 2643 12124 2688 12152
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 3344 12152 3372 12192
rect 2792 12124 3372 12152
rect 3620 12152 3648 12192
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4111 12223 4169 12229
rect 4111 12220 4123 12223
rect 3752 12192 4123 12220
rect 3752 12180 3758 12192
rect 4111 12189 4123 12192
rect 4157 12189 4169 12223
rect 4338 12220 4344 12232
rect 4299 12192 4344 12220
rect 4111 12183 4169 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4540 12229 4568 12260
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 3970 12152 3976 12164
rect 3620 12124 3976 12152
rect 2792 12096 2820 12124
rect 3970 12112 3976 12124
rect 4028 12152 4034 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 4028 12124 4261 12152
rect 4028 12112 4034 12124
rect 4249 12121 4261 12124
rect 4295 12152 4307 12155
rect 4890 12152 4896 12164
rect 4295 12124 4896 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 2774 12084 2780 12096
rect 2547 12056 2780 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 3660 12056 4629 12084
rect 3660 12044 3666 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 5000 12084 5028 12260
rect 5092 12229 5120 12328
rect 5258 12316 5264 12328
rect 5316 12356 5322 12368
rect 8205 12359 8263 12365
rect 8205 12356 8217 12359
rect 5316 12328 8217 12356
rect 5316 12316 5322 12328
rect 8205 12325 8217 12328
rect 8251 12325 8263 12359
rect 8205 12319 8263 12325
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 9490 12356 9496 12368
rect 8628 12328 9260 12356
rect 9451 12328 9496 12356
rect 8628 12316 8634 12328
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6880 12260 7389 12288
rect 6880 12248 6886 12260
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5718 12220 5724 12232
rect 5679 12192 5724 12220
rect 5077 12183 5135 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6961 12229 6989 12260
rect 7377 12257 7389 12260
rect 7423 12288 7435 12291
rect 7423 12260 8524 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7098 12229 7104 12232
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 6512 12192 6653 12220
rect 6512 12180 6518 12192
rect 6641 12189 6653 12192
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 6917 12223 6989 12229
rect 6917 12189 6929 12223
rect 6963 12192 6989 12223
rect 7061 12223 7104 12229
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7061 12189 7073 12223
rect 7061 12183 7104 12189
rect 7098 12180 7104 12183
rect 7156 12180 7162 12232
rect 8386 12229 8392 12232
rect 8384 12220 8392 12229
rect 8347 12192 8392 12220
rect 8384 12183 8392 12192
rect 8386 12180 8392 12183
rect 8444 12180 8450 12232
rect 8496 12229 8524 12260
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8736 12223 8794 12229
rect 8736 12189 8748 12223
rect 8782 12220 8794 12223
rect 8782 12214 8800 12220
rect 8846 12214 8852 12232
rect 8782 12189 8852 12214
rect 8736 12186 8852 12189
rect 8736 12183 8794 12186
rect 8846 12180 8852 12186
rect 8904 12180 8910 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9232 12220 9260 12328
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 10042 12356 10048 12368
rect 10003 12328 10048 12356
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10152 12356 10180 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 14366 12424 14372 12436
rect 12406 12396 14372 12424
rect 12406 12356 12434 12396
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 13262 12356 13268 12368
rect 10152 12328 12434 12356
rect 13223 12328 13268 12356
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9364 12260 9597 12288
rect 9364 12248 9370 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10594 12288 10600 12300
rect 10183 12260 10600 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 11848 12260 12020 12288
rect 11848 12248 11854 12260
rect 10965 12223 11023 12229
rect 9232 12192 10180 12220
rect 9125 12183 9183 12189
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 5684 12124 6009 12152
rect 5684 12112 5690 12124
rect 5997 12121 6009 12124
rect 6043 12121 6055 12155
rect 6362 12152 6368 12164
rect 6323 12124 6368 12152
rect 5997 12115 6055 12121
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 6546 12152 6552 12164
rect 6507 12124 6552 12152
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 6825 12155 6883 12161
rect 6825 12152 6837 12155
rect 6788 12124 6837 12152
rect 6788 12112 6794 12124
rect 6825 12121 6837 12124
rect 6871 12121 6883 12155
rect 7558 12152 7564 12164
rect 7519 12124 7564 12152
rect 6825 12115 6883 12121
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 7834 12152 7840 12164
rect 7668 12124 7840 12152
rect 7282 12084 7288 12096
rect 5000 12056 7288 12084
rect 4617 12047 4675 12053
rect 7282 12044 7288 12056
rect 7340 12084 7346 12096
rect 7668 12084 7696 12124
rect 7834 12112 7840 12124
rect 7892 12112 7898 12164
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8628 12124 8673 12152
rect 8628 12112 8634 12124
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 9674 12152 9680 12164
rect 8996 12124 9680 12152
rect 8996 12112 9002 12124
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 10152 12152 10180 12192
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 11606 12220 11612 12232
rect 11567 12192 11612 12220
rect 10965 12183 11023 12189
rect 10229 12155 10287 12161
rect 10229 12152 10241 12155
rect 10152 12124 10241 12152
rect 10229 12121 10241 12124
rect 10275 12121 10287 12155
rect 10229 12115 10287 12121
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10560 12124 10793 12152
rect 10560 12112 10566 12124
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10980 12152 11008 12183
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11992 12229 12020 12260
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 11977 12183 12035 12189
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 11238 12152 11244 12164
rect 10980 12124 11244 12152
rect 10781 12115 10839 12121
rect 11238 12112 11244 12124
rect 11296 12152 11302 12164
rect 12066 12152 12072 12164
rect 11296 12124 12072 12152
rect 11296 12112 11302 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 7340 12056 7696 12084
rect 7340 12044 7346 12056
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 7929 12087 7987 12093
rect 7800 12056 7845 12084
rect 7800 12044 7806 12056
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 9030 12084 9036 12096
rect 7975 12056 9036 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 10042 12084 10048 12096
rect 9548 12056 10048 12084
rect 9548 12044 9554 12056
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 10376 12056 10425 12084
rect 10376 12044 10382 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10413 12047 10471 12053
rect 10597 12087 10655 12093
rect 10597 12053 10609 12087
rect 10643 12084 10655 12087
rect 10962 12084 10968 12096
rect 10643 12056 10968 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 2958 11880 2964 11892
rect 2792 11852 2964 11880
rect 2222 11812 2228 11824
rect 2183 11784 2228 11812
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 2314 11772 2320 11824
rect 2372 11812 2378 11824
rect 2372 11784 2417 11812
rect 2372 11772 2378 11784
rect 2498 11744 2504 11756
rect 2459 11716 2504 11744
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2792 11753 2820 11852
rect 2958 11840 2964 11852
rect 3016 11880 3022 11892
rect 3016 11852 5396 11880
rect 3016 11840 3022 11852
rect 3513 11815 3571 11821
rect 3513 11781 3525 11815
rect 3559 11812 3571 11815
rect 3602 11812 3608 11824
rect 3559 11784 3608 11812
rect 3559 11781 3571 11784
rect 3513 11775 3571 11781
rect 3602 11772 3608 11784
rect 3660 11772 3666 11824
rect 4525 11815 4583 11821
rect 4525 11781 4537 11815
rect 4571 11812 4583 11815
rect 4798 11812 4804 11824
rect 4571 11784 4804 11812
rect 4571 11781 4583 11784
rect 4525 11775 4583 11781
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2866 11704 2872 11756
rect 2924 11744 2930 11756
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 2924 11716 3709 11744
rect 2924 11704 2930 11716
rect 3436 11688 3464 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4154 11744 4160 11756
rect 3835 11716 4160 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4724 11716 4905 11744
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11676 4399 11679
rect 4614 11676 4620 11688
rect 4387 11648 4620 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4724 11620 4752 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5368 11744 5396 11852
rect 5902 11840 5908 11892
rect 5960 11840 5966 11892
rect 6362 11840 6368 11892
rect 6420 11880 6426 11892
rect 6914 11880 6920 11892
rect 6420 11852 6592 11880
rect 6875 11852 6920 11880
rect 6420 11840 6426 11852
rect 5445 11815 5503 11821
rect 5445 11781 5457 11815
rect 5491 11812 5503 11815
rect 5626 11812 5632 11824
rect 5491 11784 5632 11812
rect 5491 11781 5503 11784
rect 5445 11775 5503 11781
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 5920 11775 5948 11840
rect 6564 11824 6592 11852
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 9217 11883 9275 11889
rect 7392 11852 7967 11880
rect 6546 11812 6552 11824
rect 6012 11784 6408 11812
rect 6507 11784 6552 11812
rect 5904 11769 5962 11775
rect 5368 11716 5488 11744
rect 5261 11707 5319 11713
rect 5276 11676 5304 11707
rect 4816 11648 5304 11676
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2682 11608 2688 11620
rect 2179 11580 2688 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11577 4307 11611
rect 4706 11608 4712 11620
rect 4667 11580 4712 11608
rect 4249 11571 4307 11577
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 2774 11540 2780 11552
rect 1627 11512 2780 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 4264 11540 4292 11571
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 4816 11552 4844 11648
rect 5460 11608 5488 11716
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5592 11716 5637 11744
rect 5592 11704 5598 11716
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 5812 11747 5870 11753
rect 5812 11744 5824 11747
rect 5776 11716 5824 11744
rect 5776 11704 5782 11716
rect 5812 11713 5824 11716
rect 5858 11713 5870 11747
rect 5904 11735 5916 11769
rect 5950 11735 5962 11769
rect 6012 11756 6040 11784
rect 5904 11729 5962 11735
rect 5812 11707 5870 11713
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6052 11716 6097 11744
rect 6052 11704 6058 11716
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6380 11753 6408 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 7282 11778 7288 11824
rect 7225 11772 7288 11778
rect 7340 11772 7346 11824
rect 6365 11747 6423 11753
rect 6236 11716 6281 11744
rect 6236 11704 6242 11716
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 7098 11744 7104 11756
rect 6411 11716 7104 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7225 11753 7328 11772
rect 7193 11750 7328 11753
rect 7193 11747 7253 11750
rect 7193 11713 7205 11747
rect 7239 11716 7253 11747
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 5552 11676 5580 11704
rect 7392 11676 7420 11852
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 7939 11812 7967 11852
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 10686 11880 10692 11892
rect 9263 11852 10692 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 11606 11880 11612 11892
rect 10796 11852 11008 11880
rect 11567 11852 11612 11880
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 7800 11784 7845 11812
rect 7939 11784 10149 11812
rect 7800 11772 7806 11784
rect 10137 11781 10149 11784
rect 10183 11781 10195 11815
rect 10137 11775 10195 11781
rect 10321 11815 10379 11821
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 10502 11812 10508 11824
rect 10367 11784 10508 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10796 11812 10824 11852
rect 10980 11821 11008 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 10612 11784 10824 11812
rect 10965 11815 11023 11821
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8018 11744 8024 11756
rect 7975 11716 8024 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8251 11716 8432 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 5552 11648 7420 11676
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 8128 11676 8156 11707
rect 7469 11639 7527 11645
rect 8036 11648 8156 11676
rect 8297 11679 8355 11685
rect 6546 11608 6552 11620
rect 5460 11580 6552 11608
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 7484 11608 7512 11639
rect 7248 11580 7512 11608
rect 7248 11568 7254 11580
rect 4798 11540 4804 11552
rect 4264 11512 4804 11540
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6641 11543 6699 11549
rect 6641 11540 6653 11543
rect 6512 11512 6653 11540
rect 6512 11500 6518 11512
rect 6641 11509 6653 11512
rect 6687 11540 6699 11543
rect 7282 11540 7288 11552
rect 6687 11512 7288 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 7558 11540 7564 11552
rect 7423 11512 7564 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 7558 11500 7564 11512
rect 7616 11540 7622 11552
rect 8036 11540 8064 11648
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 8312 11608 8340 11639
rect 8404 11620 8432 11716
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 8536 11716 8585 11744
rect 8536 11704 8542 11716
rect 8573 11713 8585 11716
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 8754 11744 8760 11756
rect 8711 11716 8760 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 8588 11676 8616 11707
rect 8754 11704 8760 11716
rect 8812 11744 8818 11756
rect 8938 11744 8944 11756
rect 8812 11716 8944 11744
rect 8812 11704 8818 11716
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9309 11747 9367 11753
rect 9309 11713 9321 11747
rect 9355 11744 9367 11747
rect 9674 11744 9680 11756
rect 9355 11716 9536 11744
rect 9635 11716 9680 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 9398 11676 9404 11688
rect 8588 11648 9404 11676
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 8168 11580 8340 11608
rect 8168 11568 8174 11580
rect 8202 11540 8208 11552
rect 7616 11512 8208 11540
rect 7616 11500 7622 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8312 11540 8340 11580
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 8444 11580 8489 11608
rect 8444 11568 8450 11580
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9508 11608 9536 11716
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 9824 11716 9869 11744
rect 9824 11704 9830 11716
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10612 11744 10640 11784
rect 10965 11781 10977 11815
rect 11011 11812 11023 11815
rect 11146 11812 11152 11824
rect 11011 11784 11152 11812
rect 11011 11781 11023 11784
rect 10965 11775 11023 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 12989 11815 13047 11821
rect 12989 11812 13001 11815
rect 11480 11784 13001 11812
rect 11480 11772 11486 11784
rect 12989 11781 13001 11784
rect 13035 11781 13047 11815
rect 13262 11812 13268 11824
rect 13223 11784 13268 11812
rect 12989 11775 13047 11781
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 10100 11716 10640 11744
rect 10100 11704 10106 11716
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 10870 11753 10876 11756
rect 10827 11747 10876 11753
rect 10744 11716 10789 11744
rect 10744 11704 10750 11716
rect 10827 11713 10839 11747
rect 10873 11713 10876 11747
rect 10827 11707 10876 11713
rect 10870 11704 10876 11707
rect 10928 11704 10934 11756
rect 11062 11747 11120 11753
rect 11062 11713 11074 11747
rect 11108 11744 11120 11747
rect 11330 11744 11336 11756
rect 11108 11716 11336 11744
rect 11108 11713 11120 11716
rect 11062 11707 11120 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11440 11716 11529 11744
rect 9692 11676 9720 11704
rect 10502 11676 10508 11688
rect 9692 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10410 11608 10416 11620
rect 8996 11580 9260 11608
rect 9508 11580 10416 11608
rect 8996 11568 9002 11580
rect 8754 11540 8760 11552
rect 8312 11512 8760 11540
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9122 11540 9128 11552
rect 8895 11512 9128 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9232 11540 9260 11580
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 11440 11608 11468 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11698 11704 11704 11756
rect 11756 11753 11762 11756
rect 11756 11747 11783 11753
rect 11771 11713 11783 11747
rect 11756 11707 11783 11713
rect 11756 11704 11762 11707
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12124 11716 12169 11744
rect 12124 11704 12130 11716
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12860 11716 12909 11744
rect 12860 11704 12866 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 11809 11679 11867 11685
rect 11809 11676 11821 11679
rect 11808 11645 11821 11676
rect 11855 11645 11867 11679
rect 11808 11639 11867 11645
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12710 11676 12716 11688
rect 12483 11648 12716 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 11514 11608 11520 11620
rect 10520 11580 11520 11608
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 9232 11512 9505 11540
rect 9493 11509 9505 11512
rect 9539 11509 9551 11543
rect 9493 11503 9551 11509
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10318 11540 10324 11552
rect 9999 11512 10324 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10520 11549 10548 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 11808 11608 11836 11639
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 11974 11608 11980 11620
rect 11808 11580 11980 11608
rect 11974 11568 11980 11580
rect 12032 11568 12038 11620
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11509 10563 11543
rect 11238 11540 11244 11552
rect 11199 11512 11244 11540
rect 10505 11503 10563 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 11388 11512 12081 11540
rect 11388 11500 11394 11512
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 12069 11503 12127 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 6822 11336 6828 11348
rect 5767 11308 6828 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 8018 11336 8024 11348
rect 7156 11308 8024 11336
rect 7156 11296 7162 11308
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8113 11339 8171 11345
rect 8113 11305 8125 11339
rect 8159 11336 8171 11339
rect 8159 11308 9076 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 2682 11268 2688 11280
rect 2643 11240 2688 11268
rect 2682 11228 2688 11240
rect 2740 11228 2746 11280
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 5077 11271 5135 11277
rect 5077 11268 5089 11271
rect 4856 11240 5089 11268
rect 4856 11228 4862 11240
rect 5077 11237 5089 11240
rect 5123 11237 5135 11271
rect 7006 11268 7012 11280
rect 5077 11231 5135 11237
rect 6288 11240 7012 11268
rect 1670 11200 1676 11212
rect 1412 11172 1676 11200
rect 1412 11141 1440 11172
rect 1670 11160 1676 11172
rect 1728 11200 1734 11212
rect 3513 11203 3571 11209
rect 3513 11200 3525 11203
rect 1728 11172 3525 11200
rect 1728 11160 1734 11172
rect 3513 11169 3525 11172
rect 3559 11169 3571 11203
rect 6178 11200 6184 11212
rect 3513 11163 3571 11169
rect 3712 11172 6184 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 1397 11095 1455 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 3292 11104 3341 11132
rect 3292 11092 3298 11104
rect 3329 11101 3341 11104
rect 3375 11132 3387 11135
rect 3712 11132 3740 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6288 11209 6316 11240
rect 7006 11228 7012 11240
rect 7064 11268 7070 11280
rect 7064 11240 7236 11268
rect 7064 11228 7070 11240
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 7098 11160 7104 11212
rect 7156 11160 7162 11212
rect 3375 11104 3740 11132
rect 3789 11135 3847 11141
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 3789 11101 3801 11135
rect 3835 11132 3847 11135
rect 4062 11132 4068 11144
rect 3835 11104 4068 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4706 11132 4712 11144
rect 4304 11104 4712 11132
rect 4304 11092 4310 11104
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5442 11132 5448 11144
rect 5224 11104 5448 11132
rect 5224 11092 5230 11104
rect 5442 11092 5448 11104
rect 5500 11132 5506 11144
rect 5951 11135 6009 11141
rect 5951 11132 5963 11135
rect 5500 11104 5963 11132
rect 5500 11092 5506 11104
rect 5951 11101 5963 11104
rect 5997 11101 6009 11135
rect 6454 11132 6460 11144
rect 6415 11104 6460 11132
rect 5951 11095 6009 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6604 11104 6653 11132
rect 6604 11092 6610 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6859 11135 6917 11141
rect 6859 11101 6871 11135
rect 6905 11132 6917 11135
rect 7116 11132 7144 11160
rect 7208 11141 7236 11240
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8297 11271 8355 11277
rect 8297 11268 8309 11271
rect 7892 11240 8309 11268
rect 7892 11228 7898 11240
rect 8297 11237 8309 11240
rect 8343 11237 8355 11271
rect 9048 11268 9076 11308
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 10134 11336 10140 11348
rect 9180 11308 9225 11336
rect 9324 11308 10140 11336
rect 9180 11296 9186 11308
rect 9324 11268 9352 11308
rect 10134 11296 10140 11308
rect 10192 11336 10198 11348
rect 10413 11339 10471 11345
rect 10413 11336 10425 11339
rect 10192 11308 10425 11336
rect 10192 11296 10198 11308
rect 10413 11305 10425 11308
rect 10459 11305 10471 11339
rect 10413 11299 10471 11305
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10744 11308 10793 11336
rect 10744 11296 10750 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11146 11336 11152 11348
rect 10928 11308 11152 11336
rect 10928 11296 10934 11308
rect 11146 11296 11152 11308
rect 11204 11336 11210 11348
rect 12066 11336 12072 11348
rect 11204 11308 12072 11336
rect 11204 11296 11210 11308
rect 9048 11240 9352 11268
rect 8297 11231 8355 11237
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 9858 11268 9864 11280
rect 9456 11240 9864 11268
rect 9456 11228 9462 11240
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 11606 11268 11612 11280
rect 11348 11240 11612 11268
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 8021 11203 8079 11209
rect 7340 11172 7420 11200
rect 7340 11160 7346 11172
rect 7392 11141 7420 11172
rect 7484 11172 7972 11200
rect 7484 11141 7512 11172
rect 7944 11141 7972 11172
rect 8021 11169 8033 11203
rect 8067 11200 8079 11203
rect 8110 11200 8116 11212
rect 8067 11172 8116 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 8260 11172 9965 11200
rect 8260 11160 8266 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 11348 11200 11376 11240
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 11514 11200 11520 11212
rect 10367 11172 11376 11200
rect 11475 11172 11520 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 6905 11104 7144 11132
rect 7193 11135 7251 11141
rect 6905 11101 6917 11104
rect 6859 11095 6917 11101
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7378 11135 7436 11141
rect 7378 11101 7390 11135
rect 7424 11101 7436 11135
rect 7378 11095 7436 11101
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7595 11135 7653 11141
rect 7595 11101 7607 11135
rect 7641 11101 7653 11135
rect 7595 11095 7653 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9401 11095 9459 11101
rect 9508 11104 9597 11132
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 4948 11036 5733 11064
rect 4948 11024 4954 11036
rect 5721 11033 5733 11036
rect 5767 11033 5779 11067
rect 6748 11064 6776 11095
rect 5721 11027 5779 11033
rect 6104 11036 6776 11064
rect 7101 11067 7159 11073
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3145 10999 3203 11005
rect 3145 10996 3157 10999
rect 3016 10968 3157 10996
rect 3016 10956 3022 10968
rect 3145 10965 3157 10968
rect 3191 10965 3203 10999
rect 3145 10959 3203 10965
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5994 10996 6000 11008
rect 5592 10968 6000 10996
rect 5592 10956 5598 10968
rect 5994 10956 6000 10968
rect 6052 10996 6058 11008
rect 6104 11005 6132 11036
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7282 11064 7288 11076
rect 7147 11036 7288 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 6052 10968 6101 10996
rect 6052 10956 6058 10968
rect 6089 10965 6101 10968
rect 6135 10965 6147 10999
rect 6089 10959 6147 10965
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7484 10996 7512 11095
rect 6972 10968 7512 10996
rect 7610 10996 7638 11095
rect 7837 11067 7895 11073
rect 7837 11033 7849 11067
rect 7883 11064 7895 11067
rect 8941 11067 8999 11073
rect 7883 11036 8800 11064
rect 7883 11033 7895 11036
rect 7837 11027 7895 11033
rect 7926 10996 7932 11008
rect 7610 10968 7932 10996
rect 6972 10956 6978 10968
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8168 10968 8585 10996
rect 8168 10956 8174 10968
rect 8573 10965 8585 10968
rect 8619 10996 8631 10999
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 8619 10968 8677 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 8665 10965 8677 10968
rect 8711 10965 8723 10999
rect 8772 10996 8800 11036
rect 8941 11033 8953 11067
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 8956 10996 8984 11027
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 9088 11036 9137 11064
rect 9088 11024 9094 11036
rect 9125 11033 9137 11036
rect 9171 11033 9183 11067
rect 9125 11027 9183 11033
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 9416 11064 9444 11095
rect 9508 11076 9536 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 9766 11132 9772 11144
rect 9727 11104 9772 11132
rect 9585 11095 9643 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 9916 11104 9961 11132
rect 9916 11092 9922 11104
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 10100 11104 10149 11132
rect 10100 11092 10106 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10778 11132 10784 11144
rect 10643 11104 10784 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 9272 11036 9444 11064
rect 9272 11024 9278 11036
rect 9490 11024 9496 11076
rect 9548 11024 9554 11076
rect 9784 11064 9812 11092
rect 10428 11064 10456 11095
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 11146 11132 11152 11144
rect 11107 11104 11152 11132
rect 10965 11095 11023 11101
rect 10980 11064 11008 11095
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11422 11132 11428 11144
rect 11383 11104 11428 11132
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11624 11141 11652 11228
rect 11992 11144 12020 11308
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12710 11336 12716 11348
rect 12207 11308 12716 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 11790 11141 11796 11144
rect 11624 11135 11691 11141
rect 11624 11104 11645 11135
rect 11633 11101 11645 11104
rect 11679 11101 11691 11135
rect 11633 11095 11691 11101
rect 11747 11135 11796 11141
rect 11747 11101 11759 11135
rect 11793 11101 11796 11135
rect 11747 11095 11796 11101
rect 11790 11092 11796 11095
rect 11848 11092 11854 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12360 11141 12388 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12345 11135 12403 11141
rect 12032 11104 12125 11132
rect 12032 11092 12038 11104
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12860 11104 13001 11132
rect 12860 11092 12866 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 9784 11036 10456 11064
rect 10520 11036 11008 11064
rect 8772 10968 8984 10996
rect 8665 10959 8723 10965
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 10042 10996 10048 11008
rect 9640 10968 10048 10996
rect 9640 10956 9646 10968
rect 10042 10956 10048 10968
rect 10100 10996 10106 11008
rect 10520 10996 10548 11036
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 12894 11064 12900 11076
rect 12492 11036 12900 11064
rect 12492 11024 12498 11036
rect 12894 11024 12900 11036
rect 12952 11064 12958 11076
rect 13265 11067 13323 11073
rect 13265 11064 13277 11067
rect 12952 11036 13277 11064
rect 12952 11024 12958 11036
rect 13265 11033 13277 11036
rect 13311 11033 13323 11067
rect 13265 11027 13323 11033
rect 10100 10968 10548 10996
rect 10100 10956 10106 10968
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11241 10999 11299 11005
rect 11241 10996 11253 10999
rect 11204 10968 11253 10996
rect 11204 10956 11210 10968
rect 11241 10965 11253 10968
rect 11287 10965 11299 10999
rect 11241 10959 11299 10965
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 12768 10968 13369 10996
rect 12768 10956 12774 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 13446 10956 13452 11008
rect 13504 10996 13510 11008
rect 13504 10968 13549 10996
rect 13504 10956 13510 10968
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3568 10764 3617 10792
rect 3568 10752 3574 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4614 10792 4620 10804
rect 4111 10764 4620 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 6181 10795 6239 10801
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6270 10792 6276 10804
rect 6227 10764 6276 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 10873 10795 10931 10801
rect 7668 10764 10364 10792
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 2593 10727 2651 10733
rect 2593 10724 2605 10727
rect 2556 10696 2605 10724
rect 2556 10684 2562 10696
rect 2593 10693 2605 10696
rect 2639 10693 2651 10727
rect 2593 10687 2651 10693
rect 3329 10727 3387 10733
rect 3329 10693 3341 10727
rect 3375 10724 3387 10727
rect 3694 10724 3700 10736
rect 3375 10696 3700 10724
rect 3375 10693 3387 10696
rect 3329 10687 3387 10693
rect 3694 10684 3700 10696
rect 3752 10684 3758 10736
rect 4246 10724 4252 10736
rect 4207 10696 4252 10724
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 5261 10727 5319 10733
rect 5261 10724 5273 10727
rect 5132 10696 5273 10724
rect 5132 10684 5138 10696
rect 5261 10693 5273 10696
rect 5307 10693 5319 10727
rect 7006 10724 7012 10736
rect 6967 10696 7012 10724
rect 5261 10687 5319 10693
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 7193 10727 7251 10733
rect 7193 10724 7205 10727
rect 7156 10696 7205 10724
rect 7156 10684 7162 10696
rect 7193 10693 7205 10696
rect 7239 10724 7251 10727
rect 7668 10724 7696 10764
rect 7926 10724 7932 10736
rect 7239 10696 7696 10724
rect 7839 10696 7932 10724
rect 7239 10693 7251 10696
rect 7193 10687 7251 10693
rect 1578 10616 1584 10668
rect 1636 10665 1642 10668
rect 1636 10659 1679 10665
rect 1667 10625 1679 10659
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1636 10619 1679 10625
rect 1636 10616 1642 10619
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2041 10659 2099 10665
rect 1912 10628 1957 10656
rect 1912 10616 1918 10628
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 3234 10656 3240 10668
rect 2087 10628 3240 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3418 10656 3424 10668
rect 3379 10628 3424 10656
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5215 10628 5856 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1504 10560 2145 10588
rect 1504 10529 1532 10560
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 3326 10588 3332 10600
rect 2731 10560 3332 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4172 10588 4200 10619
rect 4540 10588 4568 10619
rect 5828 10597 5856 10628
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 5960 10628 7389 10656
rect 5960 10616 5966 10628
rect 7377 10625 7389 10628
rect 7423 10656 7435 10659
rect 7558 10656 7564 10668
rect 7423 10628 7564 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 7668 10665 7696 10696
rect 7852 10665 7880 10696
rect 7926 10684 7932 10696
rect 7984 10724 7990 10736
rect 7984 10696 8156 10724
rect 7984 10684 7990 10696
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8128 10656 8156 10696
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 8260 10696 8401 10724
rect 8260 10684 8266 10696
rect 8389 10693 8401 10696
rect 8435 10724 8447 10727
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 8435 10696 8585 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 8754 10724 8760 10736
rect 8715 10696 8760 10724
rect 8573 10687 8631 10693
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9125 10727 9183 10733
rect 9125 10724 9137 10727
rect 9088 10696 9137 10724
rect 9088 10684 9094 10696
rect 9125 10693 9137 10696
rect 9171 10693 9183 10727
rect 9125 10687 9183 10693
rect 8941 10659 8999 10665
rect 8128 10628 8892 10656
rect 8021 10619 8079 10625
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 4172 10560 5365 10588
rect 5353 10557 5365 10560
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 6730 10588 6736 10600
rect 5859 10560 6736 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 8036 10588 8064 10619
rect 8754 10588 8760 10600
rect 6963 10560 7420 10588
rect 8036 10560 8760 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7392 10532 7420 10560
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 8864 10588 8892 10628
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9232 10656 9260 10764
rect 9766 10724 9772 10736
rect 9727 10696 9772 10724
rect 9766 10684 9772 10696
rect 9824 10724 9830 10736
rect 10229 10727 10287 10733
rect 10229 10724 10241 10727
rect 9824 10696 10241 10724
rect 9824 10684 9830 10696
rect 10229 10693 10241 10696
rect 10275 10693 10287 10727
rect 10229 10687 10287 10693
rect 9674 10656 9680 10668
rect 8987 10628 9260 10656
rect 9635 10628 9680 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 9950 10656 9956 10668
rect 9911 10628 9956 10656
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 9582 10588 9588 10600
rect 8864 10560 9588 10588
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 1578 10520 1584 10532
rect 1535 10492 1584 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 1578 10480 1584 10492
rect 1636 10480 1642 10532
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 6457 10523 6515 10529
rect 6457 10520 6469 10523
rect 6236 10492 6469 10520
rect 6236 10480 6242 10492
rect 6457 10489 6469 10492
rect 6503 10520 6515 10523
rect 6546 10520 6552 10532
rect 6503 10492 6552 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10489 6699 10523
rect 6641 10483 6699 10489
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10452 3022 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3016 10424 3801 10452
rect 3016 10412 3022 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5718 10452 5724 10464
rect 5132 10424 5724 10452
rect 5132 10412 5138 10424
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6362 10452 6368 10464
rect 6043 10424 6368 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6656 10452 6684 10483
rect 7374 10480 7380 10532
rect 7432 10480 7438 10532
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 7653 10523 7711 10529
rect 7653 10520 7665 10523
rect 7616 10492 7665 10520
rect 7616 10480 7622 10492
rect 7653 10489 7665 10492
rect 7699 10489 7711 10523
rect 10152 10520 10180 10619
rect 10336 10588 10364 10764
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11330 10792 11336 10804
rect 10919 10764 11336 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11514 10752 11520 10804
rect 11572 10752 11578 10804
rect 11974 10792 11980 10804
rect 11808 10764 11980 10792
rect 11532 10724 11560 10752
rect 11808 10733 11836 10764
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 10704 10696 11560 10724
rect 11793 10727 11851 10733
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 10704 10665 10732 10696
rect 11793 10693 11805 10727
rect 11839 10693 11851 10727
rect 12710 10724 12716 10736
rect 12671 10696 12716 10724
rect 11793 10687 11851 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 13446 10724 13452 10736
rect 13407 10696 13452 10724
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 10689 10659 10747 10665
rect 10468 10628 10513 10656
rect 10468 10616 10474 10628
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 11146 10656 11152 10668
rect 11107 10628 11152 10656
rect 10689 10619 10747 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11330 10656 11336 10668
rect 11291 10628 11336 10656
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11164 10588 11192 10616
rect 10336 10560 11192 10588
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11532 10588 11560 10619
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11664 10628 11713 10656
rect 11664 10616 11670 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11937 10659 11995 10665
rect 11937 10625 11949 10659
rect 11983 10656 11995 10659
rect 13170 10656 13176 10668
rect 11983 10628 13176 10656
rect 11983 10625 11995 10628
rect 11937 10619 11995 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 11296 10560 11560 10588
rect 11296 10548 11302 10560
rect 12066 10548 12072 10600
rect 12124 10588 12130 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 12124 10560 12265 10588
rect 12124 10548 12130 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12253 10551 12311 10557
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 12952 10560 12997 10588
rect 12952 10548 12958 10560
rect 10318 10520 10324 10532
rect 10152 10492 10324 10520
rect 7653 10483 7711 10489
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10594 10520 10600 10532
rect 10555 10492 10600 10520
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10704 10492 12112 10520
rect 6914 10452 6920 10464
rect 6656 10424 6920 10452
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9122 10452 9128 10464
rect 8904 10424 9128 10452
rect 8904 10412 8910 10424
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 9180 10424 9321 10452
rect 9180 10412 9186 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9309 10415 9367 10421
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9456 10424 9505 10452
rect 9456 10412 9462 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10704 10452 10732 10492
rect 9640 10424 10732 10452
rect 11057 10455 11115 10461
rect 9640 10412 9646 10424
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11698 10452 11704 10464
rect 11103 10424 11704 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12084 10461 12112 10492
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 13357 10523 13415 10529
rect 13357 10520 13369 10523
rect 13320 10492 13369 10520
rect 13320 10480 13326 10492
rect 13357 10489 13369 10492
rect 13403 10489 13415 10523
rect 13357 10483 13415 10489
rect 12069 10455 12127 10461
rect 12069 10421 12081 10455
rect 12115 10421 12127 10455
rect 12069 10415 12127 10421
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 1489 10251 1547 10257
rect 1489 10217 1501 10251
rect 1535 10248 1547 10251
rect 1762 10248 1768 10260
rect 1535 10220 1768 10248
rect 1535 10217 1547 10220
rect 1489 10211 1547 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 3326 10248 3332 10260
rect 3287 10220 3332 10248
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 3786 10248 3792 10260
rect 3651 10220 3792 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 5442 10248 5448 10260
rect 4019 10220 5448 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5592 10220 5641 10248
rect 5592 10208 5598 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 7282 10248 7288 10260
rect 6503 10220 7288 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7432 10220 7477 10248
rect 7432 10208 7438 10220
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 7708 10220 8401 10248
rect 7708 10208 7714 10220
rect 8389 10217 8401 10220
rect 8435 10217 8447 10251
rect 8389 10211 8447 10217
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8536 10220 8585 10248
rect 8536 10208 8542 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 10410 10248 10416 10260
rect 9088 10220 10416 10248
rect 9088 10208 9094 10220
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 11149 10251 11207 10257
rect 11149 10217 11161 10251
rect 11195 10248 11207 10251
rect 11330 10248 11336 10260
rect 11195 10220 11336 10248
rect 11195 10217 11207 10220
rect 11149 10211 11207 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11480 10220 11805 10248
rect 11480 10208 11486 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 2869 10183 2927 10189
rect 2869 10180 2881 10183
rect 2556 10152 2881 10180
rect 2556 10140 2562 10152
rect 2869 10149 2881 10152
rect 2915 10149 2927 10183
rect 2869 10143 2927 10149
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 6825 10183 6883 10189
rect 5040 10152 6224 10180
rect 5040 10140 5046 10152
rect 1854 10072 1860 10124
rect 1912 10112 1918 10124
rect 4617 10115 4675 10121
rect 1912 10084 4568 10112
rect 1912 10072 1918 10084
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3142 10044 3148 10056
rect 3099 10016 3148 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3660 10016 4077 10044
rect 3660 10004 3666 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4540 10044 4568 10084
rect 4617 10081 4629 10115
rect 4663 10112 4675 10115
rect 6086 10112 6092 10124
rect 4663 10084 6092 10112
rect 4663 10081 4675 10084
rect 4617 10075 4675 10081
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6196 10112 6224 10152
rect 6825 10149 6837 10183
rect 6871 10180 6883 10183
rect 7098 10180 7104 10192
rect 6871 10152 7104 10180
rect 6871 10149 6883 10152
rect 6825 10143 6883 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7193 10183 7251 10189
rect 7193 10149 7205 10183
rect 7239 10180 7251 10183
rect 13262 10180 13268 10192
rect 7239 10152 12020 10180
rect 13223 10152 13268 10180
rect 7239 10149 7251 10152
rect 7193 10143 7251 10149
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 6196 10084 6776 10112
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4540 10016 4905 10044
rect 4065 10007 4123 10013
rect 4893 10013 4905 10016
rect 4939 10044 4951 10047
rect 5261 10047 5319 10053
rect 4939 10016 5212 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 4522 9976 4528 9988
rect 4483 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5074 9976 5080 9988
rect 5035 9948 5080 9976
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5184 9976 5212 10016
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5307 10016 5917 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6270 10004 6276 10056
rect 6328 10053 6334 10056
rect 6748 10053 6776 10084
rect 7760 10084 9045 10112
rect 6328 10044 6336 10053
rect 6733 10047 6791 10053
rect 6328 10016 6373 10044
rect 6328 10007 6336 10016
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6733 10007 6791 10013
rect 6328 10004 6334 10007
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7374 10044 7380 10056
rect 7055 10016 7380 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 5534 9976 5540 9988
rect 5184 9948 5540 9976
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 5810 9976 5816 9988
rect 5771 9948 5816 9976
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 5994 9936 6000 9988
rect 6052 9976 6058 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 6052 9948 6101 9976
rect 6052 9936 6058 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 6362 9976 6368 9988
rect 6227 9948 6368 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 6362 9936 6368 9948
rect 6420 9976 6426 9988
rect 6420 9948 6776 9976
rect 6420 9936 6426 9948
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4709 9911 4767 9917
rect 4709 9908 4721 9911
rect 3844 9880 4721 9908
rect 3844 9868 3850 9880
rect 4709 9877 4721 9880
rect 4755 9877 4767 9911
rect 4709 9871 4767 9877
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5408 9880 5457 9908
rect 5408 9868 5414 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 6012 9908 6040 9936
rect 6748 9920 6776 9948
rect 5675 9880 6040 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 7024 9908 7052 10007
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7760 10053 7788 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9950 10072 9956 10124
rect 10008 10072 10014 10124
rect 10226 10121 10232 10124
rect 10212 10115 10232 10121
rect 10212 10081 10224 10115
rect 10212 10075 10232 10081
rect 10226 10072 10232 10075
rect 10284 10072 10290 10124
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10686 10112 10692 10124
rect 10551 10084 10692 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 10836 10084 11744 10112
rect 10836 10072 10842 10084
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 6788 9880 7052 9908
rect 7852 9908 7880 10007
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 7984 10016 8677 10044
rect 7984 10004 7990 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 8938 10044 8944 10056
rect 8803 10016 8944 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9214 10044 9220 10056
rect 9175 10016 9220 10044
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9398 10044 9404 10056
rect 9355 10016 9404 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 8205 9979 8263 9985
rect 8205 9945 8217 9979
rect 8251 9976 8263 9979
rect 8570 9976 8576 9988
rect 8251 9948 8576 9976
rect 8251 9945 8263 9948
rect 8205 9939 8263 9945
rect 8570 9936 8576 9948
rect 8628 9936 8634 9988
rect 8956 9976 8984 10004
rect 9508 9976 9536 10007
rect 9582 10004 9588 10056
rect 9640 10044 9646 10056
rect 9968 10044 9996 10072
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 9640 10016 10609 10044
rect 9640 10004 9646 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10870 10044 10876 10056
rect 10831 10016 10876 10044
rect 10597 10007 10655 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 9766 9976 9772 9988
rect 8956 9948 9536 9976
rect 9727 9948 9772 9976
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 9950 9976 9956 9988
rect 9911 9948 9956 9976
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 11072 9976 11100 10007
rect 10152 9948 11100 9976
rect 11256 9976 11284 10007
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11388 10016 11529 10044
rect 11388 10004 11394 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 11716 9988 11744 10084
rect 11992 10053 12020 10152
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12894 10044 12900 10056
rect 12023 10016 12900 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 11422 9976 11428 9988
rect 11256 9948 11428 9976
rect 8478 9908 8484 9920
rect 7852 9880 8484 9908
rect 6788 9868 6794 9880
rect 8478 9868 8484 9880
rect 8536 9908 8542 9920
rect 9306 9908 9312 9920
rect 8536 9880 9312 9908
rect 8536 9868 8542 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10152 9908 10180 9948
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 11698 9976 11704 9988
rect 11659 9948 11704 9976
rect 11698 9936 11704 9948
rect 11756 9936 11762 9988
rect 10318 9908 10324 9920
rect 9548 9880 10180 9908
rect 10279 9880 10324 9908
rect 9548 9868 9554 9880
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10459 9880 10885 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10873 9877 10885 9880
rect 10919 9908 10931 9911
rect 11146 9908 11152 9920
rect 10919 9880 11152 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 1486 9704 1492 9716
rect 1447 9676 1492 9704
rect 1486 9664 1492 9676
rect 1544 9664 1550 9716
rect 2884 9676 3372 9704
rect 2884 9636 2912 9676
rect 2148 9608 2912 9636
rect 2961 9639 3019 9645
rect 2148 9577 2176 9608
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 3234 9636 3240 9648
rect 3007 9608 3240 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 3344 9636 3372 9676
rect 5350 9664 5356 9716
rect 5408 9664 5414 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 5776 9676 6960 9704
rect 5776 9664 5782 9676
rect 4798 9636 4804 9648
rect 3344 9608 4804 9636
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 5368 9636 5396 9664
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 5368 9608 6837 9636
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6932 9636 6960 9676
rect 7760 9676 8340 9704
rect 6932 9608 7328 9636
rect 6825 9599 6883 9605
rect 7300 9580 7328 9608
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2406 9568 2412 9580
rect 2271 9540 2412 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9568 3206 9580
rect 3421 9571 3479 9577
rect 3200 9540 3280 9568
rect 3200 9528 3206 9540
rect 3252 9509 3280 9540
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3421 9531 3479 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9469 3295 9503
rect 3436 9500 3464 9531
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5123 9540 5273 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5261 9537 5273 9540
rect 5307 9568 5319 9571
rect 5350 9568 5356 9580
rect 5307 9540 5356 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 3436 9472 4568 9500
rect 3237 9463 3295 9469
rect 4540 9444 4568 9472
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 6196 9500 6224 9531
rect 6546 9528 6552 9580
rect 6604 9577 6610 9580
rect 6604 9571 6647 9577
rect 6635 9537 6647 9571
rect 6604 9531 6647 9537
rect 6604 9528 6610 9531
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7009 9571 7067 9577
rect 6788 9540 6833 9568
rect 6788 9528 6794 9540
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 7055 9540 7113 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 7101 9531 7159 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7760 9568 7788 9676
rect 7834 9596 7840 9648
rect 7892 9636 7898 9648
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 7892 9608 8125 9636
rect 7892 9596 7898 9608
rect 8113 9605 8125 9608
rect 8159 9605 8171 9639
rect 8312 9636 8340 9676
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 9490 9704 9496 9716
rect 8812 9676 9496 9704
rect 8812 9664 8818 9676
rect 9490 9664 9496 9676
rect 9548 9704 9554 9716
rect 9548 9676 9812 9704
rect 9548 9664 9554 9676
rect 8846 9636 8852 9648
rect 8312 9608 8852 9636
rect 8113 9599 8171 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 9784 9645 9812 9676
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10870 9704 10876 9716
rect 10008 9676 10876 9704
rect 10008 9664 10014 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11422 9704 11428 9716
rect 11164 9676 11428 9704
rect 9769 9639 9827 9645
rect 8956 9608 9444 9636
rect 7515 9540 7788 9568
rect 7924 9571 7982 9577
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7924 9537 7936 9571
rect 7970 9537 7982 9571
rect 7924 9531 7982 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8202 9568 8208 9580
rect 8067 9540 8208 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 7944 9500 7972 9531
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8570 9568 8576 9580
rect 8343 9540 8576 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8754 9568 8760 9580
rect 8715 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 8956 9577 8984 9608
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 9122 9568 9128 9580
rect 9083 9540 9128 9568
rect 8941 9531 8999 9537
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9416 9577 9444 9608
rect 9769 9605 9781 9639
rect 9815 9605 9827 9639
rect 10505 9639 10563 9645
rect 10505 9636 10517 9639
rect 9769 9599 9827 9605
rect 10060 9608 10517 9636
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 9582 9568 9588 9580
rect 9447 9540 9588 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 9732 9540 9873 9568
rect 9732 9528 9738 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10060 9577 10088 9608
rect 10505 9605 10517 9608
rect 10551 9605 10563 9639
rect 10686 9636 10692 9648
rect 10647 9608 10692 9636
rect 10505 9599 10563 9605
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 10008 9540 10057 9568
rect 10008 9528 10014 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10410 9568 10416 9580
rect 10367 9540 10416 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 8662 9500 8668 9512
rect 5224 9472 6679 9500
rect 7944 9472 8668 9500
rect 5224 9460 5230 9472
rect 1670 9432 1676 9444
rect 1583 9404 1676 9432
rect 1670 9392 1676 9404
rect 1728 9432 1734 9444
rect 2958 9432 2964 9444
rect 1728 9404 2964 9432
rect 1728 9392 1734 9404
rect 2958 9392 2964 9404
rect 3016 9432 3022 9444
rect 3786 9432 3792 9444
rect 3016 9404 3792 9432
rect 3016 9392 3022 9404
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4580 9404 4905 9432
rect 4580 9392 4586 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 6651 9432 6679 9472
rect 8496 9441 8524 9472
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 9214 9500 9220 9512
rect 9175 9472 9220 9500
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9766 9500 9772 9512
rect 9324 9472 9772 9500
rect 7745 9435 7803 9441
rect 7745 9432 7757 9435
rect 4893 9395 4951 9401
rect 6288 9404 6592 9432
rect 6651 9404 7757 9432
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 6288 9364 6316 9404
rect 6454 9364 6460 9376
rect 2464 9336 6316 9364
rect 6415 9336 6460 9364
rect 2464 9324 2470 9336
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6564 9364 6592 9404
rect 7745 9401 7757 9404
rect 7791 9401 7803 9435
rect 7745 9395 7803 9401
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9401 8539 9435
rect 9324 9432 9352 9472
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9674 9432 9680 9444
rect 8481 9395 8539 9401
rect 8680 9404 9352 9432
rect 9416 9404 9680 9432
rect 8680 9364 8708 9404
rect 6564 9336 8708 9364
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9416 9373 9444 9404
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10520 9432 10548 9599
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 11164 9577 11192 9676
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 12860 9676 13185 9704
rect 12860 9664 12866 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 13173 9667 13231 9673
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9537 11299 9571
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 11241 9531 11299 9537
rect 11256 9500 11284 9531
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 11698 9568 11704 9580
rect 11659 9540 11704 9568
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 11256 9472 11744 9500
rect 10520 9404 11008 9432
rect 9401 9367 9459 9373
rect 8812 9336 8857 9364
rect 8812 9324 8818 9336
rect 9401 9333 9413 9367
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 9585 9367 9643 9373
rect 9585 9333 9597 9367
rect 9631 9364 9643 9367
rect 10778 9364 10784 9376
rect 9631 9336 10784 9364
rect 9631 9333 9643 9336
rect 9585 9327 9643 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 10980 9364 11008 9404
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11716 9441 11744 9472
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 11112 9404 11253 9432
rect 11112 9392 11118 9404
rect 11241 9401 11253 9404
rect 11287 9401 11299 9435
rect 11241 9395 11299 9401
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 12084 9364 12112 9531
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12216 9540 12261 9568
rect 12216 9528 12222 9540
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 12768 9540 12817 9568
rect 12768 9528 12774 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13354 9568 13360 9580
rect 13127 9540 13360 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13538 9364 13544 9376
rect 10980 9336 12112 9364
rect 13499 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 1394 9160 1400 9172
rect 1355 9132 1400 9160
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 3326 9160 3332 9172
rect 3287 9132 3332 9160
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 3660 9132 4905 9160
rect 3660 9120 3666 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 6086 9160 6092 9172
rect 4893 9123 4951 9129
rect 5552 9132 5948 9160
rect 6047 9132 6092 9160
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 3234 9092 3240 9104
rect 2915 9064 3240 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 2406 9024 2412 9036
rect 2367 8996 2412 9024
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 3344 9024 3372 9120
rect 5552 9104 5580 9132
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 4249 9095 4307 9101
rect 4249 9092 4261 9095
rect 3568 9064 4261 9092
rect 3568 9052 3574 9064
rect 4249 9061 4261 9064
rect 4295 9061 4307 9095
rect 5534 9092 5540 9104
rect 5495 9064 5540 9092
rect 4249 9055 4307 9061
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 5721 9095 5779 9101
rect 5721 9092 5733 9095
rect 5644 9064 5733 9092
rect 5077 9027 5135 9033
rect 3344 8996 4476 9024
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 4448 8965 4476 8996
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 5166 9024 5172 9036
rect 5123 8996 5172 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5644 9033 5672 9064
rect 5721 9061 5733 9064
rect 5767 9061 5779 9095
rect 5721 9055 5779 9061
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5920 9024 5948 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 7742 9160 7748 9172
rect 6656 9132 7748 9160
rect 6656 9104 6684 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9309 9163 9367 9169
rect 8904 9132 9260 9160
rect 8904 9120 8910 9132
rect 6638 9092 6644 9104
rect 6564 9064 6644 9092
rect 5920 8996 6040 9024
rect 5629 8987 5687 8993
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3200 8928 3249 8956
rect 3200 8916 3206 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4433 8959 4491 8965
rect 4111 8928 4384 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 2961 8891 3019 8897
rect 2961 8857 2973 8891
rect 3007 8857 3019 8891
rect 2961 8851 3019 8857
rect 3605 8891 3663 8897
rect 3605 8857 3617 8891
rect 3651 8888 3663 8891
rect 3786 8888 3792 8900
rect 3651 8860 3792 8888
rect 3651 8857 3663 8860
rect 3605 8851 3663 8857
rect 2976 8820 3004 8851
rect 3786 8848 3792 8860
rect 3844 8888 3850 8900
rect 4356 8888 4384 8928
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5258 8956 5264 8968
rect 4755 8928 5264 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 6012 8965 6040 8996
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5408 8928 5917 8956
rect 5408 8916 5414 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6564 8956 6592 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 6972 9064 7481 9092
rect 6972 9052 6978 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 8018 9092 8024 9104
rect 7469 9055 7527 9061
rect 7576 9064 8024 9092
rect 6932 9024 6960 9052
rect 6656 8996 6960 9024
rect 6656 8965 6684 8996
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7576 9024 7604 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8754 9092 8760 9104
rect 8251 9064 8760 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 9030 9092 9036 9104
rect 8812 9064 9036 9092
rect 8812 9052 8818 9064
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9232 9092 9260 9132
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9674 9160 9680 9172
rect 9355 9132 9680 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 10134 9160 10140 9172
rect 9907 9132 10140 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 12066 9160 12072 9172
rect 11931 9132 12072 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 9398 9092 9404 9104
rect 9232 9064 9404 9092
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 9582 9092 9588 9104
rect 9543 9064 9588 9092
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 10042 9092 10048 9104
rect 9692 9064 10048 9092
rect 7926 9024 7932 9036
rect 7340 8996 7604 9024
rect 7668 8996 7932 9024
rect 7340 8984 7346 8996
rect 6503 8928 6592 8956
rect 6641 8959 6699 8965
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7006 8956 7012 8968
rect 6779 8928 7012 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7668 8965 7696 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8036 9024 8064 9052
rect 8481 9027 8539 9033
rect 8036 8996 8432 9024
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7653 8959 7711 8965
rect 7239 8928 7604 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 6825 8891 6883 8897
rect 6825 8888 6837 8891
rect 3844 8860 4292 8888
rect 4356 8860 6837 8888
rect 3844 8848 3850 8860
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2976 8792 3065 8820
rect 3053 8789 3065 8792
rect 3099 8789 3111 8823
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3053 8783 3111 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4264 8820 4292 8860
rect 6825 8857 6837 8860
rect 6871 8888 6883 8891
rect 7466 8888 7472 8900
rect 6871 8860 7472 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4264 8792 4537 8820
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6730 8820 6736 8832
rect 6420 8792 6736 8820
rect 6420 8780 6426 8792
rect 6730 8780 6736 8792
rect 6788 8820 6794 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6788 8792 7297 8820
rect 6788 8780 6794 8792
rect 7285 8789 7297 8792
rect 7331 8820 7343 8823
rect 7576 8820 7604 8928
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8404 8965 8432 8996
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 9692 9024 9720 9064
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 10505 9095 10563 9101
rect 10505 9092 10517 9095
rect 10468 9064 10517 9092
rect 10468 9052 10474 9064
rect 10505 9061 10517 9064
rect 10551 9061 10563 9095
rect 10505 9055 10563 9061
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 11330 9092 11336 9104
rect 10928 9064 11336 9092
rect 10928 9052 10934 9064
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 11609 9095 11667 9101
rect 11609 9061 11621 9095
rect 11655 9092 11667 9095
rect 11655 9064 12480 9092
rect 11655 9061 11667 9064
rect 11609 9055 11667 9061
rect 8527 8996 9720 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10744 8996 11100 9024
rect 10744 8984 10750 8996
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7800 8928 8033 8956
rect 7800 8916 7806 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8662 8956 8668 8968
rect 8435 8928 8668 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 7834 8888 7840 8900
rect 7795 8860 7840 8888
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 8312 8888 8340 8919
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8904 8928 8953 8956
rect 8904 8916 8910 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9398 8956 9404 8968
rect 9088 8928 9404 8956
rect 9088 8916 9094 8928
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9950 8956 9956 8968
rect 9732 8928 9777 8956
rect 9911 8928 9956 8956
rect 9732 8916 9738 8928
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10226 8916 10232 8968
rect 10284 8958 10290 8968
rect 11072 8965 11100 8996
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11204 8996 12112 9024
rect 11204 8984 11210 8996
rect 10413 8959 10471 8965
rect 10284 8956 10364 8958
rect 10284 8928 10377 8956
rect 10284 8916 10290 8928
rect 9122 8888 9128 8900
rect 8312 8860 9128 8888
rect 9122 8848 9128 8860
rect 9180 8888 9186 8900
rect 9858 8888 9864 8900
rect 9180 8860 9864 8888
rect 9180 8848 9186 8860
rect 9858 8848 9864 8860
rect 9916 8888 9922 8900
rect 10045 8891 10103 8897
rect 10045 8888 10057 8891
rect 9916 8860 10057 8888
rect 9916 8848 9922 8860
rect 10045 8857 10057 8860
rect 10091 8857 10103 8891
rect 10336 8888 10364 8928
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 11057 8959 11115 8965
rect 10459 8928 10916 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10888 8900 10916 8928
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 11057 8919 11115 8925
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11477 8959 11535 8965
rect 11477 8925 11489 8959
rect 11523 8956 11535 8959
rect 11974 8956 11980 8968
rect 11523 8928 11980 8956
rect 11523 8925 11535 8928
rect 11477 8919 11535 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12084 8965 12112 8996
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12452 9033 12480 9064
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 12400 8996 12449 9024
rect 12400 8984 12406 8996
rect 12437 8993 12449 8996
rect 12483 8993 12495 9027
rect 13538 9024 13544 9036
rect 12437 8987 12495 8993
rect 12636 8996 13544 9024
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 10689 8891 10747 8897
rect 10689 8888 10701 8891
rect 10336 8860 10701 8888
rect 10045 8851 10103 8857
rect 10689 8857 10701 8860
rect 10735 8857 10747 8891
rect 10870 8888 10876 8900
rect 10831 8860 10876 8888
rect 10689 8851 10747 8857
rect 8202 8820 8208 8832
rect 7331 8792 8208 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9306 8820 9312 8832
rect 9079 8792 9312 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 10594 8820 10600 8832
rect 9456 8792 10600 8820
rect 9456 8780 9462 8792
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10704 8820 10732 8851
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11241 8891 11299 8897
rect 11241 8888 11253 8891
rect 11020 8860 11253 8888
rect 11020 8848 11026 8860
rect 11241 8857 11253 8860
rect 11287 8857 11299 8891
rect 11348 8888 11376 8916
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 11348 8860 12265 8888
rect 11241 8851 11299 8857
rect 12253 8857 12265 8860
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 12345 8891 12403 8897
rect 12345 8857 12357 8891
rect 12391 8888 12403 8891
rect 12636 8888 12664 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 12894 8888 12900 8900
rect 12391 8860 12664 8888
rect 12855 8860 12900 8888
rect 12391 8857 12403 8860
rect 12345 8851 12403 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8857 13047 8891
rect 13446 8888 13452 8900
rect 13407 8860 13452 8888
rect 12989 8851 13047 8857
rect 11698 8820 11704 8832
rect 10704 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13004 8820 13032 8851
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 12492 8792 13032 8820
rect 12492 8780 12498 8792
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9916 8588 10057 8616
rect 9916 8576 9922 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10652 8588 11008 8616
rect 10652 8576 10658 8588
rect 4724 8520 5488 8548
rect 1486 8480 1492 8492
rect 1447 8452 1492 8480
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 4724 8489 4752 8520
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 4709 8443 4767 8449
rect 4816 8452 5273 8480
rect 4816 8356 4844 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5460 8480 5488 8520
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5592 8520 6009 8548
rect 5592 8508 5598 8520
rect 5997 8517 6009 8520
rect 6043 8517 6055 8551
rect 10134 8548 10140 8560
rect 5997 8511 6055 8517
rect 7944 8520 10140 8548
rect 5626 8480 5632 8492
rect 5460 8452 5632 8480
rect 5261 8443 5319 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6822 8480 6828 8492
rect 6783 8452 6828 8480
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7156 8452 7205 8480
rect 7156 8440 7162 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7558 8480 7564 8492
rect 7519 8452 7564 8480
rect 7193 8443 7251 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7944 8489 7972 8520
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10870 8548 10876 8560
rect 10284 8520 10876 8548
rect 10284 8508 10290 8520
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 9122 8480 9128 8492
rect 8619 8452 9128 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9640 8452 9873 8480
rect 9640 8440 9646 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10796 8489 10824 8520
rect 10870 8508 10876 8520
rect 10928 8508 10934 8560
rect 10980 8557 11008 8588
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11388 8588 11529 8616
rect 11388 8576 11394 8588
rect 11517 8585 11529 8588
rect 11563 8616 11575 8619
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 11563 8588 11713 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11701 8585 11713 8588
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12434 8616 12440 8628
rect 12299 8588 12440 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 10965 8551 11023 8557
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 11011 8520 11560 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 11532 8492 11560 8520
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12952 8520 13001 8548
rect 12952 8508 12958 8520
rect 12989 8517 13001 8520
rect 13035 8548 13047 8551
rect 13357 8551 13415 8557
rect 13357 8548 13369 8551
rect 13035 8520 13369 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 13357 8517 13369 8520
rect 13403 8517 13415 8551
rect 13357 8511 13415 8517
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 10008 8452 10057 8480
rect 10008 8440 10014 8452
rect 10045 8449 10057 8452
rect 10091 8480 10103 8483
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10091 8452 10609 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 11146 8480 11152 8492
rect 11107 8452 11152 8480
rect 10781 8443 10839 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11514 8440 11520 8492
rect 11572 8440 11578 8492
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12342 8480 12348 8492
rect 12303 8452 12348 8480
rect 12069 8443 12127 8449
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7374 8412 7380 8424
rect 7055 8384 7380 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 9766 8412 9772 8424
rect 9727 8384 9772 8412
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 10459 8384 10517 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 12084 8412 12112 8443
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 12894 8412 12900 8424
rect 12084 8384 12900 8412
rect 10505 8375 10563 8381
rect 12894 8372 12900 8384
rect 12952 8412 12958 8424
rect 13280 8412 13308 8443
rect 12952 8384 13308 8412
rect 12952 8372 12958 8384
rect 3326 8344 3332 8356
rect 3287 8316 3332 8344
rect 3326 8304 3332 8316
rect 3384 8304 3390 8356
rect 4798 8344 4804 8356
rect 4759 8316 4804 8344
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5718 8344 5724 8356
rect 5679 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6362 8344 6368 8356
rect 6323 8316 6368 8344
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 6914 8344 6920 8356
rect 6875 8316 6920 8344
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 10318 8344 10324 8356
rect 7892 8316 10324 8344
rect 7892 8304 7898 8316
rect 10318 8304 10324 8316
rect 10376 8344 10382 8356
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 10376 8316 11345 8344
rect 10376 8304 10382 8316
rect 11333 8313 11345 8316
rect 11379 8344 11391 8347
rect 11606 8344 11612 8356
rect 11379 8316 11612 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 11974 8344 11980 8356
rect 11935 8316 11980 8344
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 12124 8316 13461 8344
rect 12124 8304 12130 8316
rect 13449 8313 13461 8316
rect 13495 8313 13507 8347
rect 13449 8307 13507 8313
rect 6086 8276 6092 8288
rect 6047 8248 6092 8276
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 3878 8072 3884 8084
rect 3651 8044 3884 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 9306 8072 9312 8084
rect 8444 8044 9312 8072
rect 8444 8032 8450 8044
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11790 8072 11796 8084
rect 11379 8044 11796 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 4798 8004 4804 8016
rect 4571 7976 4804 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 7282 8004 7288 8016
rect 6288 7976 7288 8004
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3108 7908 3372 7936
rect 3108 7896 3114 7908
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2866 7868 2872 7880
rect 2823 7840 2872 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3344 7877 3372 7908
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3568 7908 4077 7936
rect 3568 7896 3574 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 6086 7936 6092 7948
rect 4663 7908 6092 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2924 7840 3157 7868
rect 2924 7828 2930 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5534 7868 5540 7880
rect 5491 7840 5540 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 2593 7803 2651 7809
rect 2593 7800 2605 7803
rect 2004 7772 2605 7800
rect 2004 7760 2010 7772
rect 2593 7769 2605 7772
rect 2639 7769 2651 7803
rect 2958 7800 2964 7812
rect 2919 7772 2964 7800
rect 2593 7763 2651 7769
rect 2958 7760 2964 7772
rect 3016 7760 3022 7812
rect 3053 7803 3111 7809
rect 3053 7769 3065 7803
rect 3099 7769 3111 7803
rect 4724 7800 4752 7831
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6181 7871 6239 7877
rect 5684 7840 5729 7868
rect 5684 7828 5690 7840
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6288 7868 6316 7976
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 13170 8004 13176 8016
rect 13131 7976 13176 8004
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 6822 7936 6828 7948
rect 6735 7908 6828 7936
rect 6822 7896 6828 7908
rect 6880 7936 6886 7948
rect 6880 7908 8524 7936
rect 6880 7896 6886 7908
rect 6227 7840 6316 7868
rect 6365 7871 6423 7877
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6411 7840 7205 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 4890 7800 4896 7812
rect 4724 7772 4896 7800
rect 3053 7763 3111 7769
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 3068 7732 3096 7763
rect 4890 7760 4896 7772
rect 4948 7800 4954 7812
rect 6454 7800 6460 7812
rect 4948 7772 6460 7800
rect 4948 7760 4954 7772
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 3878 7732 3884 7744
rect 2188 7704 3096 7732
rect 3839 7704 3884 7732
rect 2188 7692 2194 7704
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 7208 7732 7236 7831
rect 7392 7800 7420 7831
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 8496 7877 8524 7908
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9180 7908 9597 7936
rect 9180 7896 9186 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7524 7840 8309 7868
rect 7524 7828 7530 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 9381 7871 9439 7877
rect 9381 7837 9393 7871
rect 9427 7868 9439 7871
rect 9427 7837 9444 7868
rect 9381 7831 9444 7837
rect 8386 7800 8392 7812
rect 7392 7772 8392 7800
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 8628 7772 8953 7800
rect 8628 7760 8634 7772
rect 8941 7769 8953 7772
rect 8987 7769 8999 7803
rect 9122 7800 9128 7812
rect 9083 7772 9128 7800
rect 8941 7763 8999 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9416 7800 9444 7831
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9548 7840 9689 7868
rect 9548 7828 9554 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10100 7840 10149 7868
rect 10100 7828 10106 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11296 7840 11437 7868
rect 11296 7828 11302 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11839 7840 11897 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 11885 7837 11897 7840
rect 11931 7837 11943 7871
rect 12894 7868 12900 7880
rect 12855 7840 12900 7868
rect 11885 7831 11943 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 11609 7803 11667 7809
rect 9416 7772 10456 7800
rect 10428 7744 10456 7772
rect 11609 7769 11621 7803
rect 11655 7800 11667 7803
rect 12158 7800 12164 7812
rect 11655 7772 12164 7800
rect 11655 7769 11667 7772
rect 11609 7763 11667 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 7558 7732 7564 7744
rect 7208 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 8168 7704 8217 7732
rect 8168 7692 8174 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8662 7732 8668 7744
rect 8623 7704 8668 7732
rect 8205 7695 8263 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8812 7704 9505 7732
rect 8812 7692 8818 7704
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7528 2286 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 2280 7500 2421 7528
rect 2280 7488 2286 7500
rect 2409 7497 2421 7500
rect 2455 7497 2467 7531
rect 2409 7491 2467 7497
rect 2424 7460 2452 7491
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2924 7500 2973 7528
rect 2924 7488 2930 7500
rect 2961 7497 2973 7500
rect 3007 7528 3019 7531
rect 6546 7528 6552 7540
rect 3007 7500 6552 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8110 7528 8116 7540
rect 7975 7500 8116 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8110 7488 8116 7500
rect 8168 7528 8174 7540
rect 8846 7528 8852 7540
rect 8168 7500 8852 7528
rect 8168 7488 8174 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9398 7528 9404 7540
rect 9079 7500 9404 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9398 7488 9404 7500
rect 9456 7528 9462 7540
rect 9456 7500 9904 7528
rect 9456 7488 9462 7500
rect 2774 7460 2780 7472
rect 2424 7432 2780 7460
rect 2774 7420 2780 7432
rect 2832 7460 2838 7472
rect 4798 7460 4804 7472
rect 2832 7432 3740 7460
rect 2832 7420 2838 7432
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 3712 7401 3740 7432
rect 4540 7432 4804 7460
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3878 7392 3884 7404
rect 3743 7364 3884 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3050 7324 3056 7336
rect 3011 7296 3056 7324
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3237 7287 3295 7293
rect 3252 7256 3280 7287
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3620 7324 3648 7355
rect 3878 7352 3884 7364
rect 3936 7392 3942 7404
rect 4540 7401 4568 7432
rect 4798 7420 4804 7432
rect 4856 7420 4862 7472
rect 5353 7463 5411 7469
rect 5353 7429 5365 7463
rect 5399 7460 5411 7463
rect 5534 7460 5540 7472
rect 5399 7432 5540 7460
rect 5399 7429 5411 7432
rect 5353 7423 5411 7429
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 8662 7460 8668 7472
rect 5684 7432 6224 7460
rect 5684 7420 5690 7432
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3936 7364 3985 7392
rect 3936 7352 3942 7364
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4709 7355 4767 7361
rect 4172 7324 4200 7355
rect 3620 7296 4200 7324
rect 3712 7268 3740 7296
rect 3510 7256 3516 7268
rect 3252 7228 3516 7256
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 3694 7216 3700 7268
rect 3752 7216 3758 7268
rect 4172 7256 4200 7296
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4614 7324 4620 7336
rect 4387 7296 4620 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4724 7324 4752 7355
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6196 7401 6224 7432
rect 6840 7432 8668 7460
rect 6840 7401 6868 7432
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 9048 7432 9352 7460
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7374 7392 7380 7404
rect 6972 7364 7017 7392
rect 7335 7364 7380 7392
rect 6972 7352 6978 7364
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 7558 7392 7564 7404
rect 7519 7364 7564 7392
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 7834 7401 7840 7404
rect 7817 7395 7840 7401
rect 7817 7361 7829 7395
rect 7817 7355 7840 7361
rect 7834 7352 7840 7355
rect 7892 7352 7898 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8202 7392 8208 7404
rect 8067 7364 8208 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8478 7392 8484 7404
rect 8439 7364 8484 7392
rect 8478 7352 8484 7364
rect 8536 7392 8542 7404
rect 9048 7392 9076 7432
rect 9214 7401 9220 7404
rect 8536 7364 9076 7392
rect 9183 7395 9220 7401
rect 8536 7352 8542 7364
rect 9183 7361 9195 7395
rect 9183 7355 9220 7361
rect 9214 7352 9220 7355
rect 9272 7352 9278 7404
rect 4982 7324 4988 7336
rect 4724 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7293 5503 7327
rect 7098 7324 7104 7336
rect 7059 7296 7104 7324
rect 5445 7287 5503 7293
rect 5460 7256 5488 7287
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7282 7324 7288 7336
rect 7239 7296 7288 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7282 7284 7288 7296
rect 7340 7324 7346 7336
rect 7926 7324 7932 7336
rect 7340 7296 7932 7324
rect 7340 7284 7346 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8294 7324 8300 7336
rect 8159 7296 8300 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8294 7284 8300 7296
rect 8352 7324 8358 7336
rect 8570 7324 8576 7336
rect 8352 7296 8576 7324
rect 8352 7284 8358 7296
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 8754 7324 8760 7336
rect 8711 7296 8760 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 8754 7284 8760 7296
rect 8812 7324 8818 7336
rect 9030 7324 9036 7336
rect 8812 7296 9036 7324
rect 8812 7284 8818 7296
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9324 7324 9352 7432
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 9876 7460 9904 7500
rect 10318 7460 10324 7472
rect 9548 7432 9628 7460
rect 9876 7432 9996 7460
rect 10279 7432 10324 7460
rect 9548 7420 9554 7432
rect 9600 7401 9628 7432
rect 9590 7395 9648 7401
rect 9590 7361 9602 7395
rect 9636 7361 9648 7395
rect 9590 7355 9648 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 9677 7355 9735 7361
rect 9473 7327 9531 7333
rect 9473 7324 9485 7327
rect 9324 7296 9485 7324
rect 9473 7293 9485 7296
rect 9519 7293 9531 7327
rect 9692 7324 9720 7355
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 9968 7401 9996 7432
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12345 7463 12403 7469
rect 12345 7460 12357 7463
rect 12124 7432 12357 7460
rect 12124 7420 12130 7432
rect 12345 7429 12357 7432
rect 12391 7429 12403 7463
rect 12345 7423 12403 7429
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10046 7395 10104 7401
rect 10046 7361 10058 7395
rect 10092 7392 10104 7395
rect 10134 7392 10140 7404
rect 10092 7364 10140 7392
rect 10092 7361 10104 7364
rect 10046 7355 10104 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 9692 7296 9904 7324
rect 9473 7287 9531 7293
rect 9876 7268 9904 7296
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11296 7296 11805 7324
rect 11296 7284 11302 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12124 7296 12449 7324
rect 12124 7284 12130 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12851 7296 12909 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 5997 7259 6055 7265
rect 5997 7256 6009 7259
rect 4172 7228 5396 7256
rect 5460 7228 6009 7256
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 1946 7188 1952 7200
rect 1811 7160 1952 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2590 7188 2596 7200
rect 2551 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4798 7188 4804 7200
rect 4755 7160 4804 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5368 7188 5396 7228
rect 5997 7225 6009 7228
rect 6043 7225 6055 7259
rect 5997 7219 6055 7225
rect 9858 7216 9864 7268
rect 9916 7216 9922 7268
rect 12250 7256 12256 7268
rect 12211 7228 12256 7256
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 6454 7188 6460 7200
rect 5368 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6638 7188 6644 7200
rect 6599 7160 6644 7188
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8570 7188 8576 7200
rect 8343 7160 8576 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 12268 7188 12296 7216
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12268 7160 12817 7188
rect 12805 7157 12817 7160
rect 12851 7188 12863 7191
rect 13170 7188 13176 7200
rect 12851 7160 13176 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 2028 6987 2086 6993
rect 2028 6953 2040 6987
rect 2074 6984 2086 6987
rect 2590 6984 2596 6996
rect 2074 6956 2596 6984
rect 2074 6953 2086 6956
rect 2028 6947 2086 6953
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3513 6987 3571 6993
rect 3513 6984 3525 6987
rect 3108 6956 3525 6984
rect 3108 6944 3114 6956
rect 3513 6953 3525 6956
rect 3559 6953 3571 6987
rect 3513 6947 3571 6953
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 5902 6984 5908 6996
rect 4120 6956 5908 6984
rect 4120 6944 4126 6956
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 6076 6987 6134 6993
rect 6076 6953 6088 6987
rect 6122 6984 6134 6987
rect 6638 6984 6644 6996
rect 6122 6956 6644 6984
rect 6122 6953 6134 6956
rect 6076 6947 6134 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9950 6984 9956 6996
rect 8536 6956 9956 6984
rect 8536 6944 8542 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 9398 6916 9404 6928
rect 7156 6888 9404 6916
rect 7156 6876 7162 6888
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 1811 6820 3801 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 3789 6817 3801 6820
rect 3835 6848 3847 6851
rect 5258 6848 5264 6860
rect 3835 6820 5264 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 5258 6808 5264 6820
rect 5316 6848 5322 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5316 6820 5825 6848
rect 5316 6808 5322 6820
rect 5813 6817 5825 6820
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 7926 6848 7932 6860
rect 7607 6820 7932 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8294 6848 8300 6860
rect 8067 6820 8300 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8294 6808 8300 6820
rect 8352 6848 8358 6860
rect 8662 6848 8668 6860
rect 8352 6820 8668 6848
rect 8352 6808 8358 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9232 6857 9260 6888
rect 9398 6876 9404 6888
rect 9456 6916 9462 6928
rect 9858 6916 9864 6928
rect 9456 6888 9864 6916
rect 9456 6876 9462 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 13265 6919 13323 6925
rect 13265 6916 13277 6919
rect 12952 6888 13277 6916
rect 12952 6876 12958 6888
rect 13265 6885 13277 6888
rect 13311 6885 13323 6919
rect 13265 6879 13323 6885
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6817 9275 6851
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 9217 6811 9275 6817
rect 9416 6820 11621 6848
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9416 6789 9444 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11882 6808 11888 6860
rect 11940 6808 11946 6860
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 8812 6752 9413 6780
rect 8812 6740 8818 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9732 6752 9873 6780
rect 9732 6740 9738 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 11900 6780 11928 6808
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11900 6752 11989 6780
rect 9861 6743 9919 6749
rect 11977 6749 11989 6752
rect 12023 6780 12035 6783
rect 12342 6780 12348 6792
rect 12023 6752 12348 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 3418 6712 3424 6724
rect 3266 6684 3424 6712
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 4062 6712 4068 6724
rect 4023 6684 4068 6712
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 4614 6672 4620 6724
rect 4672 6672 4678 6724
rect 6638 6672 6644 6724
rect 6696 6672 6702 6724
rect 7374 6672 7380 6724
rect 7432 6712 7438 6724
rect 8772 6712 8800 6740
rect 7432 6684 8800 6712
rect 10137 6715 10195 6721
rect 7432 6672 7438 6684
rect 10137 6681 10149 6715
rect 10183 6681 10195 6715
rect 11882 6712 11888 6724
rect 11362 6684 11888 6712
rect 10137 6675 10195 6681
rect 1394 6644 1400 6656
rect 1355 6616 1400 6644
rect 1394 6604 1400 6616
rect 1452 6604 1458 6656
rect 1673 6647 1731 6653
rect 1673 6613 1685 6647
rect 1719 6644 1731 6647
rect 1762 6644 1768 6656
rect 1719 6616 1768 6644
rect 1719 6613 1731 6616
rect 1673 6607 1731 6613
rect 1762 6604 1768 6616
rect 1820 6604 1826 6656
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4430 6644 4436 6656
rect 3568 6616 4436 6644
rect 3568 6604 3574 6616
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 5534 6644 5540 6656
rect 5495 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 8754 6644 8760 6656
rect 8527 6616 8760 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 9088 6616 9321 6644
rect 9088 6604 9094 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10152 6644 10180 6675
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 9815 6616 10180 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 4062 6440 4068 6452
rect 2004 6412 3096 6440
rect 4023 6412 4068 6440
rect 2004 6400 2010 6412
rect 1964 6344 2360 6372
rect 1394 6264 1400 6316
rect 1452 6304 1458 6316
rect 1964 6313 1992 6344
rect 2332 6316 2360 6344
rect 1823 6307 1881 6313
rect 1823 6304 1835 6307
rect 1452 6276 1835 6304
rect 1452 6264 1458 6276
rect 1823 6273 1835 6276
rect 1869 6273 1881 6307
rect 1823 6267 1881 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2056 6236 2084 6267
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2188 6276 2237 6304
rect 2188 6264 2194 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 3068 6313 3096 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 4706 6440 4712 6452
rect 4571 6412 4712 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 4706 6400 4712 6412
rect 4764 6440 4770 6452
rect 5534 6440 5540 6452
rect 4764 6412 5540 6440
rect 4764 6400 4770 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6409 7343 6443
rect 8570 6440 8576 6452
rect 7285 6403 7343 6409
rect 7760 6412 8576 6440
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4614 6372 4620 6384
rect 4019 6344 4620 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 5169 6375 5227 6381
rect 5169 6341 5181 6375
rect 5215 6372 5227 6375
rect 5258 6372 5264 6384
rect 5215 6344 5264 6372
rect 5215 6341 5227 6344
rect 5169 6335 5227 6341
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 7300 6372 7328 6403
rect 6512 6344 6776 6372
rect 7300 6344 7512 6372
rect 6512 6332 6518 6344
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2372 6276 2417 6304
rect 2516 6276 2973 6304
rect 2372 6264 2378 6276
rect 2516 6236 2544 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 3053 6267 3111 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3384 6276 3801 6304
rect 3384 6264 3390 6276
rect 3789 6273 3801 6276
rect 3835 6304 3847 6307
rect 4062 6304 4068 6316
rect 3835 6276 4068 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 4433 6267 4491 6273
rect 2056 6208 2544 6236
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 1578 6168 1584 6180
rect 1539 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 2409 6171 2467 6177
rect 2409 6168 2421 6171
rect 1728 6140 2421 6168
rect 1728 6128 1734 6140
rect 2409 6137 2421 6140
rect 2455 6137 2467 6171
rect 2409 6131 2467 6137
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6100 1458 6112
rect 2608 6100 2636 6199
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4448 6236 4476 6267
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 6748 6313 6776 6344
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6420 6276 6561 6304
rect 6420 6264 6426 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 7098 6304 7104 6316
rect 7059 6276 7104 6304
rect 6733 6267 6791 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7484 6313 7512 6344
rect 7760 6313 7788 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 8904 6412 9812 6440
rect 8904 6400 8910 6412
rect 9030 6372 9036 6384
rect 8991 6344 9036 6372
rect 9030 6332 9036 6344
rect 9088 6332 9094 6384
rect 8668 6316 8720 6322
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8018 6304 8024 6316
rect 7883 6276 8024 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9784 6313 9812 6412
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11330 6440 11336 6452
rect 10008 6412 10640 6440
rect 11291 6412 11336 6440
rect 10008 6400 10014 6412
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 8812 6276 9505 6304
rect 8812 6264 8818 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10612 6313 10640 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11808 6412 12204 6440
rect 11348 6372 11376 6400
rect 11808 6372 11836 6412
rect 11348 6344 11836 6372
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10100 6276 10425 6304
rect 10100 6264 10106 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 11808 6313 11836 6344
rect 11882 6332 11888 6384
rect 11940 6372 11946 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11940 6344 11989 6372
rect 11940 6332 11946 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 12176 6372 12204 6412
rect 12437 6375 12495 6381
rect 12437 6372 12449 6375
rect 12176 6344 12449 6372
rect 11977 6335 12035 6341
rect 11701 6307 11759 6313
rect 10744 6276 10789 6304
rect 10744 6264 10750 6276
rect 11701 6273 11713 6307
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 3568 6208 4476 6236
rect 3568 6196 3574 6208
rect 3602 6168 3608 6180
rect 3563 6140 3608 6168
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 4448 6168 4476 6208
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4580 6208 4721 6236
rect 4580 6196 4586 6208
rect 4709 6205 4721 6208
rect 4755 6236 4767 6239
rect 5350 6236 5356 6248
rect 4755 6208 5356 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7116 6236 7144 6264
rect 8668 6258 8720 6264
rect 7558 6236 7564 6248
rect 7116 6208 7564 6236
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8772 6208 9137 6236
rect 5166 6168 5172 6180
rect 4448 6140 5172 6168
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 5960 6140 8432 6168
rect 5960 6128 5966 6140
rect 1452 6072 2636 6100
rect 2777 6103 2835 6109
rect 1452 6060 1458 6072
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2958 6100 2964 6112
rect 2823 6072 2964 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 6362 6100 6368 6112
rect 5684 6072 6368 6100
rect 5684 6060 5690 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 8404 6100 8432 6140
rect 8478 6128 8484 6180
rect 8536 6168 8542 6180
rect 8772 6168 8800 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 10318 6236 10324 6248
rect 9364 6208 10324 6236
rect 9364 6196 9370 6208
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10778 6236 10784 6248
rect 10612 6208 10784 6236
rect 8536 6140 8800 6168
rect 10505 6171 10563 6177
rect 8536 6128 8542 6140
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 10612 6168 10640 6208
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 11716 6236 11744 6267
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12268 6313 12296 6344
rect 12437 6341 12449 6344
rect 12483 6341 12495 6375
rect 12437 6335 12495 6341
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 13081 6375 13139 6381
rect 13081 6372 13093 6375
rect 13044 6344 13093 6372
rect 13044 6332 13050 6344
rect 13081 6341 13093 6344
rect 13127 6341 13139 6375
rect 13081 6335 13139 6341
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 12124 6276 12173 6304
rect 12124 6264 12130 6276
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12621 6307 12679 6313
rect 12621 6304 12633 6307
rect 12400 6276 12633 6304
rect 12400 6264 12406 6276
rect 12621 6273 12633 6276
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 13173 6239 13231 6245
rect 11716 6208 11836 6236
rect 11606 6168 11612 6180
rect 10551 6140 10640 6168
rect 11567 6140 11612 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 11808 6168 11836 6208
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 13262 6236 13268 6248
rect 13219 6208 13268 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 12066 6168 12072 6180
rect 11808 6140 12072 6168
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 9030 6100 9036 6112
rect 8404 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10376 6072 10885 6100
rect 10376 6060 10382 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 4706 5896 4712 5908
rect 3528 5868 4712 5896
rect 2225 5831 2283 5837
rect 2225 5797 2237 5831
rect 2271 5828 2283 5831
rect 2314 5828 2320 5840
rect 2271 5800 2320 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 3326 5828 3332 5840
rect 3287 5800 3332 5828
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 3528 5760 3556 5868
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5258 5896 5264 5908
rect 4816 5868 5264 5896
rect 1872 5732 2774 5760
rect 1872 5701 1900 5732
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2332 5701 2360 5732
rect 2317 5695 2375 5701
rect 2004 5664 2049 5692
rect 2004 5652 2010 5664
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2590 5692 2596 5704
rect 2551 5664 2596 5692
rect 2409 5655 2467 5661
rect 1964 5624 1992 5652
rect 2424 5624 2452 5655
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 1964 5596 2452 5624
rect 2746 5624 2774 5732
rect 3436 5732 3556 5760
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3050 5692 3056 5704
rect 3007 5664 3056 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3436 5701 3464 5732
rect 3786 5720 3792 5772
rect 3844 5760 3850 5772
rect 4816 5769 4844 5868
rect 5258 5856 5264 5868
rect 5316 5896 5322 5908
rect 6546 5896 6552 5908
rect 5316 5868 6408 5896
rect 6507 5868 6552 5896
rect 5316 5856 5322 5868
rect 6380 5828 6408 5868
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 9214 5896 9220 5908
rect 9175 5868 9220 5896
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 10594 5896 10600 5908
rect 9539 5868 10600 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11756 5868 12081 5896
rect 11756 5856 11762 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 12069 5859 12127 5865
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 6914 5828 6920 5840
rect 6380 5800 6920 5828
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 9398 5828 9404 5840
rect 8220 5800 9404 5828
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 3844 5732 4813 5760
rect 3844 5720 3850 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8220 5769 8248 5800
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 9674 5788 9680 5840
rect 9732 5788 9738 5840
rect 10042 5828 10048 5840
rect 10003 5800 10048 5828
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7984 5732 8217 5760
rect 7984 5720 7990 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8478 5760 8484 5772
rect 8343 5732 8484 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 9692 5760 9720 5788
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 9692 5732 10333 5760
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10962 5760 10968 5772
rect 10643 5732 10968 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 3421 5695 3479 5701
rect 3200 5664 3245 5692
rect 3200 5652 3206 5664
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3568 5664 3613 5692
rect 3568 5652 3574 5664
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 4120 5664 4445 5692
rect 4120 5652 4126 5664
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6696 5664 7021 5692
rect 6696 5652 6702 5664
rect 7009 5661 7021 5664
rect 7055 5692 7067 5695
rect 7098 5692 7104 5704
rect 7055 5664 7104 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 8846 5692 8852 5704
rect 7515 5664 8852 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9306 5692 9312 5704
rect 9267 5664 9312 5692
rect 9033 5655 9091 5661
rect 3234 5624 3240 5636
rect 2746 5596 3240 5624
rect 3234 5584 3240 5596
rect 3292 5624 3298 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3292 5596 3801 5624
rect 3292 5584 3298 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3970 5624 3976 5636
rect 3931 5596 3976 5624
rect 3789 5587 3847 5593
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4614 5624 4620 5636
rect 4387 5596 4620 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5074 5624 5080 5636
rect 5035 5596 5080 5624
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 5718 5584 5724 5636
rect 5776 5584 5782 5636
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 8570 5624 8576 5636
rect 8435 5596 8576 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 8570 5584 8576 5596
rect 8628 5584 8634 5636
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9048 5624 9076 5655
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 9675 5695 9733 5701
rect 9675 5692 9687 5695
rect 9456 5664 9687 5692
rect 9456 5652 9462 5664
rect 9675 5661 9687 5664
rect 9721 5692 9733 5695
rect 10137 5695 10195 5701
rect 9721 5664 9996 5692
rect 9721 5661 9733 5664
rect 9675 5655 9733 5661
rect 9858 5624 9864 5636
rect 8720 5596 9076 5624
rect 9416 5596 9864 5624
rect 8720 5584 8726 5596
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 1762 5556 1768 5568
rect 1535 5528 1768 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2685 5559 2743 5565
rect 2685 5556 2697 5559
rect 1912 5528 2697 5556
rect 1912 5516 1918 5528
rect 2685 5525 2697 5528
rect 2731 5525 2743 5559
rect 4062 5556 4068 5568
rect 4023 5528 4068 5556
rect 2685 5519 2743 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 4203 5528 4537 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 4525 5525 4537 5528
rect 4571 5525 4583 5559
rect 4525 5519 4583 5525
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 7837 5559 7895 5565
rect 7837 5556 7849 5559
rect 7800 5528 7849 5556
rect 7800 5516 7806 5528
rect 7837 5525 7849 5528
rect 7883 5525 7895 5559
rect 7837 5519 7895 5525
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 9416 5556 9444 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 9968 5624 9996 5664
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10226 5692 10232 5704
rect 10183 5664 10232 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10318 5624 10324 5636
rect 9968 5596 10324 5624
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 11606 5584 11612 5636
rect 11664 5584 11670 5636
rect 8803 5528 9444 5556
rect 9677 5559 9735 5565
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 9766 5556 9772 5568
rect 9723 5528 9772 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 2590 5352 2596 5364
rect 1820 5324 2596 5352
rect 1820 5312 1826 5324
rect 2590 5312 2596 5324
rect 2648 5352 2654 5364
rect 2685 5355 2743 5361
rect 2685 5352 2697 5355
rect 2648 5324 2697 5352
rect 2648 5312 2654 5324
rect 2685 5321 2697 5324
rect 2731 5321 2743 5355
rect 2685 5315 2743 5321
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 3660 5324 4476 5352
rect 3660 5312 3666 5324
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 2777 5287 2835 5293
rect 2777 5284 2789 5287
rect 1995 5256 2789 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 2777 5253 2789 5256
rect 2823 5284 2835 5287
rect 3050 5284 3056 5296
rect 2823 5256 3056 5284
rect 2823 5253 2835 5256
rect 2777 5247 2835 5253
rect 3050 5244 3056 5256
rect 3108 5284 3114 5296
rect 3973 5287 4031 5293
rect 3973 5284 3985 5287
rect 3108 5256 3985 5284
rect 3108 5244 3114 5256
rect 3973 5253 3985 5256
rect 4019 5253 4031 5287
rect 4249 5287 4307 5293
rect 4249 5284 4261 5287
rect 3973 5247 4031 5253
rect 4080 5256 4261 5284
rect 4080 5228 4108 5256
rect 4249 5253 4261 5256
rect 4295 5253 4307 5287
rect 4249 5247 4307 5253
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2406 5216 2412 5228
rect 2363 5188 2412 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2056 5148 2084 5179
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2792 5188 2973 5216
rect 2792 5160 2820 5188
rect 2961 5185 2973 5188
rect 3007 5216 3019 5219
rect 3237 5219 3295 5225
rect 3007 5188 3096 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3068 5160 3096 5188
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3237 5179 3295 5185
rect 2590 5157 2596 5160
rect 2576 5151 2596 5157
rect 2056 5120 2452 5148
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 2314 5080 2320 5092
rect 1627 5052 2320 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 2314 5040 2320 5052
rect 2372 5040 2378 5092
rect 2424 5080 2452 5120
rect 2576 5117 2588 5151
rect 2576 5111 2596 5117
rect 2590 5108 2596 5111
rect 2648 5108 2654 5160
rect 2774 5108 2780 5160
rect 2832 5108 2838 5160
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5117 2927 5151
rect 2869 5111 2927 5117
rect 2884 5080 2912 5111
rect 3050 5108 3056 5160
rect 3108 5108 3114 5160
rect 3252 5148 3280 5179
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 3881 5179 3939 5185
rect 3694 5148 3700 5160
rect 3252 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 3896 5148 3924 5179
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4448 5225 4476 5324
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 4893 5355 4951 5361
rect 4893 5352 4905 5355
rect 4672 5324 4905 5352
rect 4672 5312 4678 5324
rect 4893 5321 4905 5324
rect 4939 5321 4951 5355
rect 4893 5315 4951 5321
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5132 5324 5457 5352
rect 5132 5312 5138 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 6546 5312 6552 5364
rect 6604 5312 6610 5364
rect 9490 5352 9496 5364
rect 9048 5324 9496 5352
rect 5534 5284 5540 5296
rect 5092 5256 5540 5284
rect 5092 5225 5120 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 6564 5284 6592 5312
rect 8570 5284 8576 5296
rect 5920 5256 6592 5284
rect 8418 5256 8576 5284
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 3970 5148 3976 5160
rect 3896 5120 3976 5148
rect 3970 5108 3976 5120
rect 4028 5148 4034 5160
rect 4172 5148 4200 5179
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5920 5225 5948 5256
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 8846 5284 8852 5296
rect 8807 5256 8852 5284
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 5905 5219 5963 5225
rect 5224 5188 5764 5216
rect 5224 5176 5230 5188
rect 4028 5120 4200 5148
rect 4028 5108 4034 5120
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 5408 5120 5641 5148
rect 5408 5108 5414 5120
rect 5629 5117 5641 5120
rect 5675 5117 5687 5151
rect 5736 5148 5764 5188
rect 5905 5185 5917 5219
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6144 5188 6561 5216
rect 6144 5176 6150 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6914 5216 6920 5228
rect 6875 5188 6920 5216
rect 6549 5179 6607 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 9048 5225 9076 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 12262 5355 12320 5361
rect 12262 5352 12274 5355
rect 11480 5324 12274 5352
rect 11480 5312 11486 5324
rect 12262 5321 12274 5324
rect 12308 5321 12320 5355
rect 12262 5315 12320 5321
rect 9674 5284 9680 5296
rect 9508 5256 9680 5284
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8536 5188 9045 5216
rect 8536 5176 8542 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9508 5225 9536 5256
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 9769 5287 9827 5293
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 9858 5284 9864 5296
rect 9815 5256 9864 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11517 5287 11575 5293
rect 11517 5284 11529 5287
rect 11388 5256 11529 5284
rect 11388 5244 11394 5256
rect 11517 5253 11529 5256
rect 11563 5284 11575 5287
rect 11701 5287 11759 5293
rect 11701 5284 11713 5287
rect 11563 5256 11713 5284
rect 11563 5253 11575 5256
rect 11517 5247 11575 5253
rect 11701 5253 11713 5256
rect 11747 5284 11759 5287
rect 11882 5284 11888 5296
rect 11747 5256 11888 5284
rect 11747 5253 11759 5256
rect 11701 5247 11759 5253
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 13170 5244 13176 5296
rect 13228 5284 13234 5296
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 13228 5256 13277 5284
rect 13228 5244 13234 5256
rect 13265 5253 13277 5256
rect 13311 5253 13323 5287
rect 13265 5247 13323 5253
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5185 9551 5219
rect 11606 5216 11612 5228
rect 10902 5188 11612 5216
rect 9493 5179 9551 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 12618 5216 12624 5228
rect 12579 5188 12624 5216
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5736 5120 6377 5148
rect 5629 5111 5687 5117
rect 6365 5117 6377 5120
rect 6411 5148 6423 5151
rect 6454 5148 6460 5160
rect 6411 5120 6460 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 2424 5052 2912 5080
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2884 5012 2912 5052
rect 3237 5083 3295 5089
rect 3237 5049 3249 5083
rect 3283 5080 3295 5083
rect 4706 5080 4712 5092
rect 3283 5052 4712 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5644 5080 5672 5111
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7282 5148 7288 5160
rect 7239 5120 7288 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 9122 5148 9128 5160
rect 8812 5120 9128 5148
rect 8812 5108 8818 5120
rect 9122 5108 9128 5120
rect 9180 5148 9186 5160
rect 11146 5148 11152 5160
rect 9180 5120 11152 5148
rect 9180 5108 9186 5120
rect 11146 5108 11152 5120
rect 11204 5148 11210 5160
rect 11204 5120 11284 5148
rect 11204 5108 11210 5120
rect 5813 5083 5871 5089
rect 5644 5052 5764 5080
rect 3142 5012 3148 5024
rect 2884 4984 3148 5012
rect 3142 4972 3148 4984
rect 3200 5012 3206 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 3200 4984 4629 5012
rect 3200 4972 3206 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 5736 5012 5764 5052
rect 5813 5049 5825 5083
rect 5859 5080 5871 5083
rect 6733 5083 6791 5089
rect 6733 5080 6745 5083
rect 5859 5052 6745 5080
rect 5859 5049 5871 5052
rect 5813 5043 5871 5049
rect 6733 5049 6745 5052
rect 6779 5080 6791 5083
rect 6822 5080 6828 5092
rect 6779 5052 6828 5080
rect 6779 5049 6791 5052
rect 6733 5043 6791 5049
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 11256 5089 11284 5120
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 11287 5052 12296 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 5902 5012 5908 5024
rect 5736 4984 5908 5012
rect 4617 4975 4675 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 8662 5012 8668 5024
rect 8623 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 12268 5021 12296 5052
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12710 5012 12716 5024
rect 12483 4984 12716 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 3878 4808 3884 4820
rect 2746 4780 3884 4808
rect 2590 4740 2596 4752
rect 1412 4712 2596 4740
rect 1412 4480 1440 4712
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 1854 4672 1860 4684
rect 1815 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2746 4672 2774 4780
rect 3878 4768 3884 4780
rect 3936 4808 3942 4820
rect 4798 4808 4804 4820
rect 3936 4780 4804 4808
rect 3936 4768 3942 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8478 4808 8484 4820
rect 8439 4780 8484 4808
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 8812 4780 9229 4808
rect 8812 4768 8818 4780
rect 9217 4777 9229 4780
rect 9263 4808 9275 4811
rect 9306 4808 9312 4820
rect 9263 4780 9312 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9306 4768 9312 4780
rect 9364 4808 9370 4820
rect 10134 4808 10140 4820
rect 9364 4780 10140 4808
rect 9364 4768 9370 4780
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 10284 4780 12081 4808
rect 10284 4768 10290 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12069 4771 12127 4777
rect 2958 4749 2964 4752
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4709 2927 4743
rect 2869 4703 2927 4709
rect 2957 4703 2964 4749
rect 3016 4740 3022 4752
rect 3237 4743 3295 4749
rect 3016 4712 3057 4740
rect 2700 4644 2774 4672
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1728 4576 1777 4604
rect 1728 4564 1734 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2130 4604 2136 4616
rect 2087 4576 2136 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 2280 4576 2421 4604
rect 2280 4564 2286 4576
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2700 4604 2728 4644
rect 2639 4576 2728 4604
rect 2777 4607 2835 4613
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 1578 4496 1584 4548
rect 1636 4536 1642 4548
rect 2792 4536 2820 4567
rect 2884 4548 2912 4703
rect 2958 4700 2964 4703
rect 3016 4700 3022 4712
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 6638 4740 6644 4752
rect 3283 4712 3924 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 3786 4672 3792 4684
rect 3747 4644 3792 4672
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 3896 4672 3924 4712
rect 5828 4712 6644 4740
rect 5828 4672 5856 4712
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 6733 4743 6791 4749
rect 6733 4709 6745 4743
rect 6779 4709 6791 4743
rect 6733 4703 6791 4709
rect 6748 4672 6776 4703
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7064 4712 9628 4740
rect 7064 4700 7070 4712
rect 3896 4644 5856 4672
rect 5920 4644 6776 4672
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 5810 4604 5816 4616
rect 5767 4576 5816 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 1636 4508 2820 4536
rect 1636 4496 1642 4508
rect 2866 4496 2872 4548
rect 2924 4496 2930 4548
rect 1394 4468 1400 4480
rect 1355 4440 1400 4468
rect 1394 4428 1400 4440
rect 1452 4428 1458 4480
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 3068 4468 3096 4567
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5920 4613 5948 4644
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7742 4672 7748 4684
rect 6880 4644 6925 4672
rect 7703 4644 7748 4672
rect 6880 4632 6886 4644
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 7926 4672 7932 4684
rect 7887 4644 7932 4672
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 6123 4607 6181 4613
rect 5905 4567 5963 4573
rect 5998 4585 6056 4591
rect 5998 4551 6010 4585
rect 6044 4551 6056 4585
rect 6123 4573 6135 4607
rect 6169 4604 6181 4607
rect 6454 4604 6460 4616
rect 6169 4576 6460 4604
rect 6169 4573 6181 4576
rect 6123 4567 6181 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7653 4607 7711 4613
rect 6604 4576 6649 4604
rect 6604 4564 6610 4576
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 7699 4576 8585 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8573 4573 8585 4576
rect 8619 4604 8631 4607
rect 8662 4604 8668 4616
rect 8619 4576 8668 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 8662 4564 8668 4576
rect 8720 4604 8726 4616
rect 9600 4613 9628 4712
rect 9674 4700 9680 4752
rect 9732 4700 9738 4752
rect 13170 4740 13176 4752
rect 13131 4712 13176 4740
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 9692 4672 9720 4700
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9692 4644 10333 4672
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10321 4635 10379 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 11940 4644 12572 4672
rect 11940 4632 11946 4644
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 8720 4576 9229 4604
rect 8720 4564 8726 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9950 4604 9956 4616
rect 9723 4576 9956 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 10045 4567 10103 4573
rect 5998 4548 6056 4551
rect 4065 4539 4123 4545
rect 4065 4505 4077 4539
rect 4111 4536 4123 4539
rect 4338 4536 4344 4548
rect 4111 4508 4344 4536
rect 4111 4505 4123 4508
rect 4065 4499 4123 4505
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4706 4496 4712 4548
rect 4764 4496 4770 4548
rect 5626 4536 5632 4548
rect 5368 4508 5632 4536
rect 2639 4440 3096 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3513 4471 3571 4477
rect 3513 4468 3525 4471
rect 3200 4440 3525 4468
rect 3200 4428 3206 4440
rect 3513 4437 3525 4440
rect 3559 4468 3571 4471
rect 3602 4468 3608 4480
rect 3559 4440 3608 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3602 4428 3608 4440
rect 3660 4468 3666 4480
rect 5368 4468 5396 4508
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 5994 4496 6000 4548
rect 6052 4496 6058 4548
rect 6365 4539 6423 4545
rect 6365 4505 6377 4539
rect 6411 4536 6423 4539
rect 7926 4536 7932 4548
rect 6411 4508 7932 4536
rect 6411 4505 6423 4508
rect 6365 4499 6423 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8754 4536 8760 4548
rect 8715 4508 8760 4536
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 9858 4536 9864 4548
rect 9819 4508 9864 4536
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 10060 4536 10088 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12544 4613 12572 4644
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 12124 4576 12357 4604
rect 12124 4564 12130 4576
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12676 4576 12725 4604
rect 12676 4564 12682 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 12713 4567 12771 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 10134 4536 10140 4548
rect 10060 4508 10140 4536
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 11822 4508 12265 4536
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 12253 4499 12311 4505
rect 13265 4539 13323 4545
rect 13265 4505 13277 4539
rect 13311 4505 13323 4539
rect 13265 4499 13323 4505
rect 5534 4468 5540 4480
rect 3660 4440 5396 4468
rect 5495 4440 5540 4468
rect 3660 4428 3666 4440
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5644 4468 5672 4496
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 5644 4440 8125 4468
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9214 4468 9220 4480
rect 9079 4440 9220 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 13280 4468 13308 4499
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13280 4440 13369 4468
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 1489 4267 1547 4273
rect 1489 4233 1501 4267
rect 1535 4264 1547 4267
rect 1762 4264 1768 4276
rect 1535 4236 1768 4264
rect 1535 4233 1547 4236
rect 1489 4227 1547 4233
rect 1762 4224 1768 4236
rect 1820 4224 1826 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4525 4267 4583 4273
rect 4525 4264 4537 4267
rect 4396 4236 4537 4264
rect 4396 4224 4402 4236
rect 4525 4233 4537 4236
rect 4571 4233 4583 4267
rect 4525 4227 4583 4233
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5534 4264 5540 4276
rect 5031 4236 5540 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 4062 4196 4068 4208
rect 4023 4168 4068 4196
rect 4062 4156 4068 4168
rect 4120 4156 4126 4208
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 5000 4196 5028 4227
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5718 4264 5724 4276
rect 5679 4236 5724 4264
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6454 4264 6460 4276
rect 6415 4236 6460 4264
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 8570 4264 8576 4276
rect 6972 4236 8156 4264
rect 8531 4236 8576 4264
rect 6972 4224 6978 4236
rect 4479 4168 5028 4196
rect 8128 4196 8156 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 11606 4264 11612 4276
rect 11567 4236 11612 4264
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 12802 4264 12808 4276
rect 11940 4236 12808 4264
rect 11940 4224 11946 4236
rect 9674 4196 9680 4208
rect 8128 4168 8248 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 1670 4128 1676 4140
rect 1627 4100 1676 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2130 4128 2136 4140
rect 1811 4100 2136 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2866 4128 2872 4140
rect 2547 4100 2872 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3292 4100 3433 4128
rect 3292 4088 3298 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4295 4100 4905 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4893 4097 4905 4100
rect 4939 4128 4951 4131
rect 5258 4128 5264 4140
rect 4939 4100 5264 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5626 4128 5632 4140
rect 5583 4100 5632 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6362 4128 6368 4140
rect 5951 4100 6368 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6362 4088 6368 4100
rect 6420 4128 6426 4140
rect 6638 4128 6644 4140
rect 6420 4100 6644 4128
rect 6420 4088 6426 4100
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6914 4128 6920 4140
rect 6854 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 8220 4137 8248 4168
rect 9508 4168 9680 4196
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8478 4128 8484 4140
rect 8439 4100 8484 4128
rect 8205 4091 8263 4097
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2406 4060 2412 4072
rect 2004 4032 2412 4060
rect 2004 4020 2010 4032
rect 2406 4020 2412 4032
rect 2464 4060 2470 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2464 4032 2789 4060
rect 2464 4020 2470 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 2777 4023 2835 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5644 4060 5672 4088
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5644 4032 6101 4060
rect 5169 4023 5227 4029
rect 6089 4029 6101 4032
rect 6135 4060 6147 4063
rect 6454 4060 6460 4072
rect 6135 4032 6460 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 1486 3952 1492 4004
rect 1544 3992 1550 4004
rect 4890 3992 4896 4004
rect 1544 3964 4896 3992
rect 1544 3952 1550 3964
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 5184 3992 5212 4023
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 7926 4060 7932 4072
rect 7887 4032 7932 4060
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8220 4060 8248 4091
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 8386 4060 8392 4072
rect 8220 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8588 4060 8616 4091
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8720 4100 9045 4128
rect 8720 4088 8726 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9180 4100 9225 4128
rect 9180 4088 9186 4100
rect 8588 4032 8708 4060
rect 5902 3992 5908 4004
rect 5184 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 8680 3992 8708 4032
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 9508 4069 9536 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 11977 4199 12035 4205
rect 11977 4196 11989 4199
rect 10994 4168 11989 4196
rect 11977 4165 11989 4168
rect 12023 4165 12035 4199
rect 11977 4159 12035 4165
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 11480 4100 11621 4128
rect 11480 4088 11486 4100
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11609 4091 11667 4097
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 8812 4032 9505 4060
rect 8812 4020 8818 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9766 4060 9772 4072
rect 9727 4032 9772 4060
rect 9493 4023 9551 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 11624 4060 11652 4091
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12066 4128 12072 4140
rect 11979 4100 12072 4128
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12176 4128 12204 4236
rect 12802 4224 12808 4236
rect 12860 4264 12866 4276
rect 12897 4267 12955 4273
rect 12897 4264 12909 4267
rect 12860 4236 12909 4264
rect 12860 4224 12866 4236
rect 12897 4233 12909 4236
rect 12943 4264 12955 4267
rect 13081 4267 13139 4273
rect 13081 4264 13093 4267
rect 12943 4236 13093 4264
rect 12943 4233 12955 4236
rect 12897 4227 12955 4233
rect 13081 4233 13093 4236
rect 13127 4264 13139 4267
rect 13265 4267 13323 4273
rect 13265 4264 13277 4267
rect 13127 4236 13277 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 13265 4233 13277 4236
rect 13311 4233 13323 4267
rect 13265 4227 13323 4233
rect 12529 4199 12587 4205
rect 12529 4165 12541 4199
rect 12575 4196 12587 4199
rect 12618 4196 12624 4208
rect 12575 4168 12624 4196
rect 12575 4165 12587 4168
rect 12529 4159 12587 4165
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 12176 4100 12265 4128
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 12710 4128 12716 4140
rect 12671 4100 12716 4128
rect 12253 4091 12311 4097
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13538 4128 13544 4140
rect 13035 4100 13544 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 12084 4060 12112 4088
rect 11624 4032 12112 4060
rect 8938 3992 8944 4004
rect 8680 3964 8944 3992
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 1854 3924 1860 3936
rect 1811 3896 1860 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2590 3924 2596 3936
rect 1995 3896 2596 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8680 3924 8708 3964
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 9398 3992 9404 4004
rect 9359 3964 9404 3992
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 8168 3896 8708 3924
rect 8849 3927 8907 3933
rect 8168 3884 8174 3896
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9950 3924 9956 3936
rect 8895 3896 9956 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10192 3896 11253 3924
rect 10192 3884 10198 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 13538 3924 13544 3936
rect 13499 3896 13544 3924
rect 11241 3887 11299 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3720 2743 3723
rect 2958 3720 2964 3732
rect 2731 3692 2964 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 4028 3692 4077 3720
rect 4028 3680 4034 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 8662 3720 8668 3732
rect 4065 3683 4123 3689
rect 5184 3692 8668 3720
rect 1670 3652 1676 3664
rect 1631 3624 1676 3652
rect 1670 3612 1676 3624
rect 1728 3612 1734 3664
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3621 2927 3655
rect 3326 3652 3332 3664
rect 3287 3624 3332 3652
rect 2869 3615 2927 3621
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 2015 3587 2073 3593
rect 1636 3556 1900 3584
rect 1636 3544 1642 3556
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 1872 3525 1900 3556
rect 2015 3553 2027 3587
rect 2061 3584 2073 3587
rect 2590 3584 2596 3596
rect 2061 3556 2452 3584
rect 2551 3556 2596 3584
rect 2061 3553 2073 3556
rect 2015 3547 2073 3553
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2314 3516 2320 3528
rect 2271 3488 2320 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2424 3516 2452 3556
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 2884 3584 2912 3615
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 5184 3652 5212 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9306 3720 9312 3732
rect 9267 3692 9312 3720
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9766 3720 9772 3732
rect 9723 3692 9772 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10318 3720 10324 3732
rect 9876 3692 10324 3720
rect 3528 3624 5212 3652
rect 3528 3584 3556 3624
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 6273 3655 6331 3661
rect 5316 3624 5764 3652
rect 5316 3612 5322 3624
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 2884 3556 3556 3584
rect 3620 3556 5457 3584
rect 3620 3525 3648 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2424 3488 2513 3516
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3485 3663 3519
rect 4246 3516 4252 3528
rect 4207 3488 4252 3516
rect 3605 3479 3663 3485
rect 1412 3448 1440 3476
rect 3053 3451 3111 3457
rect 3053 3448 3065 3451
rect 1412 3420 3065 3448
rect 3053 3417 3065 3420
rect 3099 3417 3111 3451
rect 3436 3448 3464 3479
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4338 3476 4344 3528
rect 4396 3516 4402 3528
rect 4525 3519 4583 3525
rect 4396 3488 4441 3516
rect 4396 3476 4402 3488
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4540 3448 4568 3479
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5169 3519 5227 3525
rect 4672 3488 4717 3516
rect 4672 3476 4678 3488
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 4985 3451 5043 3457
rect 4985 3448 4997 3451
rect 3436 3420 4997 3448
rect 3053 3411 3111 3417
rect 4985 3417 4997 3420
rect 5031 3417 5043 3451
rect 5184 3448 5212 3479
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5534 3516 5540 3528
rect 5316 3488 5361 3516
rect 5495 3488 5540 3516
rect 5316 3476 5322 3488
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5736 3525 5764 3624
rect 6273 3621 6285 3655
rect 6319 3652 6331 3655
rect 7190 3652 7196 3664
rect 6319 3624 7196 3652
rect 6319 3621 6331 3624
rect 6273 3615 6331 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9876 3652 9904 3692
rect 10318 3680 10324 3692
rect 10376 3720 10382 3732
rect 11882 3720 11888 3732
rect 10376 3692 11888 3720
rect 10376 3680 10382 3692
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 12802 3680 12808 3692
rect 12860 3720 12866 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12860 3692 13001 3720
rect 12860 3680 12866 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 10042 3652 10048 3664
rect 8996 3624 9904 3652
rect 10003 3624 10048 3652
rect 8996 3612 9002 3624
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 6546 3584 6552 3596
rect 6196 3556 6552 3584
rect 6196 3525 6224 3556
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 6914 3584 6920 3596
rect 6871 3556 6920 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8754 3584 8760 3596
rect 8444 3556 8760 3584
rect 8444 3544 8450 3556
rect 8754 3544 8760 3556
rect 8812 3584 8818 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 8812 3556 10425 3584
rect 8812 3544 8818 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11480 3556 12480 3584
rect 11480 3544 11486 3556
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 5552 3448 5580 3476
rect 5184 3420 5580 3448
rect 4985 3411 5043 3417
rect 5736 3380 5764 3479
rect 6380 3448 6408 3479
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6512 3488 6557 3516
rect 6512 3476 6518 3488
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 9858 3516 9864 3528
rect 6696 3488 6741 3516
rect 9819 3488 9864 3516
rect 6696 3476 6702 3488
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 12452 3525 12480 3556
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 12802 3516 12808 3528
rect 12759 3488 12808 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 6822 3448 6828 3460
rect 6380 3420 6828 3448
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7926 3408 7932 3460
rect 7984 3408 7990 3460
rect 8481 3451 8539 3457
rect 8481 3417 8493 3451
rect 8527 3417 8539 3451
rect 8481 3411 8539 3417
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 10686 3448 10692 3460
rect 9539 3420 10548 3448
rect 10647 3420 10692 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 6914 3380 6920 3392
rect 5736 3352 6920 3380
rect 6914 3340 6920 3352
rect 6972 3380 6978 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6972 3352 7021 3380
rect 6972 3340 6978 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8496 3380 8524 3411
rect 7524 3352 8524 3380
rect 9309 3383 9367 3389
rect 7524 3340 7530 3352
rect 9309 3349 9321 3383
rect 9355 3380 9367 3383
rect 9582 3380 9588 3392
rect 9355 3352 9588 3380
rect 9355 3349 9367 3352
rect 9309 3343 9367 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10520 3380 10548 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 12345 3451 12403 3457
rect 12345 3448 12357 3451
rect 11914 3420 12357 3448
rect 12345 3417 12357 3420
rect 12391 3417 12403 3451
rect 12345 3411 12403 3417
rect 10594 3380 10600 3392
rect 10520 3352 10600 3380
rect 10594 3340 10600 3352
rect 10652 3380 10658 3392
rect 12161 3383 12219 3389
rect 12161 3380 12173 3383
rect 10652 3352 12173 3380
rect 10652 3340 10658 3352
rect 12161 3349 12173 3352
rect 12207 3349 12219 3383
rect 12161 3343 12219 3349
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 4614 3176 4620 3188
rect 3436 3148 4620 3176
rect 2866 3108 2872 3120
rect 1596 3080 2619 3108
rect 2779 3080 2872 3108
rect 1486 3040 1492 3052
rect 1447 3012 1492 3040
rect 1486 3000 1492 3012
rect 1544 3000 1550 3052
rect 1596 2981 1624 3080
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2498 3040 2504 3052
rect 1903 3012 2504 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2591 3040 2619 3080
rect 2866 3068 2872 3080
rect 2924 3108 2930 3120
rect 2961 3111 3019 3117
rect 2961 3108 2973 3111
rect 2924 3080 2973 3108
rect 2924 3068 2930 3080
rect 2961 3077 2973 3080
rect 3007 3077 3019 3111
rect 3234 3108 3240 3120
rect 3195 3080 3240 3108
rect 2961 3071 3019 3077
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 3436 3049 3464 3148
rect 4614 3136 4620 3148
rect 4672 3176 4678 3188
rect 5169 3179 5227 3185
rect 5169 3176 5181 3179
rect 4672 3148 5181 3176
rect 4672 3136 4678 3148
rect 5169 3145 5181 3148
rect 5215 3145 5227 3179
rect 5169 3139 5227 3145
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 6086 3176 6092 3188
rect 5316 3148 5764 3176
rect 6047 3148 6092 3176
rect 5316 3136 5322 3148
rect 3697 3111 3755 3117
rect 3697 3077 3709 3111
rect 3743 3108 3755 3111
rect 4893 3111 4951 3117
rect 3743 3080 4292 3108
rect 3743 3077 3755 3080
rect 3697 3071 3755 3077
rect 4264 3052 4292 3080
rect 4893 3077 4905 3111
rect 4939 3108 4951 3111
rect 4982 3108 4988 3120
rect 4939 3080 4988 3108
rect 4939 3077 4951 3080
rect 4893 3071 4951 3077
rect 3421 3043 3479 3049
rect 2591 3012 3000 3040
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1780 2972 1808 3000
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 1780 2944 2697 2972
rect 1581 2935 1639 2941
rect 2685 2941 2697 2944
rect 2731 2972 2743 2975
rect 2866 2972 2872 2984
rect 2731 2944 2872 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 2972 2972 3000 3012
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3651 3012 4169 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4172 2972 4200 3003
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4304 3012 4537 3040
rect 4304 3000 4310 3012
rect 4525 3009 4537 3012
rect 4571 3040 4583 3043
rect 4614 3040 4620 3052
rect 4571 3012 4620 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4338 2972 4344 2984
rect 2972 2944 3740 2972
rect 4172 2944 4344 2972
rect 3712 2904 3740 2944
rect 4338 2932 4344 2944
rect 4396 2972 4402 2984
rect 4706 2972 4712 2984
rect 4396 2944 4712 2972
rect 4396 2932 4402 2944
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4908 2904 4936 3071
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 5736 3117 5764 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7466 3176 7472 3188
rect 6696 3148 7328 3176
rect 7427 3148 7472 3176
rect 6696 3136 6702 3148
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 7098 3108 7104 3120
rect 5951 3080 7104 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 6380 3049 6408 3080
rect 7098 3068 7104 3080
rect 7156 3068 7162 3120
rect 7300 3108 7328 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8570 3176 8576 3188
rect 8220 3148 8576 3176
rect 8220 3108 8248 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9456 3148 10057 3176
rect 9456 3136 9462 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10594 3176 10600 3188
rect 10555 3148 10600 3176
rect 10045 3139 10103 3145
rect 8772 3108 8800 3136
rect 7300 3080 8248 3108
rect 8312 3080 8800 3108
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5316 3012 5365 3040
rect 5316 3000 5322 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6365 3003 6423 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7190 3040 7196 3052
rect 6972 3012 7017 3040
rect 7151 3012 7196 3040
rect 6972 3000 6978 3012
rect 7190 3000 7196 3012
rect 7248 3040 7254 3052
rect 7466 3040 7472 3052
rect 7248 3012 7472 3040
rect 7248 3000 7254 3012
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7944 3049 7972 3080
rect 8312 3052 8340 3080
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7929 3043 7987 3049
rect 7699 3012 7880 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 5500 2944 5549 2972
rect 5500 2932 5506 2944
rect 5537 2941 5549 2944
rect 5583 2972 5595 2975
rect 6564 2972 6592 3000
rect 5583 2944 6592 2972
rect 7009 2975 7067 2981
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 3712 2876 4936 2904
rect 2041 2839 2099 2845
rect 2041 2805 2053 2839
rect 2087 2836 2099 2839
rect 2590 2836 2596 2848
rect 2087 2808 2596 2836
rect 2087 2805 2099 2808
rect 2041 2799 2099 2805
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 5828 2836 5856 2944
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7561 2975 7619 2981
rect 7055 2944 7512 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7190 2904 7196 2916
rect 6871 2876 7196 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7484 2904 7512 2944
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7742 2972 7748 2984
rect 7607 2944 7748 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 7852 2972 7880 3012
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 8110 3040 8116 3052
rect 8071 3012 8116 3040
rect 7929 3003 7987 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8294 3040 8300 3052
rect 8207 3012 8300 3040
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 9674 3000 9680 3052
rect 9732 3000 9738 3052
rect 10060 3040 10088 3139
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 10686 3136 10692 3188
rect 10744 3176 10750 3188
rect 11057 3179 11115 3185
rect 11057 3176 11069 3179
rect 10744 3148 11069 3176
rect 10744 3136 10750 3148
rect 11057 3145 11069 3148
rect 11103 3145 11115 3179
rect 11057 3139 11115 3145
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11882 3176 11888 3188
rect 11379 3148 11888 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10060 3012 10701 3040
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11422 3040 11428 3052
rect 11020 3012 11428 3040
rect 11020 3000 11026 3012
rect 11422 3000 11428 3012
rect 11480 3040 11486 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11480 3012 11621 3040
rect 11480 3000 11486 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11609 3003 11667 3009
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12618 3040 12624 3052
rect 12579 3012 12624 3040
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 8128 2972 8156 3000
rect 7852 2944 8156 2972
rect 8202 2932 8208 2984
rect 8260 2932 8266 2984
rect 8570 2972 8576 2984
rect 8531 2944 8576 2972
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 10551 2944 11989 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 12710 2972 12716 2984
rect 12671 2944 12716 2972
rect 11977 2935 12035 2941
rect 8220 2904 8248 2932
rect 7484 2876 8248 2904
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5828 2808 5917 2836
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 10520 2836 10548 2935
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 11609 2907 11667 2913
rect 11609 2873 11621 2907
rect 11655 2904 11667 2907
rect 11698 2904 11704 2916
rect 11655 2876 11704 2904
rect 11655 2873 11667 2876
rect 11609 2867 11667 2873
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 6052 2808 10548 2836
rect 6052 2796 6058 2808
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 1489 2635 1547 2641
rect 1489 2601 1501 2635
rect 1535 2632 1547 2635
rect 2409 2635 2467 2641
rect 1535 2604 2176 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 1946 2428 1952 2440
rect 1811 2400 1952 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2148 2428 2176 2604
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2498 2632 2504 2644
rect 2455 2604 2504 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4706 2632 4712 2644
rect 4203 2604 4712 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5902 2632 5908 2644
rect 5552 2604 5908 2632
rect 4062 2564 4068 2576
rect 3252 2536 4068 2564
rect 3252 2508 3280 2536
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 5552 2564 5580 2604
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 8386 2632 8392 2644
rect 6236 2604 6868 2632
rect 8347 2604 8392 2632
rect 6236 2592 6242 2604
rect 5184 2536 5580 2564
rect 6840 2564 6868 2604
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8628 2604 8953 2632
rect 8628 2592 8634 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 8941 2595 8999 2601
rect 10318 2592 10324 2604
rect 10376 2632 10382 2644
rect 10686 2632 10692 2644
rect 10376 2604 10692 2632
rect 10376 2592 10382 2604
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 6840 2536 8432 2564
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 3234 2496 3240 2508
rect 2271 2468 2544 2496
rect 3147 2468 3240 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2516 2437 2544 2468
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 5184 2496 5212 2536
rect 3467 2468 5212 2496
rect 5537 2499 5595 2505
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 8294 2496 8300 2508
rect 5583 2468 8300 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 5264 2440 5316 2446
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2148 2400 2329 2428
rect 2041 2391 2099 2397
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 3789 2431 3847 2437
rect 3789 2430 3801 2431
rect 2501 2391 2559 2397
rect 3712 2402 3801 2430
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 2056 2360 2084 2391
rect 1627 2332 3188 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 3160 2301 3188 2332
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2096 2264 2789 2292
rect 2096 2252 2102 2264
rect 2777 2261 2789 2264
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2292 3203 2295
rect 3712 2292 3740 2402
rect 3789 2397 3801 2402
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4062 2428 4068 2440
rect 4019 2400 4068 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 5442 2428 5448 2440
rect 5399 2400 5448 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2428 8079 2431
rect 8067 2400 8248 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 5264 2382 5316 2388
rect 4614 2360 4620 2372
rect 4575 2332 4620 2360
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 5810 2360 5816 2372
rect 5771 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 6144 2332 6302 2360
rect 6144 2320 6150 2332
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7248 2332 8125 2360
rect 7248 2320 7254 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 7098 2292 7104 2304
rect 3191 2264 7104 2292
rect 3191 2261 3203 2264
rect 3145 2255 3203 2261
rect 7098 2252 7104 2264
rect 7156 2292 7162 2304
rect 7282 2292 7288 2304
rect 7156 2264 7288 2292
rect 7156 2252 7162 2264
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 7929 2295 7987 2301
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8018 2292 8024 2304
rect 7975 2264 8024 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 8220 2292 8248 2400
rect 8297 2363 8355 2369
rect 8297 2329 8309 2363
rect 8343 2360 8355 2363
rect 8404 2360 8432 2536
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 9548 2536 9904 2564
rect 9548 2524 9554 2536
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 8938 2496 8944 2508
rect 8711 2468 8944 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 9582 2496 9588 2508
rect 9495 2468 9588 2496
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9398 2428 9404 2440
rect 9355 2400 9404 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9600 2360 9628 2456
rect 9876 2437 9904 2536
rect 10336 2496 10364 2592
rect 12618 2564 12624 2576
rect 11716 2536 12624 2564
rect 10152 2468 10364 2496
rect 10689 2499 10747 2505
rect 10152 2437 10180 2468
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 11716 2496 11744 2536
rect 12618 2524 12624 2536
rect 12676 2564 12682 2576
rect 12676 2536 13216 2564
rect 12676 2524 12682 2536
rect 13188 2508 13216 2536
rect 10735 2468 11744 2496
rect 12161 2499 12219 2505
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 12161 2465 12173 2499
rect 12207 2496 12219 2499
rect 13170 2496 13176 2508
rect 12207 2468 12434 2496
rect 13083 2468 13176 2496
rect 12207 2465 12219 2468
rect 12161 2459 12219 2465
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 10137 2431 10195 2437
rect 10137 2397 10149 2431
rect 10183 2397 10195 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 10137 2391 10195 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 12406 2428 12434 2468
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 12716 2440 12768 2446
rect 12406 2400 12716 2428
rect 12716 2382 12768 2388
rect 8343 2332 8432 2360
rect 8496 2332 9720 2360
rect 8343 2329 8355 2332
rect 8297 2323 8355 2329
rect 8496 2292 8524 2332
rect 8220 2264 8524 2292
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9364 2264 9413 2292
rect 9364 2252 9370 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9692 2292 9720 2332
rect 11698 2320 11704 2372
rect 11756 2320 11762 2372
rect 12345 2363 12403 2369
rect 12345 2329 12357 2363
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 12360 2292 12388 2323
rect 9692 2264 12388 2292
rect 9401 2255 9459 2261
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 1946 2048 1952 2100
rect 2004 2088 2010 2100
rect 3234 2088 3240 2100
rect 2004 2060 3240 2088
rect 2004 2048 2010 2060
rect 3234 2048 3240 2060
rect 3292 2048 3298 2100
rect 3513 2091 3571 2097
rect 3513 2057 3525 2091
rect 3559 2088 3571 2091
rect 3602 2088 3608 2100
rect 3559 2060 3608 2088
rect 3559 2057 3571 2060
rect 3513 2051 3571 2057
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 5350 2048 5356 2100
rect 5408 2088 5414 2100
rect 5537 2091 5595 2097
rect 5537 2088 5549 2091
rect 5408 2060 5549 2088
rect 5408 2048 5414 2060
rect 5537 2057 5549 2060
rect 5583 2057 5595 2091
rect 6086 2088 6092 2100
rect 6047 2060 6092 2088
rect 5537 2051 5595 2057
rect 6086 2048 6092 2060
rect 6144 2048 6150 2100
rect 6454 2088 6460 2100
rect 6415 2060 6460 2088
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
rect 9398 2048 9404 2100
rect 9456 2088 9462 2100
rect 10229 2091 10287 2097
rect 10229 2088 10241 2091
rect 9456 2060 10241 2088
rect 9456 2048 9462 2060
rect 10229 2057 10241 2060
rect 10275 2057 10287 2091
rect 10229 2051 10287 2057
rect 10870 2048 10876 2100
rect 10928 2088 10934 2100
rect 10965 2091 11023 2097
rect 10965 2088 10977 2091
rect 10928 2060 10977 2088
rect 10928 2048 10934 2060
rect 10965 2057 10977 2060
rect 11011 2057 11023 2091
rect 10965 2051 11023 2057
rect 13170 2048 13176 2100
rect 13228 2088 13234 2100
rect 13265 2091 13323 2097
rect 13265 2088 13277 2091
rect 13228 2060 13277 2088
rect 13228 2048 13234 2060
rect 13265 2057 13277 2060
rect 13311 2057 13323 2091
rect 13265 2051 13323 2057
rect 4614 1980 4620 2032
rect 4672 1980 4678 2032
rect 6472 2020 6500 2048
rect 7834 2020 7840 2032
rect 5920 1992 6500 2020
rect 7682 1992 7840 2020
rect 3326 1952 3332 1964
rect 3239 1924 3332 1952
rect 3326 1912 3332 1924
rect 3384 1952 3390 1964
rect 3786 1952 3792 1964
rect 3384 1924 3792 1952
rect 3384 1912 3390 1924
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 5920 1961 5948 1992
rect 7834 1980 7840 1992
rect 7892 1980 7898 2032
rect 8018 1980 8024 2032
rect 8076 2020 8082 2032
rect 8113 2023 8171 2029
rect 8113 2020 8125 2023
rect 8076 1992 8125 2020
rect 8076 1980 8082 1992
rect 8113 1989 8125 1992
rect 8159 1989 8171 2023
rect 8113 1983 8171 1989
rect 10410 1980 10416 2032
rect 10468 2020 10474 2032
rect 10468 1992 11560 2020
rect 10468 1980 10474 1992
rect 5905 1955 5963 1961
rect 5905 1921 5917 1955
rect 5951 1921 5963 1955
rect 5905 1915 5963 1921
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 6638 1952 6644 1964
rect 6052 1924 6644 1952
rect 6052 1912 6058 1924
rect 6638 1912 6644 1924
rect 6696 1912 6702 1964
rect 10505 1955 10563 1961
rect 9890 1924 10456 1952
rect 2685 1887 2743 1893
rect 2685 1853 2697 1887
rect 2731 1884 2743 1887
rect 2774 1884 2780 1896
rect 2731 1856 2780 1884
rect 2731 1853 2743 1856
rect 2685 1847 2743 1853
rect 2774 1844 2780 1856
rect 2832 1844 2838 1896
rect 4062 1884 4068 1896
rect 4023 1856 4068 1884
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 8389 1887 8447 1893
rect 8389 1853 8401 1887
rect 8435 1884 8447 1887
rect 8478 1884 8484 1896
rect 8435 1856 8484 1884
rect 8435 1853 8447 1856
rect 8389 1847 8447 1853
rect 8478 1844 8484 1856
rect 8536 1844 8542 1896
rect 8754 1884 8760 1896
rect 8715 1856 8760 1884
rect 8754 1844 8760 1856
rect 8812 1844 8818 1896
rect 10428 1893 10456 1924
rect 10505 1921 10517 1955
rect 10551 1921 10563 1955
rect 10686 1952 10692 1964
rect 10647 1924 10692 1952
rect 10505 1915 10563 1921
rect 10413 1887 10471 1893
rect 10413 1853 10425 1887
rect 10459 1853 10471 1887
rect 10413 1847 10471 1853
rect 10520 1816 10548 1915
rect 10686 1912 10692 1924
rect 10744 1912 10750 1964
rect 10962 1952 10968 1964
rect 10923 1924 10968 1952
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 11532 1961 11560 1992
rect 12066 1980 12072 2032
rect 12124 2020 12130 2032
rect 12124 1992 12282 2020
rect 12124 1980 12130 1992
rect 11149 1955 11207 1961
rect 11149 1921 11161 1955
rect 11195 1921 11207 1955
rect 11149 1915 11207 1921
rect 11517 1955 11575 1961
rect 11517 1921 11529 1955
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 10962 1816 10968 1828
rect 10520 1788 10968 1816
rect 6546 1708 6552 1760
rect 6604 1748 6610 1760
rect 6641 1751 6699 1757
rect 6641 1748 6653 1751
rect 6604 1720 6653 1748
rect 6604 1708 6610 1720
rect 6641 1717 6653 1720
rect 6687 1748 6699 1751
rect 7098 1748 7104 1760
rect 6687 1720 7104 1748
rect 6687 1717 6699 1720
rect 6641 1711 6699 1717
rect 7098 1708 7104 1720
rect 7156 1708 7162 1760
rect 9490 1708 9496 1760
rect 9548 1748 9554 1760
rect 10520 1748 10548 1788
rect 10962 1776 10968 1788
rect 11020 1776 11026 1828
rect 9548 1720 10548 1748
rect 9548 1708 9554 1720
rect 10686 1708 10692 1760
rect 10744 1748 10750 1760
rect 11164 1748 11192 1915
rect 11790 1884 11796 1896
rect 11751 1856 11796 1884
rect 11790 1844 11796 1856
rect 11848 1844 11854 1896
rect 11606 1748 11612 1760
rect 10744 1720 11612 1748
rect 10744 1708 10750 1720
rect 11606 1708 11612 1720
rect 11664 1748 11670 1760
rect 11974 1748 11980 1760
rect 11664 1720 11980 1748
rect 11664 1708 11670 1720
rect 11974 1708 11980 1720
rect 12032 1708 12038 1760
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 2222 1504 2228 1556
rect 2280 1544 2286 1556
rect 3881 1547 3939 1553
rect 3881 1544 3893 1547
rect 2280 1516 3893 1544
rect 2280 1504 2286 1516
rect 3881 1513 3893 1516
rect 3927 1513 3939 1547
rect 3881 1507 3939 1513
rect 4062 1504 4068 1556
rect 4120 1544 4126 1556
rect 4709 1547 4767 1553
rect 4709 1544 4721 1547
rect 4120 1516 4721 1544
rect 4120 1504 4126 1516
rect 4709 1513 4721 1516
rect 4755 1513 4767 1547
rect 4709 1507 4767 1513
rect 5629 1547 5687 1553
rect 5629 1513 5641 1547
rect 5675 1544 5687 1547
rect 5810 1544 5816 1556
rect 5675 1516 5816 1544
rect 5675 1513 5687 1516
rect 5629 1507 5687 1513
rect 5810 1504 5816 1516
rect 5868 1504 5874 1556
rect 8481 1547 8539 1553
rect 8481 1544 8493 1547
rect 6656 1516 7052 1544
rect 3234 1436 3240 1488
rect 3292 1476 3298 1488
rect 3513 1479 3571 1485
rect 3513 1476 3525 1479
rect 3292 1448 3525 1476
rect 3292 1436 3298 1448
rect 3513 1445 3525 1448
rect 3559 1445 3571 1479
rect 5902 1476 5908 1488
rect 3513 1439 3571 1445
rect 5644 1448 5908 1476
rect 2038 1408 2044 1420
rect 1999 1380 2044 1408
rect 2038 1368 2044 1380
rect 2096 1368 2102 1420
rect 2590 1368 2596 1420
rect 2648 1408 2654 1420
rect 2648 1380 3280 1408
rect 2648 1368 2654 1380
rect 1486 1340 1492 1352
rect 1447 1312 1492 1340
rect 1486 1300 1492 1312
rect 1544 1300 1550 1352
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1309 1823 1343
rect 3252 1340 3280 1380
rect 3602 1368 3608 1420
rect 3660 1408 3666 1420
rect 5353 1411 5411 1417
rect 3660 1380 4108 1408
rect 3660 1368 3666 1380
rect 3789 1343 3847 1349
rect 3789 1340 3801 1343
rect 3252 1312 3801 1340
rect 1765 1303 1823 1309
rect 3789 1309 3801 1312
rect 3835 1309 3847 1343
rect 3970 1340 3976 1352
rect 3931 1312 3976 1340
rect 3789 1303 3847 1309
rect 1780 1204 1808 1303
rect 3970 1300 3976 1312
rect 4028 1300 4034 1352
rect 4080 1340 4108 1380
rect 5353 1377 5365 1411
rect 5399 1408 5411 1411
rect 5644 1408 5672 1448
rect 5902 1436 5908 1448
rect 5960 1436 5966 1488
rect 6546 1408 6552 1420
rect 5399 1380 5672 1408
rect 5828 1380 6552 1408
rect 5399 1377 5411 1380
rect 5353 1371 5411 1377
rect 4249 1343 4307 1349
rect 4249 1340 4261 1343
rect 4080 1312 4261 1340
rect 4249 1309 4261 1312
rect 4295 1309 4307 1343
rect 4430 1340 4436 1352
rect 4391 1312 4436 1340
rect 4249 1303 4307 1309
rect 4430 1300 4436 1312
rect 4488 1300 4494 1352
rect 4614 1340 4620 1352
rect 4575 1312 4620 1340
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1340 5135 1343
rect 5442 1340 5448 1352
rect 5123 1312 5448 1340
rect 5123 1309 5135 1312
rect 5077 1303 5135 1309
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 5537 1343 5595 1349
rect 5537 1309 5549 1343
rect 5583 1309 5595 1343
rect 5537 1303 5595 1309
rect 5169 1275 5227 1281
rect 3266 1244 5120 1272
rect 3326 1204 3332 1216
rect 1780 1176 3332 1204
rect 3326 1164 3332 1176
rect 3384 1164 3390 1216
rect 5092 1204 5120 1244
rect 5169 1241 5181 1275
rect 5215 1272 5227 1275
rect 5350 1272 5356 1284
rect 5215 1244 5356 1272
rect 5215 1241 5227 1244
rect 5169 1235 5227 1241
rect 5350 1232 5356 1244
rect 5408 1232 5414 1284
rect 5552 1272 5580 1303
rect 5828 1272 5856 1380
rect 6546 1368 6552 1380
rect 6604 1368 6610 1420
rect 5902 1300 5908 1352
rect 5960 1340 5966 1352
rect 6181 1343 6239 1349
rect 5960 1312 6005 1340
rect 5960 1300 5966 1312
rect 6181 1309 6193 1343
rect 6227 1340 6239 1343
rect 6656 1340 6684 1516
rect 7024 1476 7052 1516
rect 8404 1516 8493 1544
rect 7558 1476 7564 1488
rect 7024 1448 7564 1476
rect 7558 1436 7564 1448
rect 7616 1436 7622 1488
rect 7006 1368 7012 1420
rect 7064 1408 7070 1420
rect 7193 1411 7251 1417
rect 7193 1408 7205 1411
rect 7064 1380 7205 1408
rect 7064 1368 7070 1380
rect 7193 1377 7205 1380
rect 7239 1408 7251 1411
rect 7282 1408 7288 1420
rect 7239 1380 7288 1408
rect 7239 1377 7251 1380
rect 7193 1371 7251 1377
rect 7282 1368 7288 1380
rect 7340 1368 7346 1420
rect 7466 1368 7472 1420
rect 7524 1408 7530 1420
rect 7653 1411 7711 1417
rect 7653 1408 7665 1411
rect 7524 1380 7665 1408
rect 7524 1368 7530 1380
rect 7653 1377 7665 1380
rect 7699 1377 7711 1411
rect 7653 1371 7711 1377
rect 7834 1368 7840 1420
rect 7892 1408 7898 1420
rect 7929 1411 7987 1417
rect 7929 1408 7941 1411
rect 7892 1380 7941 1408
rect 7892 1368 7898 1380
rect 7929 1377 7941 1380
rect 7975 1377 7987 1411
rect 8404 1408 8432 1516
rect 8481 1513 8493 1516
rect 8527 1544 8539 1547
rect 9490 1544 9496 1556
rect 8527 1516 9496 1544
rect 8527 1513 8539 1516
rect 8481 1507 8539 1513
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 9756 1547 9814 1553
rect 9756 1513 9768 1547
rect 9802 1544 9814 1547
rect 11146 1544 11152 1556
rect 9802 1516 11152 1544
rect 9802 1513 9814 1516
rect 9756 1507 9814 1513
rect 11146 1504 11152 1516
rect 11204 1504 11210 1556
rect 11241 1547 11299 1553
rect 11241 1513 11253 1547
rect 11287 1544 11299 1547
rect 11790 1544 11796 1556
rect 11287 1516 11796 1544
rect 11287 1513 11299 1516
rect 11241 1507 11299 1513
rect 11790 1504 11796 1516
rect 11848 1504 11854 1556
rect 11974 1504 11980 1556
rect 12032 1544 12038 1556
rect 12529 1547 12587 1553
rect 12529 1544 12541 1547
rect 12032 1516 12541 1544
rect 12032 1504 12038 1516
rect 8754 1436 8760 1488
rect 8812 1476 8818 1488
rect 8941 1479 8999 1485
rect 8941 1476 8953 1479
rect 8812 1448 8953 1476
rect 8812 1436 8818 1448
rect 8941 1445 8953 1448
rect 8987 1445 8999 1479
rect 8941 1439 8999 1445
rect 7929 1371 7987 1377
rect 8128 1380 8432 1408
rect 8128 1352 8156 1380
rect 8478 1368 8484 1420
rect 8536 1408 8542 1420
rect 9493 1411 9551 1417
rect 9493 1408 9505 1411
rect 8536 1380 9505 1408
rect 8536 1368 8542 1380
rect 9493 1377 9505 1380
rect 9539 1408 9551 1411
rect 10410 1408 10416 1420
rect 9539 1380 10416 1408
rect 9539 1377 9551 1380
rect 9493 1371 9551 1377
rect 10410 1368 10416 1380
rect 10468 1368 10474 1420
rect 10962 1368 10968 1420
rect 11020 1408 11026 1420
rect 11020 1380 12204 1408
rect 11020 1368 11026 1380
rect 7098 1340 7104 1352
rect 6227 1312 6684 1340
rect 7059 1312 7104 1340
rect 6227 1309 6239 1312
rect 6181 1303 6239 1309
rect 7098 1300 7104 1312
rect 7156 1300 7162 1352
rect 8110 1340 8116 1352
rect 8071 1312 8116 1340
rect 8110 1300 8116 1312
rect 8168 1300 8174 1352
rect 8202 1300 8208 1352
rect 8260 1340 8266 1352
rect 8297 1343 8355 1349
rect 8297 1340 8309 1343
rect 8260 1312 8309 1340
rect 8260 1300 8266 1312
rect 8297 1309 8309 1312
rect 8343 1309 8355 1343
rect 8297 1303 8355 1309
rect 8389 1343 8447 1349
rect 8389 1309 8401 1343
rect 8435 1309 8447 1343
rect 8389 1303 8447 1309
rect 8665 1343 8723 1349
rect 8665 1309 8677 1343
rect 8711 1340 8723 1343
rect 8938 1340 8944 1352
rect 8711 1312 8944 1340
rect 8711 1309 8723 1312
rect 8665 1303 8723 1309
rect 5552 1244 5856 1272
rect 5920 1244 6679 1272
rect 5920 1204 5948 1244
rect 5092 1176 5948 1204
rect 6454 1164 6460 1216
rect 6512 1204 6518 1216
rect 6651 1204 6679 1244
rect 8018 1232 8024 1284
rect 8076 1272 8082 1284
rect 8404 1272 8432 1303
rect 8938 1300 8944 1312
rect 8996 1300 9002 1352
rect 9125 1343 9183 1349
rect 9125 1309 9137 1343
rect 9171 1340 9183 1343
rect 9398 1340 9404 1352
rect 9171 1312 9404 1340
rect 9171 1309 9183 1312
rect 9125 1303 9183 1309
rect 9398 1300 9404 1312
rect 9456 1300 9462 1352
rect 10870 1300 10876 1352
rect 10928 1300 10934 1352
rect 11606 1340 11612 1352
rect 11567 1312 11612 1340
rect 11606 1300 11612 1312
rect 11664 1300 11670 1352
rect 11808 1349 11836 1380
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1309 11851 1343
rect 11793 1303 11851 1309
rect 11977 1343 12035 1349
rect 11977 1309 11989 1343
rect 12023 1340 12035 1343
rect 12066 1340 12072 1352
rect 12023 1312 12072 1340
rect 12023 1309 12035 1312
rect 11977 1303 12035 1309
rect 12066 1300 12072 1312
rect 12124 1300 12130 1352
rect 12176 1349 12204 1380
rect 12360 1349 12388 1516
rect 12529 1513 12541 1516
rect 12575 1544 12587 1547
rect 12713 1547 12771 1553
rect 12713 1544 12725 1547
rect 12575 1516 12725 1544
rect 12575 1513 12587 1516
rect 12529 1507 12587 1513
rect 12713 1513 12725 1516
rect 12759 1544 12771 1547
rect 13081 1547 13139 1553
rect 13081 1544 13093 1547
rect 12759 1516 13093 1544
rect 12759 1513 12771 1516
rect 12713 1507 12771 1513
rect 13081 1513 13093 1516
rect 13127 1513 13139 1547
rect 13081 1507 13139 1513
rect 12161 1343 12219 1349
rect 12161 1309 12173 1343
rect 12207 1309 12219 1343
rect 12161 1303 12219 1309
rect 12345 1343 12403 1349
rect 12345 1309 12357 1343
rect 12391 1309 12403 1343
rect 12345 1303 12403 1309
rect 8076 1244 8432 1272
rect 9309 1275 9367 1281
rect 8076 1232 8082 1244
rect 9309 1241 9321 1275
rect 9355 1272 9367 1275
rect 9490 1272 9496 1284
rect 9355 1244 9496 1272
rect 9355 1241 9367 1244
rect 9309 1235 9367 1241
rect 9490 1232 9496 1244
rect 9548 1232 9554 1284
rect 11146 1232 11152 1284
rect 11204 1272 11210 1284
rect 11204 1244 12296 1272
rect 11204 1232 11210 1244
rect 12161 1207 12219 1213
rect 12161 1204 12173 1207
rect 6512 1176 6557 1204
rect 6651 1176 12173 1204
rect 6512 1164 6518 1176
rect 12161 1173 12173 1176
rect 12207 1173 12219 1207
rect 12268 1204 12296 1244
rect 12897 1207 12955 1213
rect 12897 1204 12909 1207
rect 12268 1176 12909 1204
rect 12161 1167 12219 1173
rect 12897 1173 12909 1176
rect 12943 1173 12955 1207
rect 12897 1167 12955 1173
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
rect 3694 960 3700 1012
rect 3752 1000 3758 1012
rect 6454 1000 6460 1012
rect 3752 972 6460 1000
rect 3752 960 3758 972
rect 6454 960 6460 972
rect 6512 1000 6518 1012
rect 8018 1000 8024 1012
rect 6512 972 8024 1000
rect 6512 960 6518 972
rect 8018 960 8024 972
rect 8076 960 8082 1012
rect 4430 892 4436 944
rect 4488 932 4494 944
rect 5994 932 6000 944
rect 4488 904 6000 932
rect 4488 892 4494 904
rect 5994 892 6000 904
rect 6052 932 6058 944
rect 8110 932 8116 944
rect 6052 904 8116 932
rect 6052 892 6058 904
rect 8110 892 8116 904
rect 8168 892 8174 944
<< via1 >>
rect 9404 13812 9456 13864
rect 12072 13812 12124 13864
rect 2044 13744 2096 13796
rect 9956 13744 10008 13796
rect 1676 13676 1728 13728
rect 7104 13676 7156 13728
rect 7380 13676 7432 13728
rect 7472 13676 7524 13728
rect 11796 13676 11848 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 572 13472 624 13524
rect 4068 13404 4120 13456
rect 4712 13336 4764 13388
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 2320 13268 2372 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 3976 13268 4028 13320
rect 4620 13311 4672 13320
rect 1400 13200 1452 13252
rect 2136 13243 2188 13252
rect 2136 13209 2145 13243
rect 2145 13209 2179 13243
rect 2179 13209 2188 13243
rect 2136 13200 2188 13209
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 4160 13200 4212 13252
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 6644 13404 6696 13456
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 6092 13311 6144 13320
rect 5080 13243 5132 13252
rect 5080 13209 5089 13243
rect 5089 13209 5123 13243
rect 5123 13209 5132 13243
rect 5080 13200 5132 13209
rect 5724 13243 5776 13252
rect 5724 13209 5733 13243
rect 5733 13209 5767 13243
rect 5767 13209 5776 13243
rect 5724 13200 5776 13209
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7380 13472 7432 13524
rect 9404 13472 9456 13524
rect 11336 13472 11388 13524
rect 9312 13404 9364 13456
rect 9496 13404 9548 13456
rect 9036 13336 9088 13388
rect 8116 13268 8168 13320
rect 8852 13268 8904 13320
rect 6920 13243 6972 13252
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 2780 13132 2832 13184
rect 2872 13132 2924 13184
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 6920 13209 6929 13243
rect 6929 13209 6963 13243
rect 6963 13209 6972 13243
rect 6920 13200 6972 13209
rect 7564 13243 7616 13252
rect 6828 13132 6880 13184
rect 7564 13209 7573 13243
rect 7573 13209 7607 13243
rect 7607 13209 7616 13243
rect 7564 13200 7616 13209
rect 8760 13243 8812 13252
rect 8760 13209 8769 13243
rect 8769 13209 8803 13243
rect 8803 13209 8812 13243
rect 9956 13243 10008 13252
rect 8760 13200 8812 13209
rect 7380 13132 7432 13184
rect 9496 13132 9548 13184
rect 9956 13209 9965 13243
rect 9965 13209 9999 13243
rect 9999 13209 10008 13243
rect 9956 13200 10008 13209
rect 10232 13268 10284 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 12072 13311 12124 13320
rect 10876 13200 10928 13252
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 11612 13243 11664 13252
rect 11612 13209 11621 13243
rect 11621 13209 11655 13243
rect 11655 13209 11664 13243
rect 11612 13200 11664 13209
rect 11796 13200 11848 13252
rect 12624 13243 12676 13252
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 12624 13200 12676 13209
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 13360 13243 13412 13252
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13360 13200 13412 13209
rect 13176 13132 13228 13184
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 1400 12971 1452 12980
rect 1400 12937 1409 12971
rect 1409 12937 1443 12971
rect 1443 12937 1452 12971
rect 1400 12928 1452 12937
rect 2780 12928 2832 12980
rect 4436 12928 4488 12980
rect 7012 12928 7064 12980
rect 7288 12928 7340 12980
rect 9036 12928 9088 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 2320 12835 2372 12844
rect 1400 12724 1452 12776
rect 2320 12801 2329 12835
rect 2329 12801 2363 12835
rect 2363 12801 2372 12835
rect 2320 12792 2372 12801
rect 2872 12792 2924 12844
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 5080 12860 5132 12912
rect 7564 12860 7616 12912
rect 5540 12792 5592 12844
rect 5632 12792 5684 12844
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 3976 12724 4028 12776
rect 3240 12656 3292 12708
rect 4804 12656 4856 12708
rect 4988 12588 5040 12640
rect 6644 12792 6696 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 7012 12835 7064 12844
rect 6828 12792 6880 12801
rect 7012 12801 7015 12835
rect 7015 12801 7064 12835
rect 7012 12792 7064 12801
rect 7380 12792 7432 12844
rect 6920 12656 6972 12708
rect 8944 12860 8996 12912
rect 8116 12835 8168 12844
rect 7380 12656 7432 12708
rect 6828 12588 6880 12640
rect 7472 12588 7524 12640
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9680 12860 9732 12912
rect 9128 12792 9180 12801
rect 9404 12792 9456 12844
rect 10324 12928 10376 12980
rect 10968 12928 11020 12980
rect 12624 12860 12676 12912
rect 10876 12792 10928 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 12164 12792 12216 12844
rect 11152 12724 11204 12776
rect 11888 12724 11940 12776
rect 8484 12656 8536 12708
rect 8852 12656 8904 12708
rect 10048 12656 10100 12708
rect 10876 12656 10928 12708
rect 11060 12656 11112 12708
rect 12900 12656 12952 12708
rect 9128 12588 9180 12640
rect 9588 12588 9640 12640
rect 10416 12588 10468 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 6736 12384 6788 12436
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 8484 12384 8536 12436
rect 8760 12384 8812 12436
rect 9128 12384 9180 12436
rect 10416 12427 10468 12436
rect 2872 12359 2924 12368
rect 2872 12325 2881 12359
rect 2881 12325 2915 12359
rect 2915 12325 2924 12359
rect 2872 12316 2924 12325
rect 3608 12316 3660 12368
rect 4620 12316 4672 12368
rect 2044 12248 2096 12300
rect 3516 12291 3568 12300
rect 3516 12257 3525 12291
rect 3525 12257 3559 12291
rect 3559 12257 3568 12291
rect 3516 12248 3568 12257
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 1584 12112 1636 12164
rect 2320 12155 2372 12164
rect 2320 12121 2329 12155
rect 2329 12121 2363 12155
rect 2363 12121 2372 12155
rect 2320 12112 2372 12121
rect 2688 12155 2740 12164
rect 2688 12121 2697 12155
rect 2697 12121 2731 12155
rect 2731 12121 2740 12155
rect 2688 12112 2740 12121
rect 3700 12180 3752 12232
rect 4344 12223 4396 12232
rect 4344 12189 4353 12223
rect 4353 12189 4387 12223
rect 4387 12189 4396 12223
rect 4344 12180 4396 12189
rect 3976 12112 4028 12164
rect 4896 12155 4948 12164
rect 4896 12121 4905 12155
rect 4905 12121 4939 12155
rect 4939 12121 4948 12155
rect 4896 12112 4948 12121
rect 2780 12044 2832 12096
rect 3608 12044 3660 12096
rect 5264 12316 5316 12368
rect 8576 12316 8628 12368
rect 9496 12359 9548 12368
rect 6828 12248 6880 12300
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 6460 12180 6512 12232
rect 7104 12223 7156 12232
rect 7104 12189 7107 12223
rect 7107 12189 7156 12223
rect 7104 12180 7156 12189
rect 8392 12223 8444 12232
rect 8392 12189 8396 12223
rect 8396 12189 8430 12223
rect 8430 12189 8444 12223
rect 8392 12180 8444 12189
rect 8852 12180 8904 12232
rect 9036 12180 9088 12232
rect 9496 12325 9505 12359
rect 9505 12325 9539 12359
rect 9539 12325 9548 12359
rect 9496 12316 9548 12325
rect 10048 12359 10100 12368
rect 10048 12325 10057 12359
rect 10057 12325 10091 12359
rect 10091 12325 10100 12359
rect 10048 12316 10100 12325
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 14372 12384 14424 12436
rect 13268 12359 13320 12368
rect 13268 12325 13277 12359
rect 13277 12325 13311 12359
rect 13311 12325 13320 12359
rect 13268 12316 13320 12325
rect 9312 12248 9364 12300
rect 10600 12248 10652 12300
rect 11796 12248 11848 12300
rect 5632 12112 5684 12164
rect 6368 12155 6420 12164
rect 6368 12121 6377 12155
rect 6377 12121 6411 12155
rect 6411 12121 6420 12155
rect 6368 12112 6420 12121
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 6736 12112 6788 12164
rect 7564 12155 7616 12164
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 7288 12044 7340 12096
rect 7840 12112 7892 12164
rect 8576 12155 8628 12164
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 8944 12112 8996 12164
rect 9680 12112 9732 12164
rect 11612 12223 11664 12232
rect 10508 12112 10560 12164
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 11244 12112 11296 12164
rect 12072 12112 12124 12164
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 9036 12044 9088 12096
rect 9496 12044 9548 12096
rect 10048 12044 10100 12096
rect 10324 12044 10376 12096
rect 10968 12044 11020 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 2228 11815 2280 11824
rect 2228 11781 2237 11815
rect 2237 11781 2271 11815
rect 2271 11781 2280 11815
rect 2228 11772 2280 11781
rect 2320 11815 2372 11824
rect 2320 11781 2329 11815
rect 2329 11781 2363 11815
rect 2363 11781 2372 11815
rect 2320 11772 2372 11781
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 2964 11840 3016 11892
rect 3608 11772 3660 11824
rect 4804 11772 4856 11824
rect 2872 11704 2924 11756
rect 4160 11704 4212 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 3424 11636 3476 11688
rect 4620 11636 4672 11688
rect 5908 11840 5960 11892
rect 6368 11840 6420 11892
rect 6920 11883 6972 11892
rect 5632 11772 5684 11824
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 6552 11815 6604 11824
rect 2688 11568 2740 11620
rect 4712 11611 4764 11620
rect 2780 11500 2832 11552
rect 4712 11577 4721 11611
rect 4721 11577 4755 11611
rect 4755 11577 4764 11611
rect 4712 11568 4764 11577
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5724 11704 5776 11756
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6184 11747 6236 11756
rect 6184 11713 6193 11747
rect 6193 11713 6227 11747
rect 6227 11713 6236 11747
rect 6552 11781 6561 11815
rect 6561 11781 6595 11815
rect 6595 11781 6604 11815
rect 6552 11772 6604 11781
rect 7288 11772 7340 11824
rect 6184 11704 6236 11713
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 7748 11815 7800 11824
rect 7748 11781 7757 11815
rect 7757 11781 7791 11815
rect 7791 11781 7800 11815
rect 10692 11840 10744 11892
rect 11612 11883 11664 11892
rect 7748 11772 7800 11781
rect 10508 11772 10560 11824
rect 11612 11849 11621 11883
rect 11621 11849 11655 11883
rect 11655 11849 11664 11883
rect 11612 11840 11664 11849
rect 8024 11704 8076 11756
rect 6552 11568 6604 11620
rect 7196 11568 7248 11620
rect 4804 11500 4856 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 6460 11500 6512 11552
rect 7288 11500 7340 11552
rect 7564 11500 7616 11552
rect 8116 11568 8168 11620
rect 8484 11704 8536 11756
rect 8760 11704 8812 11756
rect 8944 11704 8996 11756
rect 9680 11747 9732 11756
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 8208 11500 8260 11552
rect 8392 11611 8444 11620
rect 8392 11577 8401 11611
rect 8401 11577 8435 11611
rect 8435 11577 8444 11611
rect 8392 11568 8444 11577
rect 8944 11568 8996 11620
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 10048 11704 10100 11756
rect 11152 11772 11204 11824
rect 11428 11772 11480 11824
rect 13268 11815 13320 11824
rect 13268 11781 13277 11815
rect 13277 11781 13311 11815
rect 13311 11781 13320 11815
rect 13268 11772 13320 11781
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 10876 11704 10928 11756
rect 11336 11704 11388 11756
rect 10508 11636 10560 11688
rect 8760 11500 8812 11552
rect 9128 11500 9180 11552
rect 10416 11568 10468 11620
rect 11704 11747 11756 11756
rect 11704 11713 11737 11747
rect 11737 11713 11756 11747
rect 11704 11704 11756 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12808 11704 12860 11756
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 11520 11568 11572 11620
rect 12716 11636 12768 11688
rect 11980 11568 12032 11620
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11336 11500 11388 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 6828 11296 6880 11348
rect 7104 11296 7156 11348
rect 8024 11296 8076 11348
rect 2688 11271 2740 11280
rect 2688 11237 2697 11271
rect 2697 11237 2731 11271
rect 2731 11237 2740 11271
rect 2688 11228 2740 11237
rect 4804 11228 4856 11280
rect 1676 11160 1728 11212
rect 6184 11203 6236 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 3240 11092 3292 11144
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 7012 11228 7064 11280
rect 7104 11160 7156 11212
rect 4068 11092 4120 11144
rect 4252 11092 4304 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 5172 11092 5224 11144
rect 5448 11092 5500 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 6552 11092 6604 11144
rect 7840 11228 7892 11280
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 10140 11296 10192 11348
rect 10692 11296 10744 11348
rect 10876 11296 10928 11348
rect 11152 11296 11204 11348
rect 9404 11228 9456 11280
rect 9864 11228 9916 11280
rect 7288 11160 7340 11212
rect 8116 11160 8168 11212
rect 8208 11160 8260 11212
rect 11612 11228 11664 11280
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 4896 11024 4948 11076
rect 2964 10956 3016 11008
rect 5540 10956 5592 11008
rect 6000 10956 6052 11008
rect 7288 11024 7340 11076
rect 6920 10956 6972 11008
rect 7932 10956 7984 11008
rect 8116 10956 8168 11008
rect 9036 11024 9088 11076
rect 9220 11024 9272 11076
rect 9772 11135 9824 11144
rect 9772 11101 9780 11135
rect 9780 11101 9814 11135
rect 9814 11101 9824 11135
rect 9772 11092 9824 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10048 11092 10100 11144
rect 9496 11024 9548 11076
rect 10784 11092 10836 11144
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 12072 11296 12124 11348
rect 11796 11092 11848 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 12716 11296 12768 11348
rect 11980 11092 12032 11101
rect 12808 11092 12860 11144
rect 9588 10956 9640 11008
rect 10048 10956 10100 11008
rect 12440 11024 12492 11076
rect 12900 11024 12952 11076
rect 11152 10956 11204 11008
rect 12716 10956 12768 11008
rect 13452 10999 13504 11008
rect 13452 10965 13461 10999
rect 13461 10965 13495 10999
rect 13495 10965 13504 10999
rect 13452 10956 13504 10965
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 3516 10752 3568 10804
rect 4620 10752 4672 10804
rect 6276 10752 6328 10804
rect 2504 10684 2556 10736
rect 3700 10684 3752 10736
rect 4252 10727 4304 10736
rect 4252 10693 4261 10727
rect 4261 10693 4295 10727
rect 4295 10693 4304 10727
rect 4252 10684 4304 10693
rect 5080 10684 5132 10736
rect 7012 10727 7064 10736
rect 7012 10693 7021 10727
rect 7021 10693 7055 10727
rect 7055 10693 7064 10727
rect 7012 10684 7064 10693
rect 7104 10684 7156 10736
rect 1584 10659 1636 10668
rect 1584 10625 1633 10659
rect 1633 10625 1636 10659
rect 1768 10659 1820 10668
rect 1584 10616 1636 10625
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 3240 10616 3292 10668
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 3332 10548 3384 10600
rect 5908 10616 5960 10668
rect 7564 10616 7616 10668
rect 7932 10684 7984 10736
rect 8208 10727 8260 10736
rect 8208 10693 8217 10727
rect 8217 10693 8251 10727
rect 8251 10693 8260 10727
rect 8208 10684 8260 10693
rect 8760 10727 8812 10736
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 9036 10684 9088 10736
rect 6736 10548 6788 10600
rect 8760 10548 8812 10600
rect 9772 10727 9824 10736
rect 9772 10693 9781 10727
rect 9781 10693 9815 10727
rect 9815 10693 9824 10727
rect 9772 10684 9824 10693
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 1584 10480 1636 10532
rect 6184 10480 6236 10532
rect 6552 10480 6604 10532
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 5080 10412 5132 10464
rect 5724 10412 5776 10464
rect 6368 10412 6420 10464
rect 7380 10480 7432 10532
rect 7564 10480 7616 10532
rect 11336 10752 11388 10804
rect 11520 10752 11572 10804
rect 11980 10752 12032 10804
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 12716 10727 12768 10736
rect 12716 10693 12725 10727
rect 12725 10693 12759 10727
rect 12759 10693 12768 10727
rect 12716 10684 12768 10693
rect 13452 10727 13504 10736
rect 13452 10693 13461 10727
rect 13461 10693 13495 10727
rect 13495 10693 13504 10727
rect 13452 10684 13504 10693
rect 10416 10616 10468 10625
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 11244 10548 11296 10600
rect 11612 10616 11664 10668
rect 13176 10616 13228 10668
rect 12072 10548 12124 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 10324 10480 10376 10532
rect 10600 10523 10652 10532
rect 10600 10489 10609 10523
rect 10609 10489 10643 10523
rect 10643 10489 10652 10523
rect 10600 10480 10652 10489
rect 6920 10412 6972 10464
rect 8852 10412 8904 10464
rect 9128 10412 9180 10464
rect 9404 10412 9456 10464
rect 9588 10412 9640 10464
rect 11704 10412 11756 10464
rect 13268 10480 13320 10532
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 1768 10208 1820 10260
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3792 10208 3844 10260
rect 5448 10208 5500 10260
rect 5540 10208 5592 10260
rect 7288 10208 7340 10260
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 7656 10208 7708 10260
rect 8484 10208 8536 10260
rect 9036 10208 9088 10260
rect 10416 10208 10468 10260
rect 11336 10208 11388 10260
rect 11428 10208 11480 10260
rect 2504 10140 2556 10192
rect 4988 10140 5040 10192
rect 1860 10072 1912 10124
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 3148 10004 3200 10056
rect 3608 10004 3660 10056
rect 6092 10072 6144 10124
rect 7104 10140 7156 10192
rect 13268 10183 13320 10192
rect 4528 9979 4580 9988
rect 4528 9945 4537 9979
rect 4537 9945 4571 9979
rect 4571 9945 4580 9979
rect 4528 9936 4580 9945
rect 5080 9979 5132 9988
rect 5080 9945 5089 9979
rect 5089 9945 5123 9979
rect 5123 9945 5132 9979
rect 5080 9936 5132 9945
rect 6276 10047 6328 10056
rect 6276 10013 6290 10047
rect 6290 10013 6324 10047
rect 6324 10013 6328 10047
rect 6276 10004 6328 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 5540 9936 5592 9988
rect 5816 9979 5868 9988
rect 5816 9945 5825 9979
rect 5825 9945 5859 9979
rect 5859 9945 5868 9979
rect 5816 9936 5868 9945
rect 6000 9936 6052 9988
rect 6368 9936 6420 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3792 9868 3844 9920
rect 5356 9868 5408 9920
rect 6736 9868 6788 9920
rect 7380 10004 7432 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 9956 10072 10008 10124
rect 10232 10115 10284 10124
rect 10232 10081 10258 10115
rect 10258 10081 10284 10115
rect 10232 10072 10284 10081
rect 10692 10072 10744 10124
rect 10784 10072 10836 10124
rect 7932 10047 7984 10056
rect 7932 10013 7942 10047
rect 7942 10013 7976 10047
rect 7976 10013 7984 10047
rect 7932 10004 7984 10013
rect 8944 10004 8996 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9404 10004 9456 10056
rect 8576 9936 8628 9988
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 9772 9979 9824 9988
rect 9772 9945 9781 9979
rect 9781 9945 9815 9979
rect 9815 9945 9824 9979
rect 9772 9936 9824 9945
rect 9956 9979 10008 9988
rect 9956 9945 9965 9979
rect 9965 9945 9999 9979
rect 9999 9945 10008 9979
rect 9956 9936 10008 9945
rect 11336 10004 11388 10056
rect 13268 10149 13277 10183
rect 13277 10149 13311 10183
rect 13311 10149 13320 10183
rect 13268 10140 13320 10149
rect 12900 10004 12952 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 8484 9868 8536 9920
rect 9312 9868 9364 9920
rect 9496 9868 9548 9920
rect 11428 9936 11480 9988
rect 11704 9979 11756 9988
rect 11704 9945 11713 9979
rect 11713 9945 11747 9979
rect 11747 9945 11756 9979
rect 11704 9936 11756 9945
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 11152 9868 11204 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 1492 9707 1544 9716
rect 1492 9673 1501 9707
rect 1501 9673 1535 9707
rect 1535 9673 1544 9707
rect 1492 9664 1544 9673
rect 3240 9596 3292 9648
rect 5356 9664 5408 9716
rect 5724 9664 5776 9716
rect 4804 9596 4856 9648
rect 2412 9528 2464 9580
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 5356 9528 5408 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 5172 9460 5224 9512
rect 6552 9571 6604 9580
rect 6552 9537 6601 9571
rect 6601 9537 6604 9571
rect 6552 9528 6604 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7840 9596 7892 9648
rect 8760 9664 8812 9716
rect 9496 9664 9548 9716
rect 8852 9596 8904 9648
rect 9956 9664 10008 9716
rect 10876 9707 10928 9716
rect 10876 9673 10885 9707
rect 10885 9673 10919 9707
rect 10919 9673 10928 9707
rect 10876 9664 10928 9673
rect 8208 9528 8260 9580
rect 8576 9528 8628 9580
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 9588 9528 9640 9580
rect 9680 9528 9732 9580
rect 9956 9528 10008 9580
rect 10692 9639 10744 9648
rect 10416 9528 10468 9580
rect 1676 9435 1728 9444
rect 1676 9401 1685 9435
rect 1685 9401 1719 9435
rect 1719 9401 1728 9435
rect 1676 9392 1728 9401
rect 2964 9392 3016 9444
rect 3792 9392 3844 9444
rect 4528 9392 4580 9444
rect 8668 9460 8720 9512
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2412 9324 2464 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 9772 9460 9824 9512
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 9680 9392 9732 9444
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 11428 9664 11480 9716
rect 12808 9664 12860 9716
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 8760 9324 8812 9333
rect 10784 9324 10836 9376
rect 11060 9392 11112 9444
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12716 9528 12768 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 3608 9120 3660 9172
rect 6092 9163 6144 9172
rect 3240 9052 3292 9104
rect 2412 9027 2464 9036
rect 2412 8993 2421 9027
rect 2421 8993 2455 9027
rect 2455 8993 2464 9027
rect 2412 8984 2464 8993
rect 3516 9052 3568 9104
rect 5540 9095 5592 9104
rect 5540 9061 5549 9095
rect 5549 9061 5583 9095
rect 5583 9061 5592 9095
rect 5540 9052 5592 9061
rect 3148 8916 3200 8968
rect 5172 8984 5224 9036
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 7748 9120 7800 9172
rect 8852 9120 8904 9172
rect 3792 8891 3844 8900
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 5264 8916 5316 8968
rect 5356 8916 5408 8968
rect 6644 9052 6696 9104
rect 6920 9052 6972 9104
rect 7288 8984 7340 9036
rect 8024 9052 8076 9104
rect 8760 9052 8812 9104
rect 9036 9052 9088 9104
rect 9680 9120 9732 9172
rect 10140 9120 10192 9172
rect 12072 9120 12124 9172
rect 9404 9052 9456 9104
rect 9588 9095 9640 9104
rect 9588 9061 9597 9095
rect 9597 9061 9631 9095
rect 9631 9061 9640 9095
rect 9588 9052 9640 9061
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 7932 8984 7984 9036
rect 3792 8848 3844 8857
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 7472 8848 7524 8900
rect 6368 8780 6420 8832
rect 6736 8780 6788 8832
rect 7748 8916 7800 8968
rect 10048 9052 10100 9104
rect 10416 9052 10468 9104
rect 10876 9052 10928 9104
rect 11336 9052 11388 9104
rect 10692 8984 10744 9036
rect 7840 8891 7892 8900
rect 7840 8857 7849 8891
rect 7849 8857 7883 8891
rect 7883 8857 7892 8891
rect 7840 8848 7892 8857
rect 8668 8916 8720 8968
rect 8852 8916 8904 8968
rect 9036 8916 9088 8968
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9956 8959 10008 8968
rect 9680 8916 9732 8925
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 11152 8984 11204 9036
rect 10232 8916 10284 8925
rect 9128 8848 9180 8900
rect 9864 8848 9916 8900
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11980 8916 12032 8968
rect 12348 8984 12400 9036
rect 10876 8891 10928 8900
rect 8208 8780 8260 8832
rect 9312 8780 9364 8832
rect 9404 8780 9456 8832
rect 10600 8780 10652 8832
rect 10876 8857 10885 8891
rect 10885 8857 10919 8891
rect 10919 8857 10928 8891
rect 10876 8848 10928 8857
rect 10968 8848 11020 8900
rect 13544 8984 13596 9036
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 12900 8891 12952 8900
rect 12900 8857 12909 8891
rect 12909 8857 12943 8891
rect 12943 8857 12952 8891
rect 12900 8848 12952 8857
rect 13452 8891 13504 8900
rect 11704 8780 11756 8832
rect 12440 8780 12492 8832
rect 13452 8857 13461 8891
rect 13461 8857 13495 8891
rect 13495 8857 13504 8891
rect 13452 8848 13504 8857
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 9864 8576 9916 8628
rect 10600 8576 10652 8628
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 5540 8508 5592 8560
rect 5632 8440 5684 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7104 8440 7156 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 10140 8508 10192 8560
rect 10232 8508 10284 8560
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 9588 8440 9640 8492
rect 9956 8440 10008 8492
rect 10876 8508 10928 8560
rect 11336 8576 11388 8628
rect 12440 8576 12492 8628
rect 12900 8508 12952 8560
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11520 8440 11572 8492
rect 12348 8483 12400 8492
rect 7380 8372 7432 8424
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12900 8372 12952 8424
rect 3332 8347 3384 8356
rect 3332 8313 3341 8347
rect 3341 8313 3375 8347
rect 3375 8313 3384 8347
rect 3332 8304 3384 8313
rect 4804 8347 4856 8356
rect 4804 8313 4813 8347
rect 4813 8313 4847 8347
rect 4847 8313 4856 8347
rect 4804 8304 4856 8313
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 6920 8347 6972 8356
rect 6920 8313 6929 8347
rect 6929 8313 6963 8347
rect 6963 8313 6972 8347
rect 6920 8304 6972 8313
rect 7840 8304 7892 8356
rect 10324 8304 10376 8356
rect 11612 8304 11664 8356
rect 11980 8347 12032 8356
rect 11980 8313 11989 8347
rect 11989 8313 12023 8347
rect 12023 8313 12032 8347
rect 11980 8304 12032 8313
rect 12072 8304 12124 8356
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 3884 8032 3936 8084
rect 8392 8032 8444 8084
rect 9312 8032 9364 8084
rect 11796 8032 11848 8084
rect 4804 7964 4856 8016
rect 3056 7896 3108 7948
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 2872 7828 2924 7880
rect 3516 7896 3568 7948
rect 6092 7896 6144 7948
rect 1952 7760 2004 7812
rect 2964 7803 3016 7812
rect 2964 7769 2973 7803
rect 2973 7769 3007 7803
rect 3007 7769 3016 7803
rect 2964 7760 3016 7769
rect 5540 7828 5592 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 7288 7964 7340 8016
rect 13176 8007 13228 8016
rect 13176 7973 13185 8007
rect 13185 7973 13219 8007
rect 13219 7973 13228 8007
rect 13176 7964 13228 7973
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 2136 7692 2188 7744
rect 4896 7760 4948 7812
rect 6460 7760 6512 7812
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 7472 7828 7524 7880
rect 9128 7896 9180 7948
rect 8392 7760 8444 7812
rect 8576 7760 8628 7812
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 9496 7828 9548 7880
rect 10048 7828 10100 7880
rect 10324 7828 10376 7880
rect 11244 7828 11296 7880
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 12164 7760 12216 7812
rect 7564 7692 7616 7744
rect 8116 7692 8168 7744
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 8760 7692 8812 7744
rect 10416 7692 10468 7744
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 2872 7488 2924 7540
rect 6552 7488 6604 7540
rect 8116 7488 8168 7540
rect 8852 7488 8904 7540
rect 9404 7488 9456 7540
rect 2780 7420 2832 7472
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3884 7352 3936 7404
rect 4804 7420 4856 7472
rect 5540 7420 5592 7472
rect 5632 7463 5684 7472
rect 5632 7429 5641 7463
rect 5641 7429 5675 7463
rect 5675 7429 5684 7463
rect 5632 7420 5684 7429
rect 4896 7395 4948 7404
rect 3516 7216 3568 7268
rect 3700 7216 3752 7268
rect 4620 7284 4672 7336
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 8668 7420 8720 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 7380 7395 7432 7404
rect 6920 7352 6972 7361
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 7840 7395 7892 7404
rect 7840 7361 7863 7395
rect 7863 7361 7892 7395
rect 7840 7352 7892 7361
rect 8208 7352 8260 7404
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 9220 7395 9272 7404
rect 8484 7352 8536 7361
rect 9220 7361 9229 7395
rect 9229 7361 9272 7395
rect 9220 7352 9272 7361
rect 4988 7284 5040 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 7288 7284 7340 7336
rect 7932 7284 7984 7336
rect 8300 7284 8352 7336
rect 8576 7284 8628 7336
rect 8760 7284 8812 7336
rect 9036 7284 9088 7336
rect 9496 7420 9548 7472
rect 10324 7463 10376 7472
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10324 7429 10333 7463
rect 10333 7429 10367 7463
rect 10367 7429 10376 7463
rect 10324 7420 10376 7429
rect 12072 7420 12124 7472
rect 10140 7352 10192 7404
rect 11244 7284 11296 7336
rect 12072 7284 12124 7336
rect 1952 7148 2004 7200
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 4804 7148 4856 7200
rect 9864 7216 9916 7268
rect 12256 7259 12308 7268
rect 12256 7225 12265 7259
rect 12265 7225 12299 7259
rect 12299 7225 12308 7259
rect 12256 7216 12308 7225
rect 6460 7148 6512 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 8576 7148 8628 7200
rect 13176 7148 13228 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 2596 6944 2648 6996
rect 3056 6944 3108 6996
rect 4068 6944 4120 6996
rect 5908 6944 5960 6996
rect 6644 6944 6696 6996
rect 8484 6944 8536 6996
rect 9956 6944 10008 6996
rect 7104 6876 7156 6928
rect 5264 6808 5316 6860
rect 7932 6808 7984 6860
rect 8300 6808 8352 6860
rect 8668 6808 8720 6860
rect 9404 6876 9456 6928
rect 9864 6876 9916 6928
rect 12900 6876 12952 6928
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6740 8812 6792
rect 11888 6808 11940 6860
rect 9680 6740 9732 6792
rect 12348 6740 12400 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 3424 6672 3476 6724
rect 4068 6715 4120 6724
rect 4068 6681 4077 6715
rect 4077 6681 4111 6715
rect 4111 6681 4120 6715
rect 4068 6672 4120 6681
rect 4620 6672 4672 6724
rect 6644 6672 6696 6724
rect 7380 6672 7432 6724
rect 1400 6647 1452 6656
rect 1400 6613 1409 6647
rect 1409 6613 1443 6647
rect 1443 6613 1452 6647
rect 1400 6604 1452 6613
rect 1768 6604 1820 6656
rect 3516 6604 3568 6656
rect 4436 6604 4488 6656
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 8760 6604 8812 6656
rect 9036 6604 9088 6656
rect 11888 6672 11940 6724
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 1952 6400 2004 6452
rect 4068 6443 4120 6452
rect 1400 6264 1452 6316
rect 2136 6264 2188 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 4712 6400 4764 6452
rect 5540 6400 5592 6452
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 4620 6332 4672 6384
rect 5264 6332 5316 6384
rect 6460 6332 6512 6384
rect 2320 6264 2372 6273
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3332 6264 3384 6316
rect 4068 6264 4120 6316
rect 5724 6307 5776 6316
rect 1584 6171 1636 6180
rect 1584 6137 1593 6171
rect 1593 6137 1627 6171
rect 1627 6137 1636 6171
rect 1584 6128 1636 6137
rect 1676 6128 1728 6180
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 3516 6196 3568 6248
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6368 6264 6420 6316
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8576 6400 8628 6452
rect 8852 6400 8904 6452
rect 9036 6375 9088 6384
rect 9036 6341 9045 6375
rect 9045 6341 9079 6375
rect 9079 6341 9088 6375
rect 9036 6332 9088 6341
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8668 6264 8720 6316
rect 8760 6264 8812 6316
rect 9956 6400 10008 6452
rect 11336 6443 11388 6452
rect 10048 6264 10100 6316
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 11888 6332 11940 6384
rect 10692 6264 10744 6273
rect 3608 6171 3660 6180
rect 3608 6137 3617 6171
rect 3617 6137 3651 6171
rect 3651 6137 3660 6171
rect 3608 6128 3660 6137
rect 4528 6196 4580 6248
rect 5356 6196 5408 6248
rect 7564 6196 7616 6248
rect 5172 6128 5224 6180
rect 5908 6128 5960 6180
rect 1400 6060 1452 6069
rect 2964 6060 3016 6112
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5632 6060 5684 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 8484 6128 8536 6180
rect 9312 6196 9364 6248
rect 10324 6196 10376 6248
rect 10784 6196 10836 6248
rect 12072 6264 12124 6316
rect 12992 6332 13044 6384
rect 12348 6264 12400 6316
rect 11612 6171 11664 6180
rect 11612 6137 11621 6171
rect 11621 6137 11655 6171
rect 11655 6137 11664 6171
rect 11612 6128 11664 6137
rect 13268 6196 13320 6248
rect 12072 6128 12124 6180
rect 9036 6060 9088 6112
rect 10324 6060 10376 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 2320 5788 2372 5840
rect 3332 5831 3384 5840
rect 3332 5797 3341 5831
rect 3341 5797 3375 5831
rect 3375 5797 3384 5831
rect 3332 5788 3384 5797
rect 4712 5856 4764 5908
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 3056 5652 3108 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3792 5720 3844 5772
rect 5264 5856 5316 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 10600 5856 10652 5908
rect 11704 5856 11756 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 6920 5788 6972 5840
rect 7932 5720 7984 5772
rect 9404 5788 9456 5840
rect 9680 5788 9732 5840
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 8484 5720 8536 5772
rect 10968 5720 11020 5772
rect 3148 5652 3200 5661
rect 3516 5695 3568 5704
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 4068 5652 4120 5704
rect 6644 5652 6696 5704
rect 7104 5652 7156 5704
rect 8852 5652 8904 5704
rect 9312 5695 9364 5704
rect 3240 5584 3292 5636
rect 3976 5627 4028 5636
rect 3976 5593 3985 5627
rect 3985 5593 4019 5627
rect 4019 5593 4028 5627
rect 3976 5584 4028 5593
rect 4620 5584 4672 5636
rect 5080 5627 5132 5636
rect 5080 5593 5089 5627
rect 5089 5593 5123 5627
rect 5123 5593 5132 5627
rect 5080 5584 5132 5593
rect 5724 5584 5776 5636
rect 8576 5584 8628 5636
rect 8668 5584 8720 5636
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9404 5652 9456 5704
rect 1768 5516 1820 5568
rect 1860 5516 1912 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 7748 5516 7800 5568
rect 9864 5584 9916 5636
rect 10232 5652 10284 5704
rect 10324 5584 10376 5636
rect 11612 5584 11664 5636
rect 9772 5516 9824 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 1768 5312 1820 5364
rect 2596 5312 2648 5364
rect 3608 5312 3660 5364
rect 3056 5244 3108 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 2412 5176 2464 5228
rect 3608 5219 3660 5228
rect 2596 5151 2648 5160
rect 2320 5040 2372 5092
rect 2596 5117 2622 5151
rect 2622 5117 2648 5151
rect 2596 5108 2648 5117
rect 2780 5108 2832 5160
rect 3056 5108 3108 5160
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4068 5219 4120 5228
rect 3700 5108 3752 5160
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 4620 5312 4672 5364
rect 5080 5312 5132 5364
rect 6552 5312 6604 5364
rect 5540 5244 5592 5296
rect 3976 5108 4028 5160
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 8576 5244 8628 5296
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 5172 5176 5224 5185
rect 5356 5108 5408 5160
rect 6092 5176 6144 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 8484 5176 8536 5228
rect 9496 5312 9548 5364
rect 11428 5312 11480 5364
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 9680 5244 9732 5296
rect 9864 5244 9916 5296
rect 11336 5244 11388 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 13176 5244 13228 5296
rect 11612 5176 11664 5228
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 4712 5040 4764 5092
rect 6460 5108 6512 5160
rect 7288 5108 7340 5160
rect 8760 5108 8812 5160
rect 9128 5108 9180 5160
rect 11152 5108 11204 5160
rect 3148 4972 3200 5024
rect 6828 5040 6880 5092
rect 5908 4972 5960 5024
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 12716 4972 12768 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2596 4700 2648 4752
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 3884 4768 3936 4820
rect 4804 4768 4856 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 8484 4811 8536 4820
rect 8484 4777 8493 4811
rect 8493 4777 8527 4811
rect 8527 4777 8536 4811
rect 8484 4768 8536 4777
rect 8760 4768 8812 4820
rect 9312 4768 9364 4820
rect 10140 4768 10192 4820
rect 10232 4768 10284 4820
rect 2964 4743 3016 4752
rect 2964 4709 2969 4743
rect 2969 4709 3003 4743
rect 3003 4709 3016 4743
rect 1676 4564 1728 4616
rect 2136 4564 2188 4616
rect 2228 4564 2280 4616
rect 1584 4496 1636 4548
rect 2964 4700 3016 4709
rect 3792 4675 3844 4684
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 6644 4700 6696 4752
rect 7012 4700 7064 4752
rect 2872 4496 2924 4548
rect 1400 4471 1452 4480
rect 1400 4437 1409 4471
rect 1409 4437 1443 4471
rect 1443 4437 1452 4471
rect 1400 4428 1452 4437
rect 5816 4564 5868 4616
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 7748 4675 7800 4684
rect 6828 4632 6880 4641
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 6460 4564 6512 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 8668 4564 8720 4616
rect 9680 4700 9732 4752
rect 13176 4743 13228 4752
rect 13176 4709 13185 4743
rect 13185 4709 13219 4743
rect 13219 4709 13228 4743
rect 13176 4700 13228 4709
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 11888 4632 11940 4684
rect 9956 4564 10008 4616
rect 10232 4607 10284 4616
rect 4344 4496 4396 4548
rect 4712 4496 4764 4548
rect 3148 4428 3200 4480
rect 3608 4428 3660 4480
rect 5632 4496 5684 4548
rect 6000 4496 6052 4548
rect 7932 4496 7984 4548
rect 8760 4539 8812 4548
rect 8760 4505 8769 4539
rect 8769 4505 8803 4539
rect 8803 4505 8812 4539
rect 8760 4496 8812 4505
rect 9864 4539 9916 4548
rect 9864 4505 9873 4539
rect 9873 4505 9907 4539
rect 9907 4505 9916 4539
rect 9864 4496 9916 4505
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 12072 4564 12124 4616
rect 12624 4564 12676 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 10140 4496 10192 4548
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 9220 4428 9272 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 1768 4224 1820 4276
rect 4344 4224 4396 4276
rect 4068 4199 4120 4208
rect 4068 4165 4077 4199
rect 4077 4165 4111 4199
rect 4111 4165 4120 4199
rect 4068 4156 4120 4165
rect 5540 4224 5592 4276
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 6920 4224 6972 4276
rect 8576 4267 8628 4276
rect 8576 4233 8585 4267
rect 8585 4233 8619 4267
rect 8619 4233 8628 4267
rect 8576 4224 8628 4233
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 11612 4267 11664 4276
rect 11612 4233 11621 4267
rect 11621 4233 11655 4267
rect 11655 4233 11664 4267
rect 11612 4224 11664 4233
rect 11888 4224 11940 4276
rect 1676 4088 1728 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2872 4088 2924 4140
rect 3240 4088 3292 4140
rect 5264 4088 5316 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6368 4088 6420 4140
rect 6644 4088 6696 4140
rect 6920 4088 6972 4140
rect 8484 4131 8536 4140
rect 1952 4020 2004 4072
rect 2412 4020 2464 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 1492 3952 1544 4004
rect 4896 3952 4948 4004
rect 6460 4020 6512 4072
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 8392 4020 8444 4072
rect 8668 4088 8720 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 5908 3952 5960 4004
rect 8760 4020 8812 4072
rect 9680 4156 9732 4208
rect 11428 4088 11480 4140
rect 11888 4131 11940 4140
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 12808 4224 12860 4276
rect 12624 4156 12676 4208
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 13544 4088 13596 4140
rect 1860 3884 1912 3936
rect 2596 3884 2648 3936
rect 8116 3884 8168 3936
rect 8944 3952 8996 4004
rect 9404 3995 9456 4004
rect 9404 3961 9413 3995
rect 9413 3961 9447 3995
rect 9447 3961 9456 3995
rect 9404 3952 9456 3961
rect 9956 3884 10008 3936
rect 10140 3884 10192 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 2964 3680 3016 3732
rect 3976 3680 4028 3732
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 3332 3655 3384 3664
rect 1584 3544 1636 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 1768 3476 1820 3528
rect 2596 3587 2648 3596
rect 2320 3476 2372 3528
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 8668 3680 8720 3732
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 9772 3680 9824 3732
rect 10324 3723 10376 3732
rect 5264 3612 5316 3664
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5540 3519 5592 3528
rect 5264 3476 5316 3485
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7196 3612 7248 3664
rect 8944 3612 8996 3664
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 11888 3680 11940 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 10048 3655 10100 3664
rect 10048 3621 10057 3655
rect 10057 3621 10091 3655
rect 10091 3621 10100 3655
rect 10048 3612 10100 3621
rect 6552 3544 6604 3596
rect 6920 3544 6972 3596
rect 8392 3544 8444 3596
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 11428 3544 11480 3596
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 9864 3519 9916 3528
rect 6644 3476 6696 3485
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 12808 3476 12860 3528
rect 6828 3408 6880 3460
rect 7932 3408 7984 3460
rect 10692 3451 10744 3460
rect 6920 3340 6972 3392
rect 7472 3340 7524 3392
rect 9588 3340 9640 3392
rect 10692 3417 10701 3451
rect 10701 3417 10735 3451
rect 10735 3417 10744 3451
rect 10692 3408 10744 3417
rect 10600 3340 10652 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 2872 3111 2924 3120
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2872 3077 2881 3111
rect 2881 3077 2915 3111
rect 2915 3077 2924 3111
rect 2872 3068 2924 3077
rect 3240 3111 3292 3120
rect 3240 3077 3249 3111
rect 3249 3077 3283 3111
rect 3283 3077 3292 3111
rect 3240 3068 3292 3077
rect 4620 3136 4672 3188
rect 5264 3136 5316 3188
rect 6092 3179 6144 3188
rect 2872 2932 2924 2984
rect 4252 3000 4304 3052
rect 4620 3000 4672 3052
rect 4344 2932 4396 2984
rect 4712 2932 4764 2984
rect 4988 3068 5040 3120
rect 6092 3145 6101 3179
rect 6101 3145 6135 3179
rect 6135 3145 6144 3179
rect 6092 3136 6144 3145
rect 6644 3136 6696 3188
rect 7472 3179 7524 3188
rect 5264 3000 5316 3052
rect 7104 3068 7156 3120
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 8576 3136 8628 3188
rect 8760 3136 8812 3188
rect 9404 3136 9456 3188
rect 10600 3179 10652 3188
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 7196 3043 7248 3052
rect 6920 3000 6972 3009
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7472 3000 7524 3052
rect 5448 2932 5500 2984
rect 2596 2796 2648 2848
rect 7196 2864 7248 2916
rect 7748 2932 7800 2984
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 9680 3000 9732 3052
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 10692 3136 10744 3188
rect 11888 3136 11940 3188
rect 10968 3000 11020 3052
rect 11428 3000 11480 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 8208 2932 8260 2984
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 12716 2975 12768 2984
rect 6000 2796 6052 2848
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 11704 2864 11756 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 2504 2592 2556 2644
rect 4712 2592 4764 2644
rect 4068 2524 4120 2576
rect 5908 2592 5960 2644
rect 6184 2592 6236 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 8576 2592 8628 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 10692 2592 10744 2644
rect 3240 2499 3292 2508
rect 3240 2465 3249 2499
rect 3249 2465 3283 2499
rect 3283 2465 3292 2499
rect 3240 2456 3292 2465
rect 8300 2456 8352 2508
rect 2044 2252 2096 2304
rect 4068 2388 4120 2440
rect 5264 2388 5316 2440
rect 5448 2388 5500 2440
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7564 2388 7616 2440
rect 7748 2388 7800 2440
rect 4620 2363 4672 2372
rect 4620 2329 4629 2363
rect 4629 2329 4663 2363
rect 4663 2329 4672 2363
rect 4620 2320 4672 2329
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6092 2320 6144 2372
rect 7196 2320 7248 2372
rect 7104 2252 7156 2304
rect 7288 2295 7340 2304
rect 7288 2261 7297 2295
rect 7297 2261 7331 2295
rect 7331 2261 7340 2295
rect 7288 2252 7340 2261
rect 8024 2252 8076 2304
rect 9496 2524 9548 2576
rect 8944 2456 8996 2508
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 9680 2456 9732 2508
rect 9404 2388 9456 2440
rect 12624 2524 12676 2576
rect 13176 2499 13228 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 12716 2388 12768 2440
rect 9312 2252 9364 2304
rect 11704 2320 11756 2372
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 1952 2048 2004 2100
rect 3240 2048 3292 2100
rect 3608 2091 3660 2100
rect 3608 2057 3617 2091
rect 3617 2057 3651 2091
rect 3651 2057 3660 2091
rect 3608 2048 3660 2057
rect 5356 2048 5408 2100
rect 6092 2091 6144 2100
rect 6092 2057 6101 2091
rect 6101 2057 6135 2091
rect 6135 2057 6144 2091
rect 6092 2048 6144 2057
rect 6460 2091 6512 2100
rect 6460 2057 6469 2091
rect 6469 2057 6503 2091
rect 6503 2057 6512 2091
rect 6460 2048 6512 2057
rect 9404 2048 9456 2100
rect 10876 2048 10928 2100
rect 13176 2048 13228 2100
rect 4620 1980 4672 2032
rect 3332 1955 3384 1964
rect 3332 1921 3341 1955
rect 3341 1921 3375 1955
rect 3375 1921 3384 1955
rect 3792 1955 3844 1964
rect 3332 1912 3384 1921
rect 3792 1921 3801 1955
rect 3801 1921 3835 1955
rect 3835 1921 3844 1955
rect 3792 1912 3844 1921
rect 7840 1980 7892 2032
rect 8024 1980 8076 2032
rect 10416 1980 10468 2032
rect 6000 1955 6052 1964
rect 6000 1921 6009 1955
rect 6009 1921 6043 1955
rect 6043 1921 6052 1955
rect 6000 1912 6052 1921
rect 6644 1912 6696 1964
rect 2780 1844 2832 1896
rect 4068 1887 4120 1896
rect 4068 1853 4077 1887
rect 4077 1853 4111 1887
rect 4111 1853 4120 1887
rect 4068 1844 4120 1853
rect 8484 1887 8536 1896
rect 8484 1853 8493 1887
rect 8493 1853 8527 1887
rect 8527 1853 8536 1887
rect 8484 1844 8536 1853
rect 8760 1887 8812 1896
rect 8760 1853 8769 1887
rect 8769 1853 8803 1887
rect 8803 1853 8812 1887
rect 8760 1844 8812 1853
rect 10692 1955 10744 1964
rect 10692 1921 10701 1955
rect 10701 1921 10735 1955
rect 10735 1921 10744 1955
rect 10692 1912 10744 1921
rect 10968 1955 11020 1964
rect 10968 1921 10977 1955
rect 10977 1921 11011 1955
rect 11011 1921 11020 1955
rect 10968 1912 11020 1921
rect 12072 1980 12124 2032
rect 6552 1708 6604 1760
rect 7104 1708 7156 1760
rect 9496 1708 9548 1760
rect 10968 1776 11020 1828
rect 10692 1708 10744 1760
rect 11796 1887 11848 1896
rect 11796 1853 11805 1887
rect 11805 1853 11839 1887
rect 11839 1853 11848 1887
rect 11796 1844 11848 1853
rect 11612 1708 11664 1760
rect 11980 1708 12032 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 2228 1504 2280 1556
rect 4068 1504 4120 1556
rect 5816 1504 5868 1556
rect 3240 1436 3292 1488
rect 2044 1411 2096 1420
rect 2044 1377 2053 1411
rect 2053 1377 2087 1411
rect 2087 1377 2096 1411
rect 2044 1368 2096 1377
rect 2596 1368 2648 1420
rect 1492 1343 1544 1352
rect 1492 1309 1501 1343
rect 1501 1309 1535 1343
rect 1535 1309 1544 1343
rect 1492 1300 1544 1309
rect 3608 1368 3660 1420
rect 3976 1343 4028 1352
rect 3976 1309 3985 1343
rect 3985 1309 4019 1343
rect 4019 1309 4028 1343
rect 3976 1300 4028 1309
rect 5908 1436 5960 1488
rect 4436 1343 4488 1352
rect 4436 1309 4445 1343
rect 4445 1309 4479 1343
rect 4479 1309 4488 1343
rect 4436 1300 4488 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 5448 1300 5500 1352
rect 3332 1164 3384 1216
rect 5356 1232 5408 1284
rect 6552 1368 6604 1420
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 7564 1436 7616 1488
rect 7012 1368 7064 1420
rect 7288 1368 7340 1420
rect 7472 1368 7524 1420
rect 7840 1368 7892 1420
rect 9496 1504 9548 1556
rect 11152 1504 11204 1556
rect 11796 1504 11848 1556
rect 11980 1504 12032 1556
rect 8760 1436 8812 1488
rect 8484 1368 8536 1420
rect 10416 1368 10468 1420
rect 10968 1368 11020 1420
rect 7104 1343 7156 1352
rect 7104 1309 7113 1343
rect 7113 1309 7147 1343
rect 7147 1309 7156 1343
rect 7104 1300 7156 1309
rect 8116 1343 8168 1352
rect 8116 1309 8125 1343
rect 8125 1309 8159 1343
rect 8159 1309 8168 1343
rect 8116 1300 8168 1309
rect 8208 1300 8260 1352
rect 6460 1207 6512 1216
rect 6460 1173 6469 1207
rect 6469 1173 6503 1207
rect 6503 1173 6512 1207
rect 8024 1232 8076 1284
rect 8944 1300 8996 1352
rect 9404 1300 9456 1352
rect 10876 1300 10928 1352
rect 11612 1343 11664 1352
rect 11612 1309 11621 1343
rect 11621 1309 11655 1343
rect 11655 1309 11664 1343
rect 11612 1300 11664 1309
rect 12072 1300 12124 1352
rect 9496 1232 9548 1284
rect 11152 1232 11204 1284
rect 6460 1164 6512 1173
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 3700 960 3752 1012
rect 6460 960 6512 1012
rect 8024 960 8076 1012
rect 4436 892 4488 944
rect 6000 892 6052 944
rect 8116 892 8168 944
<< metal2 >>
rect 570 14200 626 15000
rect 1674 14200 1730 15000
rect 2870 14200 2926 15000
rect 3698 14512 3754 14521
rect 3698 14447 3754 14456
rect 584 13530 612 14200
rect 1688 13734 1716 14200
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 572 13524 624 13530
rect 572 13466 624 13472
rect 2056 13326 2084 13738
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1412 12986 1440 13194
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12617 1440 12718
rect 1398 12608 1454 12617
rect 1398 12543 1454 12552
rect 1412 9178 1440 12543
rect 1596 12170 1624 12786
rect 2056 12306 2084 13262
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2148 12238 2176 13194
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 2240 11830 2268 13126
rect 2332 12850 2360 13262
rect 2884 13190 2912 14200
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2792 12986 2820 13126
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2332 11830 2360 12106
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1688 11218 1716 11630
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 2332 11150 2360 11766
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2516 10742 2544 11698
rect 2700 11626 2728 12106
rect 2792 12102 2820 12922
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12374 2912 12786
rect 3252 12714 3280 13194
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2700 11286 2728 11562
rect 2792 11558 2820 12038
rect 2884 11762 2912 12310
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11898 3004 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 3424 11688 3476 11694
rect 3054 11656 3110 11665
rect 3424 11630 3476 11636
rect 3054 11591 3110 11600
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2792 10996 2820 11494
rect 3068 11150 3096 11591
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2964 11008 3016 11014
rect 2792 10968 2964 10996
rect 2964 10950 3016 10956
rect 2504 10736 2556 10742
rect 1582 10704 1638 10713
rect 2504 10678 2556 10684
rect 1504 10648 1582 10656
rect 1504 10628 1584 10648
rect 1504 9722 1532 10628
rect 1636 10639 1638 10648
rect 1768 10668 1820 10674
rect 1584 10610 1636 10616
rect 1768 10610 1820 10616
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1596 10062 1624 10474
rect 1780 10266 1808 10610
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1492 9716 1544 9722
rect 1780 9674 1808 10202
rect 1872 10130 1900 10610
rect 2516 10198 2544 10678
rect 2976 10470 3004 10950
rect 3068 10810 3096 11086
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3252 10674 3280 11086
rect 3436 10674 3464 11630
rect 3528 10810 3556 12242
rect 3620 12102 3648 12310
rect 3712 12238 3740 14447
rect 3974 14362 4030 15000
rect 3974 14334 4108 14362
rect 3974 14200 4030 14334
rect 3790 13560 3846 13569
rect 3790 13495 3846 13504
rect 3804 13326 3832 13495
rect 4080 13462 4108 14334
rect 5170 14200 5226 15000
rect 6274 14200 6330 15000
rect 7470 14362 7526 15000
rect 8574 14362 8630 15000
rect 7470 14334 7696 14362
rect 7470 14200 7526 14334
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11830 3648 12038
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3712 10742 3740 12174
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1492 9658 1544 9664
rect 1688 9646 1808 9674
rect 1688 9450 1716 9646
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 2424 9382 2452 9522
rect 2976 9450 3004 10406
rect 3344 10266 3372 10542
rect 3804 10266 3832 13262
rect 3988 12782 4016 13262
rect 4080 12850 4108 13398
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12776 4028 12782
rect 4172 12730 4200 13194
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12986 4476 13126
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4632 12850 4660 13262
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 3976 12718 4028 12724
rect 3988 12170 4016 12718
rect 4080 12702 4200 12730
rect 4080 12434 4108 12702
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4080 12406 4200 12434
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 4172 11762 4200 12406
rect 4632 12374 4660 12786
rect 4724 12442 4752 13330
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5092 12918 5120 13194
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4356 12073 4384 12174
rect 4342 12064 4398 12073
rect 4342 11999 4398 12008
rect 4816 11830 4844 12650
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4172 11642 4200 11698
rect 4080 11614 4200 11642
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4080 11150 4108 11614
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10742 4292 11086
rect 4632 10810 4660 11630
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4724 11150 4752 11562
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11286 4844 11494
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3160 9586 3188 9998
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9654 3280 9862
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1504 8090 1532 8434
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 2148 7886 2176 9318
rect 2424 9042 2452 9318
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 3160 8974 3188 9522
rect 3252 9110 3280 9590
rect 3344 9178 3372 9687
rect 3620 9586 3648 9998
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3620 9178 3648 9522
rect 3804 9450 3832 9862
rect 4540 9450 4568 9930
rect 4816 9654 4844 11222
rect 4908 11082 4936 12106
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 5000 10198 5028 12582
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 10742 5120 11494
rect 5184 11150 5212 14200
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 5276 12374 5304 13262
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5354 12880 5410 12889
rect 5354 12815 5410 12824
rect 5540 12844 5592 12850
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 5092 9994 5120 10406
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5368 9926 5396 12815
rect 5540 12786 5592 12792
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5552 11762 5580 12786
rect 5644 12170 5672 12786
rect 5736 12238 5764 13194
rect 6104 12850 6132 13262
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11830 5672 12106
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10266 5488 11086
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10266 5580 10950
rect 5736 10470 5764 11698
rect 5920 10674 5948 11834
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6012 11014 6040 11698
rect 6196 11218 6224 11698
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5552 9994 5580 10202
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9722 5396 9862
rect 5736 9722 5764 10406
rect 5816 9988 5868 9994
rect 5920 9976 5948 10610
rect 6196 10538 6224 11154
rect 6288 10810 6316 14200
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6656 12850 6684 13398
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6748 12442 6776 13262
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12850 6868 13126
rect 6932 12889 6960 13194
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6918 12880 6974 12889
rect 6828 12844 6880 12850
rect 7024 12850 7052 12922
rect 6918 12815 6974 12824
rect 7012 12844 7064 12850
rect 6828 12786 6880 12792
rect 7012 12786 7064 12792
rect 6840 12646 6868 12786
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6840 12306 6868 12582
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6550 12200 6606 12209
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6380 11898 6408 12106
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 11558 6500 12174
rect 6736 12164 6788 12170
rect 6550 12135 6552 12144
rect 6604 12135 6606 12144
rect 6552 12106 6604 12112
rect 6656 12124 6736 12152
rect 6552 11824 6604 11830
rect 6550 11792 6552 11801
rect 6604 11792 6606 11801
rect 6550 11727 6606 11736
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6460 11552 6512 11558
rect 6564 11529 6592 11562
rect 6460 11494 6512 11500
rect 6550 11520 6606 11529
rect 6472 11150 6500 11494
rect 6550 11455 6606 11464
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6552 11144 6604 11150
rect 6656 11132 6684 12124
rect 6736 12106 6788 12112
rect 6932 11898 6960 12650
rect 7116 12238 7144 13670
rect 7392 13530 7420 13670
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7194 12472 7250 12481
rect 7194 12407 7196 12416
rect 7248 12407 7250 12416
rect 7196 12378 7248 12384
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7300 12102 7328 12922
rect 7392 12850 7420 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7286 11928 7342 11937
rect 6920 11892 6972 11898
rect 7286 11863 7342 11872
rect 6920 11834 6972 11840
rect 7300 11830 7328 11863
rect 7288 11824 7340 11830
rect 6734 11792 6790 11801
rect 7194 11792 7250 11801
rect 6734 11727 6790 11736
rect 7104 11756 7156 11762
rect 6604 11104 6684 11132
rect 6552 11086 6604 11092
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 10418 6224 10474
rect 6012 10390 6224 10418
rect 6012 9994 6040 10390
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5868 9948 5948 9976
rect 6000 9988 6052 9994
rect 5816 9930 5868 9936
rect 6000 9930 6052 9936
rect 5356 9716 5408 9722
rect 5276 9664 5356 9674
rect 5276 9658 5408 9664
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 5276 9646 5396 9658
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3528 8498 3556 9046
rect 3804 8906 3832 9386
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5184 9042 5212 9454
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5276 8974 5304 9646
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5368 8974 5396 9522
rect 5552 9110 5580 9522
rect 6104 9178 6132 10066
rect 6288 10062 6316 10746
rect 6564 10538 6592 11086
rect 6748 11064 6776 11727
rect 7288 11766 7340 11772
rect 7194 11727 7250 11736
rect 7104 11698 7156 11704
rect 7116 11665 7144 11698
rect 7102 11656 7158 11665
rect 7208 11626 7236 11727
rect 7102 11591 7158 11600
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 6826 11384 6882 11393
rect 6826 11319 6828 11328
rect 6880 11319 6882 11328
rect 7104 11348 7156 11354
rect 6828 11290 6880 11296
rect 7104 11290 7156 11296
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6656 11036 6776 11064
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6380 9994 6408 10406
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6550 9616 6606 9625
rect 6550 9551 6552 9560
rect 6604 9551 6606 9560
rect 6552 9522 6604 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 2226 7984 2282 7993
rect 2226 7919 2282 7928
rect 3056 7948 3108 7954
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7410 1992 7754
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7410 2176 7686
rect 2240 7546 2268 7919
rect 3056 7890 3108 7896
rect 2872 7880 2924 7886
rect 3068 7834 3096 7890
rect 2872 7822 2924 7828
rect 2884 7546 2912 7822
rect 2976 7818 3096 7834
rect 2964 7812 3096 7818
rect 3016 7806 3096 7812
rect 2964 7754 3016 7760
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1412 6322 1440 6598
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 6118 1440 6258
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1400 6112 1452 6118
rect 1398 6080 1400 6089
rect 1452 6080 1454 6089
rect 1398 6015 1454 6024
rect 1596 4554 1624 6122
rect 1688 5914 1716 6122
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1780 5574 1808 6598
rect 1964 6458 1992 7142
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1964 5710 1992 6394
rect 2148 6322 2176 7346
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 7002 2636 7142
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5846 2360 6258
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1780 5370 1808 5510
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1780 5234 1808 5306
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1780 5137 1808 5170
rect 1766 5128 1822 5137
rect 1766 5063 1822 5072
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1584 4548 1636 4554
rect 1584 4490 1636 4496
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 4185 1440 4422
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 1412 3534 1440 4111
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1504 3233 1532 3946
rect 1596 3602 1624 4490
rect 1688 4146 1716 4558
rect 1780 4282 1808 5063
rect 1872 4690 1900 5510
rect 2608 5370 2636 5646
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3670 1716 4082
rect 1872 3942 1900 4626
rect 2148 4622 2176 4966
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2148 4146 2176 4558
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1964 3754 1992 4014
rect 1780 3726 1992 3754
rect 2240 3738 2268 4558
rect 2332 4146 2360 5034
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2424 4078 2452 5170
rect 2792 5166 2820 7414
rect 3068 7342 3096 7806
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 7002 3096 7278
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3344 6474 3372 8298
rect 3528 7954 3556 8434
rect 3804 7970 3832 8842
rect 3884 8832 3936 8838
rect 3882 8800 3884 8809
rect 3936 8800 3938 8809
rect 3882 8735 3938 8744
rect 3896 8090 3924 8735
rect 5368 8634 5396 8910
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 4816 8022 4844 8298
rect 4804 8016 4856 8022
rect 3516 7948 3568 7954
rect 3804 7942 3924 7970
rect 4804 7958 4856 7964
rect 3516 7890 3568 7896
rect 3896 7750 3924 7942
rect 5552 7886 5580 8502
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5644 7886 5672 8434
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7410 3924 7686
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4816 7290 4844 7414
rect 4908 7410 4936 7754
rect 5552 7478 5580 7822
rect 5644 7478 5672 7822
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4988 7336 5040 7342
rect 3436 6730 3464 7278
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3528 6662 3556 7210
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3344 6446 3464 6474
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2608 4758 2636 5102
rect 2976 4758 3004 6054
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3068 5302 3096 5646
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4842 3096 5102
rect 3160 5030 3188 5646
rect 3252 5642 3280 6258
rect 3344 5846 3372 6258
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3068 4814 3188 4842
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2884 4146 2912 4490
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2228 3732 2280 3738
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1780 3534 1808 3726
rect 2228 3674 2280 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1504 3058 1532 3159
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1504 1358 1532 2994
rect 1780 2281 1808 2994
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1766 2272 1822 2281
rect 1766 2207 1822 2216
rect 1964 2106 1992 2382
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1952 2100 2004 2106
rect 1952 2042 2004 2048
rect 2056 1426 2084 2246
rect 2240 1562 2268 3674
rect 2608 3602 2636 3878
rect 2976 3738 3004 4694
rect 3160 4486 3188 4814
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2332 3194 2360 3470
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 3252 3126 3280 4082
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3344 3670 3372 4014
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2516 2650 2544 2994
rect 2884 2990 2912 3062
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 2608 1426 2636 2790
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3252 2106 3280 2450
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2044 1420 2096 1426
rect 2044 1362 2096 1368
rect 2596 1420 2648 1426
rect 2596 1362 2648 1368
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 2792 513 2820 1838
rect 3252 1494 3280 2042
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3240 1488 3292 1494
rect 3240 1430 3292 1436
rect 3344 1222 3372 1906
rect 3436 1329 3464 6446
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3528 5710 3556 6190
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3620 5370 3648 6122
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3620 5234 3648 5306
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 5166 3740 7210
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4066 7032 4122 7041
rect 4214 7035 4522 7044
rect 4066 6967 4068 6976
rect 4120 6967 4122 6976
rect 4068 6938 4120 6944
rect 4632 6730 4660 7278
rect 4816 7262 4936 7290
rect 4988 7278 5040 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4080 6458 4108 6666
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 4690 3832 5714
rect 4080 5710 4108 6258
rect 4448 6236 4476 6598
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4528 6248 4580 6254
rect 4448 6208 4528 6236
rect 4528 6190 4580 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4632 5642 4660 6326
rect 4724 5914 4752 6394
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 3988 5166 4016 5578
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5234 4108 5510
rect 4632 5370 4660 5578
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 2106 3648 4422
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3620 1426 3648 2042
rect 3804 1970 3832 4626
rect 3896 2774 3924 4762
rect 3988 3738 4016 5102
rect 4080 4214 4108 5170
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4724 4554 4752 5034
rect 4816 4826 4844 7142
rect 4908 6118 4936 7262
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4356 4282 4384 4490
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4908 4010 4936 6054
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4264 3058 4292 3470
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4356 2990 4384 3470
rect 4632 3194 4660 3470
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 5000 3126 5028 7278
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5276 6390 5304 6802
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6458 5580 6598
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 5092 5370 5120 5578
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5184 5234 5212 6122
rect 5276 5914 5304 6326
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5368 5166 5396 6190
rect 5552 5302 5580 6394
rect 5736 6322 5764 8298
rect 5828 7410 5856 8434
rect 6380 8362 6408 8774
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7954 6132 8230
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 7313 5856 7346
rect 5814 7304 5870 7313
rect 5814 7239 5870 7248
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5920 6186 5948 6938
rect 6380 6322 6408 8298
rect 6472 7818 6500 9318
rect 6656 9110 6684 11036
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10441 6776 10542
rect 6932 10470 6960 10950
rect 7024 10742 7052 11222
rect 7116 11218 7144 11290
rect 7300 11218 7328 11494
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7288 11076 7340 11082
rect 7392 11064 7420 12650
rect 7484 12646 7512 13670
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7576 12918 7604 13194
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 12073 7604 12106
rect 7562 12064 7618 12073
rect 7340 11036 7420 11064
rect 7288 11018 7340 11024
rect 7392 10985 7420 11036
rect 7484 12022 7562 12050
rect 7378 10976 7434 10985
rect 7378 10911 7434 10920
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 6920 10464 6972 10470
rect 6734 10432 6790 10441
rect 6920 10406 6972 10412
rect 6734 10367 6790 10376
rect 6932 10062 6960 10406
rect 7116 10198 7144 10678
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7392 10305 7420 10474
rect 7378 10296 7434 10305
rect 7288 10260 7340 10266
rect 7378 10231 7380 10240
rect 7288 10202 7340 10208
rect 7432 10231 7434 10240
rect 7380 10202 7432 10208
rect 7104 10192 7156 10198
rect 7300 10169 7328 10202
rect 7104 10134 7156 10140
rect 7286 10160 7342 10169
rect 7286 10095 7342 10104
rect 7392 10062 7420 10202
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9586 6776 9862
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6748 8838 6776 9522
rect 6932 9110 6960 9998
rect 7378 9616 7434 9625
rect 7288 9580 7340 9586
rect 7378 9551 7434 9560
rect 7288 9522 7340 9528
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7300 9042 7328 9522
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6840 7954 6868 8434
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6390 6500 7142
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 6380 6118 6408 6258
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5644 4554 5672 6054
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3670 5304 4082
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5276 3534 5304 3606
rect 5552 3534 5580 4218
rect 5644 4146 5672 4490
rect 5736 4282 5764 5578
rect 6472 5250 6500 6326
rect 6564 5914 6592 7482
rect 6932 7410 6960 8298
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 7002 6684 7142
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6656 6458 6684 6666
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6564 5370 6592 5850
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6380 5222 6500 5250
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5816 4616 5868 4622
rect 5920 4604 5948 4966
rect 5868 4576 5948 4604
rect 5816 4558 5868 4564
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5920 4010 5948 4576
rect 6104 4570 6132 5170
rect 6012 4554 6132 4570
rect 6000 4548 6132 4554
rect 6052 4542 6132 4548
rect 6000 4490 6052 4496
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5276 3194 5304 3470
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 3896 2746 4016 2774
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3988 1358 4016 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4080 2446 4108 2518
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4632 2378 4660 2994
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2650 4752 2926
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5276 2446 5304 2994
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 2446 5488 2926
rect 5920 2836 5948 3946
rect 6104 3194 6132 4542
rect 6380 4146 6408 5222
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4622 6500 5102
rect 6564 4622 6592 5306
rect 6656 4758 6684 5646
rect 6932 5234 6960 5782
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6840 4690 6868 5034
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6472 4282 6500 4558
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6472 3534 6500 4014
rect 6564 3602 6592 4558
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6656 3534 6684 4082
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6000 2848 6052 2854
rect 5920 2808 6000 2836
rect 5920 2650 5948 2808
rect 6000 2790 6052 2796
rect 6104 2774 6132 3130
rect 6104 2746 6224 2774
rect 6196 2650 6224 2746
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 5264 2440 5316 2446
rect 5448 2440 5500 2446
rect 5316 2400 5396 2428
rect 5264 2382 5316 2388
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 5368 2106 5396 2400
rect 5448 2382 5500 2388
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4080 1562 4108 1838
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4068 1556 4120 1562
rect 4068 1498 4120 1504
rect 4632 1358 4660 1974
rect 3976 1352 4028 1358
rect 3422 1320 3478 1329
rect 3976 1294 4028 1300
rect 4436 1352 4488 1358
rect 4436 1294 4488 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 3422 1255 3478 1264
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3700 1012 3752 1018
rect 3700 954 3752 960
rect 3712 800 3740 954
rect 4448 950 4476 1294
rect 5368 1290 5396 2042
rect 5460 1358 5488 2382
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5828 1562 5856 2314
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 5920 1494 5948 2586
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6104 2106 6132 2314
rect 6472 2106 6500 3470
rect 6656 3194 6684 3470
rect 6840 3466 6868 4626
rect 6932 4282 6960 5170
rect 7024 4758 7052 8910
rect 7392 8634 7420 9551
rect 7484 8906 7512 12022
rect 7562 11999 7618 12008
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 10674 7604 11494
rect 7668 10826 7696 14334
rect 8574 14334 8708 14362
rect 8574 14200 8630 14334
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12850 8156 13262
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8574 12880 8630 12889
rect 8116 12844 8168 12850
rect 8574 12815 8630 12824
rect 8116 12786 8168 12792
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8496 12442 8524 12650
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8588 12374 8616 12815
rect 8576 12368 8628 12374
rect 8390 12336 8446 12345
rect 8576 12310 8628 12316
rect 8390 12271 8446 12280
rect 8404 12238 8432 12271
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8588 12170 8616 12310
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11830 7788 12038
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7852 11286 7880 12106
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8022 11928 8078 11937
rect 8214 11931 8522 11940
rect 8022 11863 8078 11872
rect 8036 11762 8064 11863
rect 8024 11756 8076 11762
rect 8484 11756 8536 11762
rect 8076 11716 8484 11744
rect 8024 11698 8076 11704
rect 8484 11698 8536 11704
rect 8390 11656 8446 11665
rect 8116 11620 8168 11626
rect 8446 11600 8616 11608
rect 8390 11591 8392 11600
rect 8116 11562 8168 11568
rect 8444 11580 8616 11600
rect 8392 11562 8444 11568
rect 8024 11348 8076 11354
rect 8128 11336 8156 11562
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8076 11308 8156 11336
rect 8024 11290 8076 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 8220 11218 8248 11494
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7930 11112 7986 11121
rect 8128 11098 8156 11154
rect 7930 11047 7986 11056
rect 8036 11070 8156 11098
rect 7944 11014 7972 11047
rect 7932 11008 7984 11014
rect 7838 10976 7894 10985
rect 7932 10950 7984 10956
rect 7838 10911 7894 10920
rect 7668 10798 7788 10826
rect 7564 10668 7616 10674
rect 7616 10628 7696 10656
rect 7564 10610 7616 10616
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 10062 7604 10474
rect 7668 10266 7696 10628
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7760 9625 7788 10798
rect 7852 9654 7880 10911
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7944 10062 7972 10678
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9648 7892 9654
rect 7746 9616 7802 9625
rect 7840 9590 7892 9596
rect 7746 9551 7802 9560
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8974 7788 9114
rect 7944 9042 7972 9998
rect 8036 9110 8064 11070
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10724 8156 10950
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8588 10792 8616 11580
rect 8312 10764 8616 10792
rect 8208 10736 8260 10742
rect 8128 10696 8208 10724
rect 8128 10305 8156 10696
rect 8208 10678 8260 10684
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 8312 9908 8340 10764
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8496 9926 8524 10202
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8128 9880 8340 9908
rect 8484 9920 8536 9926
rect 8128 9674 8156 9880
rect 8484 9862 8536 9868
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8128 9646 8340 9674
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7116 7342 7144 8434
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7300 7342 7328 7958
rect 7392 7834 7420 8366
rect 7472 7880 7524 7886
rect 7392 7828 7472 7834
rect 7392 7822 7524 7828
rect 7392 7806 7512 7822
rect 7392 7410 7420 7806
rect 7576 7750 7604 8434
rect 7852 8362 7880 8842
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7449 7604 7686
rect 7562 7440 7618 7449
rect 7380 7404 7432 7410
rect 7852 7410 7880 8298
rect 7562 7375 7564 7384
rect 7380 7346 7432 7352
rect 7616 7375 7618 7384
rect 7840 7404 7892 7410
rect 7564 7346 7616 7352
rect 7840 7346 7892 7352
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7116 6934 7144 7278
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7392 6322 7420 6666
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7116 5710 7144 6258
rect 7576 6254 7604 7346
rect 7944 7342 7972 8978
rect 8220 8838 8248 9522
rect 8312 9364 8340 9646
rect 8588 9586 8616 9930
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8680 9518 8708 14334
rect 9770 14200 9826 15000
rect 10874 14200 10930 15000
rect 12070 14200 12126 15000
rect 13174 14200 13230 15000
rect 14370 14200 14426 15000
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 8956 13518 9260 13546
rect 9416 13530 9444 13806
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12442 8800 13194
rect 8864 12850 8892 13262
rect 8956 12918 8984 13518
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9048 12986 9076 13330
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 9048 12850 9076 12922
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8864 12238 8892 12650
rect 8942 12472 8998 12481
rect 8942 12407 8998 12416
rect 8852 12232 8904 12238
rect 8758 12200 8814 12209
rect 8852 12174 8904 12180
rect 8956 12170 8984 12407
rect 9048 12238 9076 12786
rect 9140 12646 9168 12786
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9140 12345 9168 12378
rect 9126 12336 9182 12345
rect 9126 12271 9182 12280
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8758 12135 8814 12144
rect 8944 12164 8996 12170
rect 8772 11762 8800 12135
rect 8944 12106 8996 12112
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 11626 8984 11698
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8760 11552 8812 11558
rect 8812 11512 8892 11540
rect 8760 11494 8812 11500
rect 8758 10976 8814 10985
rect 8758 10911 8814 10920
rect 8772 10742 8800 10911
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8760 10600 8812 10606
rect 8864 10588 8892 11512
rect 8956 10724 8984 11562
rect 9048 11082 9076 12038
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11354 9168 11494
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9232 11082 9260 13518
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9678 13424 9734 13433
rect 9324 12832 9352 13398
rect 9508 13190 9536 13398
rect 9678 13359 9734 13368
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12844 9456 12850
rect 9324 12804 9404 12832
rect 9324 12306 9352 12804
rect 9404 12786 9456 12792
rect 9508 12374 9536 13126
rect 9692 12918 9720 13359
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9678 12744 9734 12753
rect 9678 12679 9734 12688
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9508 12102 9536 12310
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11286 9444 11630
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9600 11200 9628 12582
rect 9692 12170 9720 12679
rect 9784 12186 9812 14200
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 13258 9996 13738
rect 10232 13320 10284 13326
rect 10284 13280 10364 13308
rect 10232 13262 10284 13268
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 10336 12986 10364 13280
rect 10888 13258 10916 14200
rect 12084 13870 12112 14200
rect 12072 13864 12124 13870
rect 11992 13824 12072 13852
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12374 10088 12650
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10428 12442 10456 12582
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10612 12306 10640 13126
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10888 12714 10916 12786
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 9784 12170 10548 12186
rect 9680 12164 9732 12170
rect 9784 12164 10560 12170
rect 9784 12158 10508 12164
rect 9680 12106 9732 12112
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9678 11792 9734 11801
rect 10060 11762 10088 12038
rect 9678 11727 9680 11736
rect 9732 11727 9734 11736
rect 9772 11756 9824 11762
rect 9680 11698 9732 11704
rect 9772 11698 9824 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9508 11172 9628 11200
rect 9508 11082 9536 11172
rect 9586 11112 9642 11121
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9496 11076 9548 11082
rect 9586 11047 9642 11056
rect 9496 11018 9548 11024
rect 9508 10985 9536 11018
rect 9600 11014 9628 11047
rect 9588 11008 9640 11014
rect 9494 10976 9550 10985
rect 9588 10950 9640 10956
rect 9494 10911 9550 10920
rect 9692 10826 9720 11698
rect 9784 11150 9812 11698
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 11150 9904 11222
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10048 11144 10100 11150
rect 10152 11121 10180 11290
rect 10048 11086 10100 11092
rect 10138 11112 10194 11121
rect 9508 10798 9720 10826
rect 9036 10736 9088 10742
rect 8956 10696 9036 10724
rect 9508 10690 9536 10798
rect 9784 10742 9812 11086
rect 9088 10684 9168 10690
rect 9036 10678 9168 10684
rect 9048 10662 9168 10678
rect 8864 10560 9076 10588
rect 8760 10542 8812 10548
rect 8772 9722 8800 10542
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8772 9586 8800 9658
rect 8864 9654 8892 10406
rect 9048 10266 9076 10560
rect 9140 10470 9168 10662
rect 9232 10662 9536 10690
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10668 9732 10674
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8760 9376 8812 9382
rect 8312 9336 8760 9364
rect 8760 9318 8812 9324
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8668 8968 8720 8974
rect 8666 8936 8668 8945
rect 8720 8936 8722 8945
rect 8666 8871 8722 8880
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8404 7818 8432 8026
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7546 8156 7686
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8482 7440 8538 7449
rect 8208 7404 8260 7410
rect 8482 7375 8484 7384
rect 8208 7346 8260 7352
rect 8536 7375 8538 7384
rect 8484 7346 8536 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 6866 7972 7278
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8220 6798 8248 7346
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6866 8340 7278
rect 8496 7002 8524 7346
rect 8588 7342 8616 7754
rect 8772 7750 8800 9046
rect 8864 8974 8892 9114
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8956 8922 8984 9998
rect 9048 9110 9076 10202
rect 9232 10062 9260 10662
rect 9680 10610 9732 10616
rect 9588 10600 9640 10606
rect 9586 10568 9588 10577
rect 9640 10568 9642 10577
rect 9586 10503 9642 10512
rect 9404 10464 9456 10470
rect 9324 10412 9404 10418
rect 9588 10464 9640 10470
rect 9324 10406 9456 10412
rect 9586 10432 9588 10441
rect 9640 10432 9642 10441
rect 9324 10390 9444 10406
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9324 9926 9352 10390
rect 9586 10367 9642 10376
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 9036 8968 9088 8974
rect 8956 8916 9036 8922
rect 8956 8910 9088 8916
rect 8864 8820 8892 8910
rect 8956 8894 9076 8910
rect 9140 8906 9168 9522
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8864 8792 8984 8820
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8680 7478 8708 7686
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8588 6798 8616 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8208 6792 8260 6798
rect 8036 6740 8208 6746
rect 8036 6734 8260 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8036 6718 8248 6734
rect 8036 6322 8064 6718
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8588 6458 8616 6734
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8680 6322 8708 6802
rect 8772 6798 8800 7278
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6322 8800 6598
rect 8864 6458 8892 7482
rect 8956 7188 8984 8792
rect 9048 7342 9076 8894
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9140 7954 9168 8434
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9140 7449 9168 7754
rect 9126 7440 9182 7449
rect 9232 7410 9260 9454
rect 9324 8838 9352 9862
rect 9416 9625 9444 9998
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9722 9536 9862
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9402 9616 9458 9625
rect 9600 9586 9628 9998
rect 9692 9586 9720 10610
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9402 9551 9458 9560
rect 9588 9580 9640 9586
rect 9416 9110 9444 9551
rect 9588 9522 9640 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9600 9110 9628 9522
rect 9692 9450 9720 9522
rect 9784 9518 9812 9930
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 9178 9720 9386
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9692 8974 9720 9007
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9416 8838 9444 8910
rect 9876 8906 9904 11086
rect 10060 11014 10088 11086
rect 10138 11047 10194 11056
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10130 9996 10610
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9968 9722 9996 9930
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9954 9616 10010 9625
rect 9954 9551 9956 9560
rect 10008 9551 10010 9560
rect 9956 9522 10008 9528
rect 10060 9110 10088 10950
rect 10152 9178 10180 11047
rect 10244 10130 10272 12158
rect 10508 12106 10560 12112
rect 10980 12102 11008 12922
rect 11164 12782 11192 13262
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10336 11558 10364 12038
rect 10690 11928 10746 11937
rect 10690 11863 10692 11872
rect 10744 11863 10746 11872
rect 10692 11834 10744 11840
rect 10508 11824 10560 11830
rect 10414 11792 10470 11801
rect 10560 11784 10640 11812
rect 10508 11766 10560 11772
rect 10414 11727 10470 11736
rect 10428 11626 10456 11727
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10336 9926 10364 10474
rect 10428 10266 10456 10610
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9404 8832 9456 8838
rect 9968 8809 9996 8910
rect 9404 8774 9456 8780
rect 9954 8800 10010 8809
rect 9324 8090 9352 8774
rect 9954 8735 10010 8744
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9126 7375 9182 7384
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8956 7160 9168 7188
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 9048 6390 9076 6598
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8496 5778 8524 6122
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8588 5766 8800 5794
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 4826 7328 5102
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7760 4690 7788 5510
rect 7944 4690 7972 5714
rect 8588 5642 8616 5766
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4826 8524 5170
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6932 3602 6960 4082
rect 7944 4078 7972 4490
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8588 4282 8616 5238
rect 8680 5030 8708 5578
rect 8772 5166 8800 5766
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5302 8892 5646
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4622 8708 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8772 4554 8800 4762
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 4140 8536 4146
rect 8668 4140 8720 4146
rect 8536 4100 8616 4128
rect 8484 4082 8536 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 5908 1488 5960 1494
rect 5908 1430 5960 1436
rect 5920 1358 5948 1430
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 5356 1284 5408 1290
rect 5356 1226 5408 1232
rect 6012 950 6040 1906
rect 6564 1766 6592 2994
rect 6656 1970 6684 3130
rect 6932 3058 6960 3334
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7116 2310 7144 3062
rect 7208 3058 7236 3606
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3194 7512 3334
rect 7944 3194 7972 3402
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8128 3058 8156 3878
rect 8404 3602 8432 4014
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8588 3194 8616 4100
rect 8668 4082 8720 4088
rect 8680 3738 8708 4082
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8772 3602 8800 4014
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8956 3670 8984 3946
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3194 8800 3538
rect 8576 3188 8628 3194
rect 8220 3148 8432 3176
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2378 7236 2858
rect 7484 2774 7512 2994
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7484 2746 7604 2774
rect 7576 2446 7604 2746
rect 7760 2446 7788 2926
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 6552 1420 6604 1426
rect 6552 1362 6604 1368
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 6564 1306 6592 1362
rect 7024 1306 7052 1362
rect 7116 1358 7144 1702
rect 7300 1426 7328 2246
rect 7484 1426 7512 2382
rect 7576 1494 7604 2382
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8036 2038 8064 2246
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 8024 2032 8076 2038
rect 8024 1974 8076 1980
rect 7564 1488 7616 1494
rect 7564 1430 7616 1436
rect 7852 1426 7880 1974
rect 8128 1850 8156 2994
rect 8220 2990 8248 3148
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8312 2514 8340 2994
rect 8404 2650 8432 3148
rect 8576 3130 8628 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8588 2650 8616 2926
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8772 1986 8800 3130
rect 9048 2774 9076 6054
rect 9140 5166 9168 7160
rect 9232 5914 9260 7346
rect 9324 6254 9352 8026
rect 9416 7868 9444 8434
rect 9496 7880 9548 7886
rect 9416 7840 9496 7868
rect 9416 7546 9444 7840
rect 9496 7822 9548 7828
rect 9600 7698 9628 8434
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9508 7670 9628 7698
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9508 7478 9536 7670
rect 9496 7472 9548 7478
rect 9416 7420 9496 7426
rect 9416 7414 9548 7420
rect 9416 7398 9536 7414
rect 9416 7018 9444 7398
rect 9416 6990 9536 7018
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9232 5234 9260 5850
rect 9416 5846 9444 6870
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9416 5710 9444 5782
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9324 4826 9352 5646
rect 9508 5370 9536 6990
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 5846 9720 6734
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9692 5302 9720 5782
rect 9784 5574 9812 8366
rect 9876 7410 9904 8570
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6934 9904 7210
rect 9968 7002 9996 8434
rect 10060 7886 10088 9046
rect 10152 8566 10180 9114
rect 10232 8968 10284 8974
rect 10230 8936 10232 8945
rect 10284 8936 10286 8945
rect 10230 8871 10286 8880
rect 10230 8800 10286 8809
rect 10230 8735 10286 8744
rect 10244 8566 10272 8735
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10152 7410 10180 8502
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9968 6458 9996 6938
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9876 5302 9904 5578
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9692 4758 9720 5238
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 4282 9260 4422
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9692 4214 9720 4694
rect 9968 4622 9996 6394
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5846 10088 6258
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3738 9168 4082
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 8956 2746 9076 2774
rect 8956 2514 8984 2746
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8496 1958 8800 1986
rect 8496 1902 8524 1958
rect 8484 1896 8536 1902
rect 8128 1822 8248 1850
rect 8484 1838 8536 1844
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 7288 1420 7340 1426
rect 7288 1362 7340 1368
rect 7472 1420 7524 1426
rect 7472 1362 7524 1368
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 8220 1358 8248 1822
rect 8496 1426 8524 1838
rect 8772 1494 8800 1838
rect 8760 1488 8812 1494
rect 8760 1430 8812 1436
rect 8484 1420 8536 1426
rect 8484 1362 8536 1368
rect 8956 1358 8984 2450
rect 9324 2310 9352 3674
rect 9416 3194 9444 3946
rect 9784 3738 9812 4014
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9876 3534 9904 4490
rect 9956 3936 10008 3942
rect 10060 3924 10088 5782
rect 10244 5710 10272 8502
rect 10336 8362 10364 9862
rect 10416 9580 10468 9586
rect 10520 9568 10548 11630
rect 10612 10538 10640 11784
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10876 11756 10928 11762
rect 10980 11744 11008 12038
rect 10928 11716 11008 11744
rect 10876 11698 10928 11704
rect 10704 11354 10732 11698
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10468 9540 10548 9568
rect 10416 9522 10468 9528
rect 10428 9110 10456 9522
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7478 10364 7822
rect 10428 7750 10456 9046
rect 10612 9024 10640 10474
rect 10796 10130 10824 11086
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10704 9654 10732 10066
rect 10888 10062 10916 11290
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9722 10916 9998
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 9036 10744 9042
rect 10612 8996 10692 9024
rect 10692 8978 10744 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8634 10640 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10692 6316 10744 6322
rect 10612 6276 10692 6304
rect 10324 6248 10376 6254
rect 10612 6236 10640 6276
rect 10692 6258 10744 6264
rect 10796 6254 10824 9318
rect 10888 9110 10916 9658
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10980 8906 11008 11716
rect 11072 9450 11100 12650
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11164 11354 11192 11766
rect 11256 11558 11284 12106
rect 11348 11762 11376 13466
rect 11808 13258 11836 13670
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12753 11560 12786
rect 11518 12744 11574 12753
rect 11518 12679 11574 12688
rect 11624 12238 11652 13194
rect 11808 12306 11836 13194
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11900 12238 11928 12718
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11665 11376 11698
rect 11334 11656 11390 11665
rect 11334 11591 11390 11600
rect 11244 11552 11296 11558
rect 11336 11552 11388 11558
rect 11244 11494 11296 11500
rect 11334 11520 11336 11529
rect 11388 11520 11390 11529
rect 11334 11455 11390 11464
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11440 11234 11468 11766
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11348 11206 11468 11234
rect 11532 11218 11560 11562
rect 11624 11286 11652 11834
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11520 11212 11572 11218
rect 11152 11144 11204 11150
rect 11150 11112 11152 11121
rect 11204 11112 11206 11121
rect 11150 11047 11206 11056
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10674 11192 10950
rect 11348 10810 11376 11206
rect 11520 11154 11572 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11244 10600 11296 10606
rect 11164 10548 11244 10554
rect 11164 10542 11296 10548
rect 11164 10526 11284 10542
rect 11164 9926 11192 10526
rect 11348 10266 11376 10610
rect 11440 10266 11468 11086
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11532 10713 11560 10746
rect 11518 10704 11574 10713
rect 11518 10639 11574 10648
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11164 9042 11192 9862
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10888 8566 10916 8842
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10376 6208 10640 6236
rect 10784 6248 10836 6254
rect 10324 6190 10376 6196
rect 10784 6190 10836 6196
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 4826 10272 5646
rect 10336 5642 10364 6054
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10152 4554 10180 4762
rect 10232 4616 10284 4622
rect 10336 4604 10364 5578
rect 10612 4690 10640 5850
rect 10980 5778 11008 7686
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11164 5166 11192 8434
rect 11256 7886 11284 10095
rect 11348 10062 11376 10202
rect 11532 10146 11560 10503
rect 11440 10118 11560 10146
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11440 9994 11468 10118
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11440 9722 11468 9930
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11336 9104 11388 9110
rect 11440 9081 11468 9658
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11336 9046 11388 9052
rect 11426 9072 11482 9081
rect 11348 8974 11376 9046
rect 11426 9007 11482 9016
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8634 11376 8910
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7342 11284 7822
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11348 6458 11376 8570
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11348 5302 11376 6394
rect 11440 5370 11468 9007
rect 11532 8498 11560 9522
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11624 8362 11652 10610
rect 11716 10470 11744 11698
rect 11992 11626 12020 13824
rect 12072 13806 12124 13812
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12084 12170 12112 13262
rect 12176 12850 12204 13262
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12918 12664 13194
rect 13188 13190 13216 14200
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 12912 12238 12940 12650
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12806 11792 12862 11801
rect 12072 11756 12124 11762
rect 12806 11727 12808 11736
rect 12072 11698 12124 11704
rect 12860 11727 12862 11736
rect 12808 11698 12860 11704
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11886 11384 11942 11393
rect 12084 11354 12112 11698
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 12728 11354 12756 11630
rect 11886 11319 11942 11328
rect 12072 11348 12124 11354
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9586 11744 9930
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 8838 11744 9522
rect 11704 8832 11756 8838
rect 11808 8809 11836 11086
rect 11704 8774 11756 8780
rect 11794 8800 11850 8809
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5642 11652 6122
rect 11716 5914 11744 8774
rect 11794 8735 11850 8744
rect 11808 8090 11836 8735
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11900 6866 11928 11319
rect 12072 11290 12124 11296
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12820 11150 12848 11698
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 11992 10810 12020 11086
rect 12912 11082 12940 12174
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12452 10713 12480 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10742 12756 10950
rect 12716 10736 12768 10742
rect 12438 10704 12494 10713
rect 12716 10678 12768 10684
rect 12438 10639 12494 10648
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12084 9568 12112 10542
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12728 9586 12756 10678
rect 13188 10674 13216 13126
rect 13280 12374 13308 13194
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13280 11830 13308 12310
rect 13372 11937 13400 13194
rect 14384 12442 14412 14200
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 13358 11928 13414 11937
rect 13358 11863 13414 11872
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12820 9722 12848 10542
rect 12912 10062 12940 10542
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 10198 13308 10474
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12164 9580 12216 9586
rect 12084 9540 12164 9568
rect 12084 9178 12112 9540
rect 12164 9522 12216 9528
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8362 12020 8910
rect 12360 8498 12388 8978
rect 13280 8974 13308 10134
rect 13372 10062 13400 11494
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10742 13492 10950
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13372 9586 13400 9998
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9042 13584 9318
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8634 12480 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12912 8566 12940 8842
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6390 11928 6666
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10284 4576 10364 4604
rect 10232 4558 10284 4564
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10152 3942 10180 4490
rect 11624 4282 11652 5170
rect 11900 4690 11928 5238
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4282 11928 4626
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11900 4146 11928 4218
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 10008 3896 10088 3924
rect 9956 3878 10008 3884
rect 10060 3670 10088 3896
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10152 3534 10180 3878
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9416 2446 9444 3130
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 2122 9352 2246
rect 9324 2106 9444 2122
rect 9324 2100 9456 2106
rect 9324 2094 9404 2100
rect 9404 2042 9456 2048
rect 9416 1358 9444 2042
rect 9508 1766 9536 2518
rect 9600 2514 9628 3334
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2514 9720 2994
rect 10336 2650 10364 3674
rect 11440 3602 11468 4082
rect 11900 3738 11928 4082
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3194 10640 3334
rect 10704 3194 10732 3402
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 11440 3058 11468 3538
rect 11900 3194 11928 3674
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 3058 11928 3130
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9496 1760 9548 1766
rect 9496 1702 9548 1708
rect 9508 1562 9536 1702
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 6564 1278 7052 1306
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8944 1352 8996 1358
rect 8944 1294 8996 1300
rect 9404 1352 9456 1358
rect 9600 1306 9628 2450
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10428 2038 10456 2382
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10428 1426 10456 1974
rect 10704 1970 10732 2586
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10692 1964 10744 1970
rect 10692 1906 10744 1912
rect 10704 1766 10732 1906
rect 10692 1760 10744 1766
rect 10692 1702 10744 1708
rect 10416 1420 10468 1426
rect 10416 1362 10468 1368
rect 10888 1358 10916 2042
rect 10980 1970 11008 2994
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11716 2378 11744 2858
rect 11992 2774 12020 8298
rect 12084 7478 12112 8298
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12912 7886 12940 8366
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12072 7336 12124 7342
rect 12176 7324 12204 7754
rect 12124 7296 12204 7324
rect 12254 7304 12310 7313
rect 12072 7278 12124 7284
rect 12084 6322 12112 7278
rect 12254 7239 12256 7248
rect 12308 7239 12310 7248
rect 12256 7210 12308 7216
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12912 6934 12940 7822
rect 13188 7206 13216 7958
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12900 6928 12952 6934
rect 12952 6886 13032 6914
rect 12900 6870 12952 6876
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12360 6322 12388 6734
rect 13004 6390 13032 6886
rect 13464 6798 13492 8842
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12084 6186 12112 6258
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12084 4622 12112 6122
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 13280 5914 13308 6190
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5302 13216 5510
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12636 4622 12664 5170
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12084 4146 12112 4558
rect 12636 4214 12664 4558
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12728 4146 12756 4966
rect 13188 4758 13216 5238
rect 13464 5216 13492 6734
rect 13556 6225 13584 8978
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13544 5228 13596 5234
rect 13464 5188 13544 5216
rect 13544 5170 13596 5176
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13556 4622 13584 5170
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 12820 3738 12848 4218
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3942 13584 4082
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3777 13584 3878
rect 13542 3768 13598 3777
rect 12808 3732 12860 3738
rect 13542 3703 13598 3712
rect 12808 3674 12860 3680
rect 12820 3534 12848 3674
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 11900 2746 12020 2774
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 10980 1834 11008 1906
rect 11796 1896 11848 1902
rect 11796 1838 11848 1844
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 10980 1426 11008 1770
rect 11612 1760 11664 1766
rect 11612 1702 11664 1708
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 9404 1294 9456 1300
rect 8024 1284 8076 1290
rect 8024 1226 8076 1232
rect 6460 1216 6512 1222
rect 6460 1158 6512 1164
rect 6472 1018 6500 1158
rect 8036 1018 8064 1226
rect 6460 1012 6512 1018
rect 6460 954 6512 960
rect 8024 1012 8076 1018
rect 8024 954 8076 960
rect 8128 950 8156 1294
rect 9508 1290 9628 1306
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 11164 1290 11192 1498
rect 11624 1358 11652 1702
rect 11808 1562 11836 1838
rect 11796 1556 11848 1562
rect 11796 1498 11848 1504
rect 11612 1352 11664 1358
rect 11900 1329 11928 2746
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12636 2582 12664 2994
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12728 2446 12756 2926
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13188 2106 13216 2450
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11992 1562 12020 1702
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 12084 1358 12112 1974
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 12072 1352 12124 1358
rect 11612 1294 11664 1300
rect 11886 1320 11942 1329
rect 9496 1284 9628 1290
rect 9548 1278 9628 1284
rect 11152 1284 11204 1290
rect 9496 1226 9548 1232
rect 12072 1294 12124 1300
rect 11886 1255 11942 1264
rect 11152 1226 11204 1232
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 4436 944 4488 950
rect 4436 886 4488 892
rect 6000 944 6052 950
rect 6000 886 6052 892
rect 8116 944 8168 950
rect 8116 886 8168 892
rect 11164 800 11192 1226
rect 2778 504 2834 513
rect 2778 439 2834 448
rect 3698 0 3754 800
rect 11150 0 11206 800
<< via2 >>
rect 3698 14456 3754 14512
rect 1398 12552 1454 12608
rect 3054 11600 3110 11656
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 3790 13504 3846 13560
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4342 12008 4398 12064
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 3330 9696 3386 9752
rect 5354 12824 5410 12880
rect 6918 12824 6974 12880
rect 6550 12164 6606 12200
rect 6550 12144 6552 12164
rect 6552 12144 6604 12164
rect 6604 12144 6606 12164
rect 6550 11772 6552 11792
rect 6552 11772 6604 11792
rect 6604 11772 6606 11792
rect 6550 11736 6606 11772
rect 6550 11464 6606 11520
rect 7194 12436 7250 12472
rect 7194 12416 7196 12436
rect 7196 12416 7248 12436
rect 7248 12416 7250 12436
rect 7286 11872 7342 11928
rect 6734 11736 6790 11792
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 7194 11736 7250 11792
rect 7102 11600 7158 11656
rect 6826 11348 6882 11384
rect 6826 11328 6828 11348
rect 6828 11328 6880 11348
rect 6880 11328 6882 11348
rect 6550 9580 6606 9616
rect 6550 9560 6552 9580
rect 6552 9560 6604 9580
rect 6604 9560 6606 9580
rect 2226 7928 2282 7984
rect 1398 6060 1400 6080
rect 1400 6060 1452 6080
rect 1452 6060 1454 6080
rect 1398 6024 1454 6060
rect 1766 5072 1822 5128
rect 1398 4120 1454 4176
rect 3882 8780 3884 8800
rect 3884 8780 3936 8800
rect 3936 8780 3938 8800
rect 3882 8744 3938 8780
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1490 3168 1546 3224
rect 1766 2216 1822 2272
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6996 4122 7032
rect 4066 6976 4068 6996
rect 4068 6976 4120 6996
rect 4120 6976 4122 6996
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5814 7248 5870 7304
rect 7378 10920 7434 10976
rect 6734 10376 6790 10432
rect 7378 10260 7434 10296
rect 7378 10240 7380 10260
rect 7380 10240 7432 10260
rect 7432 10240 7434 10260
rect 7286 10104 7342 10160
rect 7378 9560 7434 9616
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 3422 1264 3478 1320
rect 7562 12008 7618 12064
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8574 12824 8630 12880
rect 8390 12280 8446 12336
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 8022 11872 8078 11928
rect 8390 11620 8446 11656
rect 8390 11600 8392 11620
rect 8392 11600 8444 11620
rect 8444 11600 8446 11620
rect 7930 11056 7986 11112
rect 7838 10920 7894 10976
rect 7746 9560 7802 9616
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8114 10240 8170 10296
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 7562 7404 7618 7440
rect 7562 7384 7564 7404
rect 7564 7384 7616 7404
rect 7616 7384 7618 7404
rect 8942 12416 8998 12472
rect 8758 12144 8814 12200
rect 9126 12280 9182 12336
rect 8758 10920 8814 10976
rect 9678 13368 9734 13424
rect 9678 12688 9734 12744
rect 9678 11756 9734 11792
rect 9678 11736 9680 11756
rect 9680 11736 9732 11756
rect 9732 11736 9734 11756
rect 9586 11056 9642 11112
rect 9494 10920 9550 10976
rect 8666 8916 8668 8936
rect 8668 8916 8720 8936
rect 8720 8916 8722 8936
rect 8666 8880 8722 8916
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8482 7404 8538 7440
rect 8482 7384 8484 7404
rect 8484 7384 8536 7404
rect 8536 7384 8538 7404
rect 9586 10548 9588 10568
rect 9588 10548 9640 10568
rect 9640 10548 9642 10568
rect 9586 10512 9642 10548
rect 9586 10412 9588 10432
rect 9588 10412 9640 10432
rect 9640 10412 9642 10432
rect 9586 10376 9642 10412
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 9126 7384 9182 7440
rect 9402 9560 9458 9616
rect 9678 9016 9734 9072
rect 10138 11056 10194 11112
rect 9954 9580 10010 9616
rect 9954 9560 9956 9580
rect 9956 9560 10008 9580
rect 10008 9560 10010 9580
rect 10690 11892 10746 11928
rect 10690 11872 10692 11892
rect 10692 11872 10744 11892
rect 10744 11872 10746 11892
rect 10414 11736 10470 11792
rect 9954 8744 10010 8800
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 10230 8916 10232 8936
rect 10232 8916 10284 8936
rect 10284 8916 10286 8936
rect 10230 8880 10286 8916
rect 10230 8744 10286 8800
rect 11518 12688 11574 12744
rect 11334 11600 11390 11656
rect 11334 11500 11336 11520
rect 11336 11500 11388 11520
rect 11388 11500 11390 11520
rect 11334 11464 11390 11500
rect 11150 11092 11152 11112
rect 11152 11092 11204 11112
rect 11204 11092 11206 11112
rect 11150 11056 11206 11092
rect 11518 10648 11574 10704
rect 11518 10512 11574 10568
rect 11242 10104 11298 10160
rect 11426 9016 11482 9072
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 12806 11756 12862 11792
rect 12806 11736 12808 11756
rect 12808 11736 12860 11756
rect 12860 11736 12862 11756
rect 11886 11328 11942 11384
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 11794 8744 11850 8800
rect 12438 10648 12494 10704
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 13358 11872 13414 11928
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12254 7268 12310 7304
rect 12254 7248 12256 7268
rect 12256 7248 12308 7268
rect 12308 7248 12310 7268
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 13542 6160 13598 6216
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 13542 3712 13598 3768
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 11886 1264 11942 1320
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 2778 448 2834 504
<< metal3 >>
rect 0 14514 800 14544
rect 3693 14514 3759 14517
rect 0 14512 3759 14514
rect 0 14456 3698 14512
rect 3754 14456 3759 14512
rect 0 14454 3759 14456
rect 0 14424 800 14454
rect 3693 14451 3759 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 3785 13562 3851 13565
rect 0 13560 3851 13562
rect 0 13504 3790 13560
rect 3846 13504 3851 13560
rect 0 13502 3851 13504
rect 0 13472 800 13502
rect 3785 13499 3851 13502
rect 9673 13426 9739 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 9673 13424 12818 13426
rect 9673 13368 9678 13424
rect 9734 13368 12818 13424
rect 9673 13366 12818 13368
rect 9673 13363 9739 13366
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 5349 12882 5415 12885
rect 6913 12882 6979 12885
rect 8569 12882 8635 12885
rect 5349 12880 8635 12882
rect 5349 12824 5354 12880
rect 5410 12824 6918 12880
rect 6974 12824 8574 12880
rect 8630 12824 8635 12880
rect 5349 12822 8635 12824
rect 5349 12819 5415 12822
rect 6913 12819 6979 12822
rect 8569 12819 8635 12822
rect 9673 12746 9739 12749
rect 11513 12746 11579 12749
rect 9673 12744 11579 12746
rect 9673 12688 9678 12744
rect 9734 12688 11518 12744
rect 11574 12688 11579 12744
rect 9673 12686 11579 12688
rect 9673 12683 9739 12686
rect 11513 12683 11579 12686
rect 0 12610 800 12640
rect 1393 12610 1459 12613
rect 0 12608 1459 12610
rect 0 12552 1398 12608
rect 1454 12552 1459 12608
rect 0 12550 1459 12552
rect 0 12520 800 12550
rect 1393 12547 1459 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 7189 12474 7255 12477
rect 8937 12474 9003 12477
rect 7189 12472 9003 12474
rect 7189 12416 7194 12472
rect 7250 12416 8942 12472
rect 8998 12416 9003 12472
rect 7189 12414 9003 12416
rect 7189 12411 7255 12414
rect 8937 12411 9003 12414
rect 8385 12338 8451 12341
rect 9121 12338 9187 12341
rect 8385 12336 9187 12338
rect 8385 12280 8390 12336
rect 8446 12280 9126 12336
rect 9182 12280 9187 12336
rect 8385 12278 9187 12280
rect 8385 12275 8451 12278
rect 9121 12275 9187 12278
rect 6545 12202 6611 12205
rect 8753 12202 8819 12205
rect 6545 12200 8819 12202
rect 6545 12144 6550 12200
rect 6606 12144 8758 12200
rect 8814 12144 8819 12200
rect 6545 12142 8819 12144
rect 6545 12139 6611 12142
rect 8753 12139 8819 12142
rect 4337 12066 4403 12069
rect 7557 12066 7623 12069
rect 4337 12064 7623 12066
rect 4337 12008 4342 12064
rect 4398 12008 7562 12064
rect 7618 12008 7623 12064
rect 4337 12006 7623 12008
rect 4337 12003 4403 12006
rect 7557 12003 7623 12006
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 7281 11930 7347 11933
rect 8017 11930 8083 11933
rect 7281 11928 8083 11930
rect 7281 11872 7286 11928
rect 7342 11872 8022 11928
rect 8078 11872 8083 11928
rect 7281 11870 8083 11872
rect 7281 11867 7347 11870
rect 8017 11867 8083 11870
rect 10685 11930 10751 11933
rect 13353 11930 13419 11933
rect 10685 11928 13419 11930
rect 10685 11872 10690 11928
rect 10746 11872 13358 11928
rect 13414 11872 13419 11928
rect 10685 11870 13419 11872
rect 10685 11867 10751 11870
rect 13353 11867 13419 11870
rect 6545 11794 6611 11797
rect 6729 11794 6795 11797
rect 7189 11794 7255 11797
rect 9673 11794 9739 11797
rect 6545 11792 9739 11794
rect 6545 11736 6550 11792
rect 6606 11736 6734 11792
rect 6790 11736 7194 11792
rect 7250 11736 9678 11792
rect 9734 11736 9739 11792
rect 6545 11734 9739 11736
rect 6545 11731 6611 11734
rect 6729 11731 6795 11734
rect 7189 11731 7255 11734
rect 9673 11731 9739 11734
rect 10409 11794 10475 11797
rect 12801 11794 12867 11797
rect 10409 11792 12867 11794
rect 10409 11736 10414 11792
rect 10470 11736 12806 11792
rect 12862 11736 12867 11792
rect 10409 11734 12867 11736
rect 10409 11731 10475 11734
rect 12801 11731 12867 11734
rect 0 11658 800 11688
rect 3049 11658 3115 11661
rect 0 11656 3115 11658
rect 0 11600 3054 11656
rect 3110 11600 3115 11656
rect 0 11598 3115 11600
rect 0 11568 800 11598
rect 3049 11595 3115 11598
rect 7097 11658 7163 11661
rect 8385 11658 8451 11661
rect 7097 11656 8451 11658
rect 7097 11600 7102 11656
rect 7158 11600 8390 11656
rect 8446 11600 8451 11656
rect 7097 11598 8451 11600
rect 7097 11595 7163 11598
rect 8385 11595 8451 11598
rect 11329 11658 11395 11661
rect 11329 11656 12082 11658
rect 11329 11600 11334 11656
rect 11390 11600 12082 11656
rect 11329 11598 12082 11600
rect 11329 11595 11395 11598
rect 6545 11522 6611 11525
rect 11329 11522 11395 11525
rect 6545 11520 11395 11522
rect 6545 11464 6550 11520
rect 6606 11464 11334 11520
rect 11390 11464 11395 11520
rect 6545 11462 11395 11464
rect 6545 11459 6611 11462
rect 11329 11459 11395 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 6821 11386 6887 11389
rect 11881 11386 11947 11389
rect 6821 11384 11947 11386
rect 6821 11328 6826 11384
rect 6882 11328 11886 11384
rect 11942 11328 11947 11384
rect 6821 11326 11947 11328
rect 6821 11323 6887 11326
rect 11881 11323 11947 11326
rect 12022 11250 12082 11598
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 14200 11250 15000 11280
rect 12022 11190 15000 11250
rect 14200 11160 15000 11190
rect 7925 11114 7991 11117
rect 9581 11114 9647 11117
rect 7925 11112 9647 11114
rect 7925 11056 7930 11112
rect 7986 11056 9586 11112
rect 9642 11056 9647 11112
rect 7925 11054 9647 11056
rect 7925 11051 7991 11054
rect 9581 11051 9647 11054
rect 10133 11114 10199 11117
rect 11145 11114 11211 11117
rect 10133 11112 11211 11114
rect 10133 11056 10138 11112
rect 10194 11056 11150 11112
rect 11206 11056 11211 11112
rect 10133 11054 11211 11056
rect 10133 11051 10199 11054
rect 11145 11051 11211 11054
rect 7373 10978 7439 10981
rect 7833 10978 7899 10981
rect 7373 10976 7899 10978
rect 7373 10920 7378 10976
rect 7434 10920 7838 10976
rect 7894 10920 7899 10976
rect 7373 10918 7899 10920
rect 7373 10915 7439 10918
rect 7833 10915 7899 10918
rect 8753 10978 8819 10981
rect 9489 10978 9555 10981
rect 8753 10976 9555 10978
rect 8753 10920 8758 10976
rect 8814 10920 9494 10976
rect 9550 10920 9555 10976
rect 8753 10918 9555 10920
rect 8753 10915 8819 10918
rect 9489 10915 9555 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 0 10706 800 10736
rect 1577 10706 1643 10709
rect 0 10704 1643 10706
rect 0 10648 1582 10704
rect 1638 10648 1643 10704
rect 0 10646 1643 10648
rect 0 10616 800 10646
rect 1577 10643 1643 10646
rect 11513 10706 11579 10709
rect 12433 10706 12499 10709
rect 11513 10704 12499 10706
rect 11513 10648 11518 10704
rect 11574 10648 12438 10704
rect 12494 10648 12499 10704
rect 11513 10646 12499 10648
rect 11513 10643 11579 10646
rect 12433 10643 12499 10646
rect 9581 10570 9647 10573
rect 11513 10570 11579 10573
rect 9581 10568 11579 10570
rect 9581 10512 9586 10568
rect 9642 10512 11518 10568
rect 11574 10512 11579 10568
rect 9581 10510 11579 10512
rect 9581 10507 9647 10510
rect 11513 10507 11579 10510
rect 6729 10434 6795 10437
rect 9581 10434 9647 10437
rect 6729 10432 9647 10434
rect 6729 10376 6734 10432
rect 6790 10376 9586 10432
rect 9642 10376 9647 10432
rect 6729 10374 9647 10376
rect 6729 10371 6795 10374
rect 9581 10371 9647 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 7373 10298 7439 10301
rect 8109 10298 8175 10301
rect 7373 10296 8175 10298
rect 7373 10240 7378 10296
rect 7434 10240 8114 10296
rect 8170 10240 8175 10296
rect 7373 10238 8175 10240
rect 7373 10235 7439 10238
rect 8109 10235 8175 10238
rect 7281 10162 7347 10165
rect 11237 10162 11303 10165
rect 7281 10160 11303 10162
rect 7281 10104 7286 10160
rect 7342 10104 11242 10160
rect 11298 10104 11303 10160
rect 7281 10102 11303 10104
rect 7281 10099 7347 10102
rect 11237 10099 11303 10102
rect 8210 9824 8526 9825
rect 0 9754 800 9784
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 3325 9754 3391 9757
rect 0 9752 3391 9754
rect 0 9696 3330 9752
rect 3386 9696 3391 9752
rect 0 9694 3391 9696
rect 0 9664 800 9694
rect 3325 9691 3391 9694
rect 6545 9618 6611 9621
rect 7373 9618 7439 9621
rect 7741 9618 7807 9621
rect 6545 9616 7807 9618
rect 6545 9560 6550 9616
rect 6606 9560 7378 9616
rect 7434 9560 7746 9616
rect 7802 9560 7807 9616
rect 6545 9558 7807 9560
rect 6545 9555 6611 9558
rect 7373 9555 7439 9558
rect 7741 9555 7807 9558
rect 9397 9618 9463 9621
rect 9949 9618 10015 9621
rect 9397 9616 10015 9618
rect 9397 9560 9402 9616
rect 9458 9560 9954 9616
rect 10010 9560 10015 9616
rect 9397 9558 10015 9560
rect 9397 9555 9463 9558
rect 9949 9555 10015 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 9673 9074 9739 9077
rect 11421 9074 11487 9077
rect 9673 9072 11487 9074
rect 9673 9016 9678 9072
rect 9734 9016 11426 9072
rect 11482 9016 11487 9072
rect 9673 9014 11487 9016
rect 9673 9011 9739 9014
rect 11421 9011 11487 9014
rect 8661 8938 8727 8941
rect 10225 8938 10291 8941
rect 8661 8936 10291 8938
rect 8661 8880 8666 8936
rect 8722 8880 10230 8936
rect 10286 8880 10291 8936
rect 8661 8878 10291 8880
rect 8661 8875 8727 8878
rect 10225 8875 10291 8878
rect 0 8802 800 8832
rect 3877 8802 3943 8805
rect 0 8800 3943 8802
rect 0 8744 3882 8800
rect 3938 8744 3943 8800
rect 0 8742 3943 8744
rect 0 8712 800 8742
rect 3877 8739 3943 8742
rect 9949 8802 10015 8805
rect 10225 8802 10291 8805
rect 9949 8800 10291 8802
rect 9949 8744 9954 8800
rect 10010 8744 10230 8800
rect 10286 8744 10291 8800
rect 9949 8742 10291 8744
rect 9949 8739 10015 8742
rect 10225 8739 10291 8742
rect 11789 8802 11855 8805
rect 14200 8802 15000 8832
rect 11789 8800 15000 8802
rect 11789 8744 11794 8800
rect 11850 8744 15000 8800
rect 11789 8742 15000 8744
rect 11789 8739 11855 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 14200 8712 15000 8742
rect 8210 8671 8526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 0 7986 800 8016
rect 2221 7986 2287 7989
rect 0 7984 2287 7986
rect 0 7928 2226 7984
rect 2282 7928 2287 7984
rect 0 7926 2287 7928
rect 0 7896 800 7926
rect 2221 7923 2287 7926
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 7557 7442 7623 7445
rect 8477 7442 8543 7445
rect 9121 7442 9187 7445
rect 7557 7440 9187 7442
rect 7557 7384 7562 7440
rect 7618 7384 8482 7440
rect 8538 7384 9126 7440
rect 9182 7384 9187 7440
rect 7557 7382 9187 7384
rect 7557 7379 7623 7382
rect 8477 7379 8543 7382
rect 9121 7379 9187 7382
rect 5809 7306 5875 7309
rect 12249 7306 12315 7309
rect 5809 7304 12315 7306
rect 5809 7248 5814 7304
rect 5870 7248 12254 7304
rect 12310 7248 12315 7304
rect 5809 7246 12315 7248
rect 5809 7243 5875 7246
rect 12249 7243 12315 7246
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 4061 7034 4127 7037
rect 0 7032 4127 7034
rect 0 6976 4066 7032
rect 4122 6976 4127 7032
rect 0 6974 4127 6976
rect 0 6944 800 6974
rect 4061 6971 4127 6974
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 13537 6218 13603 6221
rect 14200 6218 15000 6248
rect 13537 6216 15000 6218
rect 13537 6160 13542 6216
rect 13598 6160 15000 6216
rect 13537 6158 15000 6160
rect 13537 6155 13603 6158
rect 14200 6128 15000 6158
rect 0 6082 800 6112
rect 1393 6082 1459 6085
rect 0 6080 1459 6082
rect 0 6024 1398 6080
rect 1454 6024 1459 6080
rect 0 6022 1459 6024
rect 0 5992 800 6022
rect 1393 6019 1459 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 0 5130 800 5160
rect 1761 5130 1827 5133
rect 0 5128 1827 5130
rect 0 5072 1766 5128
rect 1822 5072 1827 5128
rect 0 5070 1827 5072
rect 0 5040 800 5070
rect 1761 5067 1827 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 13537 3770 13603 3773
rect 14200 3770 15000 3800
rect 13537 3768 15000 3770
rect 13537 3712 13542 3768
rect 13598 3712 15000 3768
rect 13537 3710 15000 3712
rect 13537 3707 13603 3710
rect 14200 3680 15000 3710
rect 8210 3296 8526 3297
rect 0 3226 800 3256
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 1485 3226 1551 3229
rect 0 3224 1551 3226
rect 0 3168 1490 3224
rect 1546 3168 1551 3224
rect 0 3166 1551 3168
rect 0 3136 800 3166
rect 1485 3163 1551 3166
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 0 2274 800 2304
rect 1761 2274 1827 2277
rect 0 2272 1827 2274
rect 0 2216 1766 2272
rect 1822 2216 1827 2272
rect 0 2214 1827 2216
rect 0 2184 800 2214
rect 1761 2211 1827 2214
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 0 1322 800 1352
rect 3417 1322 3483 1325
rect 0 1320 3483 1322
rect 0 1264 3422 1320
rect 3478 1264 3483 1320
rect 0 1262 3483 1264
rect 0 1232 800 1262
rect 3417 1259 3483 1262
rect 11881 1322 11947 1325
rect 14200 1322 15000 1352
rect 11881 1320 15000 1322
rect 11881 1264 11886 1320
rect 11942 1264 15000 1320
rect 11881 1262 15000 1264
rect 11881 1259 11947 1262
rect 14200 1232 15000 1262
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 0 506 800 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 800 446
rect 2773 443 2839 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 8250 8252 8486 8488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 12250 4252 12486 4488
<< metal5 >>
rect 1056 12488 13940 12530
rect 1056 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13940 12488
rect 1056 12210 13940 12252
rect 1056 8488 13940 8530
rect 1056 8252 8250 8488
rect 8486 8252 13940 8488
rect 1056 8210 13940 8252
rect 1056 4488 13940 4530
rect 1056 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13940 4488
rect 1056 4210 13940 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A1 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1665323087
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B1
timestamp 1665323087
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B1
timestamp 1665323087
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B1
timestamp 1665323087
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1665323087
transform -1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1665323087
transform -1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1665323087
transform -1 0 1564 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B2
timestamp 1665323087
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B1
timestamp 1665323087
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1665323087
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1665323087
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 1665323087
transform -1 0 3680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A2
timestamp 1665323087
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A_N
timestamp 1665323087
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1665323087
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A2
timestamp 1665323087
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__B
timestamp 1665323087
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A1
timestamp 1665323087
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A2
timestamp 1665323087
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A1
timestamp 1665323087
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A2
timestamp 1665323087
transform -1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A1
timestamp 1665323087
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A2
timestamp 1665323087
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A1
timestamp 1665323087
transform 1 0 1472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A2
timestamp 1665323087
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A1
timestamp 1665323087
transform 1 0 2392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A2
timestamp 1665323087
transform -1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A1
timestamp 1665323087
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A2
timestamp 1665323087
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A1
timestamp 1665323087
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A2
timestamp 1665323087
transform -1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A1
timestamp 1665323087
transform 1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A2
timestamp 1665323087
transform 1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A_N
timestamp 1665323087
transform -1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__B
timestamp 1665323087
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A1
timestamp 1665323087
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__B1
timestamp 1665323087
transform -1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__B2
timestamp 1665323087
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A1
timestamp 1665323087
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A2
timestamp 1665323087
transform -1 0 6256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A1
timestamp 1665323087
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A2
timestamp 1665323087
transform -1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A1
timestamp 1665323087
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A2
timestamp 1665323087
transform -1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__B1
timestamp 1665323087
transform -1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__B2
timestamp 1665323087
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A1
timestamp 1665323087
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A2
timestamp 1665323087
transform -1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B1
timestamp 1665323087
transform -1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B2
timestamp 1665323087
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1665323087
transform 1 0 8372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A2
timestamp 1665323087
transform -1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1665323087
transform 1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A2
timestamp 1665323087
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B1
timestamp 1665323087
transform -1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B2
timestamp 1665323087
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A1
timestamp 1665323087
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A2
timestamp 1665323087
transform -1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__B1
timestamp 1665323087
transform -1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__B2
timestamp 1665323087
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1665323087
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A2
timestamp 1665323087
transform -1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A_N
timestamp 1665323087
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1665323087
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A2
timestamp 1665323087
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A1
timestamp 1665323087
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A2
timestamp 1665323087
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1665323087
transform 1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B
timestamp 1665323087
transform -1 0 6624 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1665323087
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1665323087
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1665323087
transform 1 0 12972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1665323087
transform 1 0 3588 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1665323087
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1665323087
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1665323087
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1665323087
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1665323087
transform 1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1665323087
transform 1 0 8096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1665323087
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1665323087
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1665323087
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1665323087
transform 1 0 13064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1665323087
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1665323087
transform 1 0 12512 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1665323087
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1665323087
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1665323087
transform 1 0 13064 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1665323087
transform 1 0 3404 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1665323087
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1665323087
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1665323087
transform 1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__D
timestamp 1665323087
transform -1 0 13064 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1665323087
transform 1 0 7820 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90
timestamp 1665323087
transform 1 0 9384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1665323087
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_50
timestamp 1665323087
transform 1 0 5704 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1665323087
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1665323087
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1665323087
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1665323087
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1665323087
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1665323087
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_42
timestamp 1665323087
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_49
timestamp 1665323087
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1665323087
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_109
timestamp 1665323087
transform 1 0 11132 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1665323087
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1665323087
transform 1 0 13524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1665323087
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 1665323087
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1665323087
transform 1 0 5888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1665323087
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1665323087
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_135
timestamp 1665323087
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp 1665323087
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1665323087
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_46
timestamp 1665323087
transform 1 0 5336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1665323087
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1665323087
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1665323087
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1665323087
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1665323087
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_39
timestamp 1665323087
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1665323087
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1665323087
transform 1 0 10212 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_121 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1665323087
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1665323087
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1665323087
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1665323087
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1665323087
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_50
timestamp 1665323087
transform 1 0 5704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 1665323087
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1665323087
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1665323087
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp 1665323087
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1665323087
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1665323087
transform 1 0 3864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1665323087
transform 1 0 5520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1665323087
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 1665323087
transform 1 0 7268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1665323087
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1665323087
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1665323087
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1665323087
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1665323087
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1665323087
transform 1 0 13524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_31
timestamp 1665323087
transform 1 0 3956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1665323087
transform 1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_94
timestamp 1665323087
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1665323087
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1665323087
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1665323087
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1665323087
transform 1 0 5520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_59
timestamp 1665323087
transform 1 0 6532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_5
timestamp 1665323087
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1665323087
transform 1 0 2300 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1665323087
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1665323087
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_107
timestamp 1665323087
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_130
timestamp 1665323087
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1665323087
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1665323087
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1665323087
transform 1 0 7544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1665323087
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1665323087
transform 1 0 10212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1665323087
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1665323087
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_18
timestamp 1665323087
transform 1 0 2760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1665323087
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_78
timestamp 1665323087
transform 1 0 8280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1665323087
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1665323087
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1665323087
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1665323087
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1665323087
transform 1 0 12236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1665323087
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_17
timestamp 1665323087
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_40
timestamp 1665323087
transform 1 0 4784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1665323087
transform 1 0 7544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1665323087
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_122
timestamp 1665323087
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1665323087
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1665323087
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1665323087
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1665323087
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_54
timestamp 1665323087
transform 1 0 6072 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1665323087
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1665323087
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1665323087
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_25
timestamp 1665323087
transform 1 0 3404 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1665323087
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_60
timestamp 1665323087
transform 1 0 6624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_105
timestamp 1665323087
transform 1 0 10764 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _176_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1665323087
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1665323087
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1665323087
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1665323087
transform -1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _181_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13156 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _182_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13524 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _183_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1665323087
transform 1 0 4048 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1665323087
transform 1 0 4508 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1665323087
transform 1 0 4692 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1665323087
transform 1 0 2760 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _188_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3496 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _189_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _190_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2208 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _191_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3680 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1665323087
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _193_
timestamp 1665323087
transform -1 0 5336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _194_
timestamp 1665323087
transform -1 0 5888 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _195_
timestamp 1665323087
transform -1 0 4508 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _196_
timestamp 1665323087
transform -1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _197_
timestamp 1665323087
transform -1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _198_
timestamp 1665323087
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _199_
timestamp 1665323087
transform 1 0 1840 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _200_
timestamp 1665323087
transform -1 0 5520 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _201_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3128 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _202_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _203_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _204_
timestamp 1665323087
transform -1 0 2576 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _205_
timestamp 1665323087
transform -1 0 2116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _206_
timestamp 1665323087
transform -1 0 3404 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _207_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1665323087
transform -1 0 3680 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _209_
timestamp 1665323087
transform -1 0 3956 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _210_
timestamp 1665323087
transform -1 0 4048 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _211_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _212_
timestamp 1665323087
transform -1 0 4784 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _213_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2116 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _214_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _215_
timestamp 1665323087
transform 1 0 1472 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _216_
timestamp 1665323087
transform 1 0 1380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _217_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _218_
timestamp 1665323087
transform 1 0 3772 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _219_
timestamp 1665323087
transform -1 0 4876 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _220_
timestamp 1665323087
transform -1 0 1840 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _221_
timestamp 1665323087
transform 1 0 2300 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _222_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _223_
timestamp 1665323087
transform 1 0 3772 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _224_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _225_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2944 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _226_
timestamp 1665323087
transform 1 0 2116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _227_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3404 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _228_
timestamp 1665323087
transform -1 0 10948 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _229_
timestamp 1665323087
transform 1 0 10948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _230_
timestamp 1665323087
transform -1 0 7912 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _231_
timestamp 1665323087
transform 1 0 6348 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1665323087
transform -1 0 8832 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _233_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9844 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _234_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9568 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _235_
timestamp 1665323087
transform -1 0 2760 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _236_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1840 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _237_
timestamp 1665323087
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _238_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _239_
timestamp 1665323087
transform -1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _240_
timestamp 1665323087
transform 1 0 10948 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _241_
timestamp 1665323087
transform -1 0 10488 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _242_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9108 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _243_
timestamp 1665323087
transform -1 0 11040 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _244_
timestamp 1665323087
transform 1 0 7084 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _245_
timestamp 1665323087
transform -1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _246_
timestamp 1665323087
transform -1 0 8740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _247_
timestamp 1665323087
transform 1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _248_
timestamp 1665323087
transform -1 0 8372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _249_
timestamp 1665323087
transform -1 0 10948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _250_
timestamp 1665323087
transform 1 0 7452 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_2  _251_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _252_
timestamp 1665323087
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _253_
timestamp 1665323087
transform 1 0 7360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _254_
timestamp 1665323087
transform 1 0 5704 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _255_
timestamp 1665323087
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _256_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6624 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _257_
timestamp 1665323087
transform 1 0 6532 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _258_
timestamp 1665323087
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _259_
timestamp 1665323087
transform -1 0 10304 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1665323087
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _261_
timestamp 1665323087
transform 1 0 7912 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1665323087
transform -1 0 9844 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _263_
timestamp 1665323087
transform 1 0 9844 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _264_
timestamp 1665323087
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _265_
timestamp 1665323087
transform 1 0 9844 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _266_
timestamp 1665323087
transform 1 0 8648 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _267_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9384 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _268_
timestamp 1665323087
transform -1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _269_
timestamp 1665323087
transform 1 0 6716 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1665323087
transform 1 0 7268 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _271_
timestamp 1665323087
transform -1 0 10304 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _272_
timestamp 1665323087
transform 1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _273_
timestamp 1665323087
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _274_
timestamp 1665323087
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _275_
timestamp 1665323087
transform 1 0 5336 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _276_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6440 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _277_
timestamp 1665323087
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _278_
timestamp 1665323087
transform -1 0 6440 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _279_
timestamp 1665323087
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _280_
timestamp 1665323087
transform 1 0 8096 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _281_
timestamp 1665323087
transform 1 0 6992 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _282_
timestamp 1665323087
transform 1 0 6624 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _283_
timestamp 1665323087
transform 1 0 7452 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _284_
timestamp 1665323087
transform 1 0 5520 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1665323087
transform -1 0 11132 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1665323087
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _287_
timestamp 1665323087
transform -1 0 9384 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _288_
timestamp 1665323087
transform -1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _289_
timestamp 1665323087
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _290_
timestamp 1665323087
transform -1 0 8832 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _291_
timestamp 1665323087
transform -1 0 10212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _292_
timestamp 1665323087
transform 1 0 8648 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _293_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _294_
timestamp 1665323087
transform -1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _295_
timestamp 1665323087
transform -1 0 5060 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _296_
timestamp 1665323087
transform 1 0 10580 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _297_
timestamp 1665323087
transform 1 0 4876 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _298_
timestamp 1665323087
transform 1 0 7912 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _299_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _300_
timestamp 1665323087
transform -1 0 3680 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _301_
timestamp 1665323087
transform -1 0 6256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _302_
timestamp 1665323087
transform -1 0 2300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _303_
timestamp 1665323087
transform 1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _304_
timestamp 1665323087
transform 1 0 6440 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _305_
timestamp 1665323087
transform -1 0 4416 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _306_
timestamp 1665323087
transform -1 0 4600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _307_
timestamp 1665323087
transform -1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _308_
timestamp 1665323087
transform -1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _309_
timestamp 1665323087
transform 1 0 6716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _310_
timestamp 1665323087
transform 1 0 6624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _311_
timestamp 1665323087
transform 1 0 6808 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _312_
timestamp 1665323087
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _313_
timestamp 1665323087
transform 1 0 3956 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _314_
timestamp 1665323087
transform -1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _315_
timestamp 1665323087
transform -1 0 7452 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _316_
timestamp 1665323087
transform 1 0 5520 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _317_
timestamp 1665323087
transform 1 0 5888 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _318_
timestamp 1665323087
transform -1 0 7544 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _319_
timestamp 1665323087
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _320_
timestamp 1665323087
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _321_
timestamp 1665323087
transform 1 0 7452 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _322_
timestamp 1665323087
transform 1 0 7544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _323_
timestamp 1665323087
transform 1 0 11040 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _324_
timestamp 1665323087
transform -1 0 10212 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _325_
timestamp 1665323087
transform -1 0 11408 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _326_
timestamp 1665323087
transform -1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _327_
timestamp 1665323087
transform 1 0 10304 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _328_
timestamp 1665323087
transform -1 0 9200 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _329_
timestamp 1665323087
transform 1 0 7636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _330_
timestamp 1665323087
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _331_
timestamp 1665323087
transform -1 0 9016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _332_
timestamp 1665323087
transform 1 0 7544 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _333_
timestamp 1665323087
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _334_
timestamp 1665323087
transform 1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _335_
timestamp 1665323087
transform -1 0 10120 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _336_
timestamp 1665323087
transform 1 0 10212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _337_
timestamp 1665323087
transform 1 0 9844 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _338_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9568 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _339_
timestamp 1665323087
transform 1 0 10212 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _340_
timestamp 1665323087
transform 1 0 10120 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _341_
timestamp 1665323087
transform -1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _342_
timestamp 1665323087
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _343_
timestamp 1665323087
transform -1 0 8832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _344_
timestamp 1665323087
transform 1 0 11500 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _345_
timestamp 1665323087
transform -1 0 11408 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _346_
timestamp 1665323087
transform 1 0 7268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _347_
timestamp 1665323087
transform 1 0 10396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _348_
timestamp 1665323087
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _349_
timestamp 1665323087
transform 1 0 11500 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _350_
timestamp 1665323087
transform -1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _351_
timestamp 1665323087
transform 1 0 11776 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _352_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _353_
timestamp 1665323087
transform 1 0 12420 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _354_
timestamp 1665323087
transform 1 0 11040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _355_
timestamp 1665323087
transform 1 0 8372 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _356_
timestamp 1665323087
transform -1 0 10856 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _357_
timestamp 1665323087
transform -1 0 10212 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _358_
timestamp 1665323087
transform -1 0 12788 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _359_
timestamp 1665323087
transform 1 0 5796 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _360_
timestamp 1665323087
transform -1 0 8372 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _361_
timestamp 1665323087
transform -1 0 8280 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _362_
timestamp 1665323087
transform 1 0 6440 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _363_
timestamp 1665323087
transform 1 0 5612 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _364_
timestamp 1665323087
transform -1 0 12420 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _365_
timestamp 1665323087
transform -1 0 8740 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _366_
timestamp 1665323087
transform -1 0 12696 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _367_
timestamp 1665323087
transform -1 0 11960 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _368_
timestamp 1665323087
transform -1 0 12420 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _369_
timestamp 1665323087
transform -1 0 11960 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _370_
timestamp 1665323087
transform 1 0 6532 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _371_
timestamp 1665323087
transform -1 0 11316 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _372_
timestamp 1665323087
transform 1 0 11592 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _373_
timestamp 1665323087
transform -1 0 11960 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _374_
timestamp 1665323087
transform -1 0 12512 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _375_
timestamp 1665323087
transform 1 0 4232 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _376_
timestamp 1665323087
transform 1 0 2944 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _377_
timestamp 1665323087
transform 1 0 3956 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _378_
timestamp 1665323087
transform -1 0 3864 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _379_ $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8464 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _380_
timestamp 1665323087
transform 1 0 8280 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _381_
timestamp 1665323087
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _382_
timestamp 1665323087
transform 1 0 5520 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _383_
timestamp 1665323087
transform -1 0 8464 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _384_
timestamp 1665323087
transform -1 0 8832 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1665323087
transform -1 0 8280 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _386_
timestamp 1665323087
transform 1 0 4784 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1665323087
transform 1 0 9476 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1665323087
transform 1 0 6900 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _389_
timestamp 1665323087
transform 1 0 10304 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _390_
timestamp 1665323087
transform 1 0 10304 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1665323087
transform 1 0 9844 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1665323087
transform 1 0 9476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1665323087
transform 1 0 5796 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1665323087
transform 1 0 9476 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1665323087
transform 1 0 11500 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _396_
timestamp 1665323087
transform 1 0 10396 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _397_
timestamp 1665323087
transform 1 0 1748 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _398_
timestamp 1665323087
transform 1 0 3772 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _399_
timestamp 1665323087
transform 1 0 3772 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _400_
timestamp 1665323087
transform 1 0 3772 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _401_
timestamp 1665323087
transform 1 0 1748 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_16  clockp_buffer_0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3404 0 -1 2176
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  clockp_buffer_1
timestamp 1665323087
transform 1 0 1380 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4048 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1665323087
transform 1 0 4876 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3496 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4692 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1665323087
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1665323087
transform 1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1665323087
transform 1 0 4048 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1665323087
transform 1 0 5060 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1665323087
transform 1 0 3588 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1665323087
transform -1 0 6256 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1665323087
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1665323087
transform -1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1665323087
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1665323087
transform 1 0 2116 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1665323087
transform 1 0 2392 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1665323087
transform 1 0 1564 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1665323087
transform 1 0 2208 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1665323087
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1665323087
transform -1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1665323087
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1665323087
transform 1 0 1656 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1665323087
transform -1 0 2116 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1665323087
transform 1 0 1380 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1665323087
transform 1 0 1380 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1665323087
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1665323087
transform 1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1665323087
transform -1 0 3680 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1665323087
transform 1 0 2760 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1665323087
transform 1 0 2944 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1665323087
transform 1 0 2300 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1665323087
transform 1 0 2760 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1665323087
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1665323087
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1665323087
transform -1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1665323087
transform 1 0 3772 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1665323087
transform -1 0 5888 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1665323087
transform 1 0 3772 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1665323087
transform -1 0 5244 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1665323087
transform -1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1665323087
transform 1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1665323087
transform 1 0 5888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1665323087
transform 1 0 4600 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1665323087
transform 1 0 5244 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1665323087
transform 1 0 4600 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1665323087
transform 1 0 5060 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1665323087
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1665323087
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1665323087
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1665323087
transform 1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1665323087
transform 1 0 8188 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1665323087
transform 1 0 9292 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1665323087
transform 1 0 8096 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1665323087
transform 1 0 10488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1665323087
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1665323087
transform -1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1665323087
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1665323087
transform -1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1665323087
transform 1 0 11500 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1665323087
transform 1 0 10948 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1665323087
transform -1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1665323087
transform -1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1665323087
transform -1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1665323087
transform 1 0 12788 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1665323087
transform 1 0 12420 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1665323087
transform 1 0 12328 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1665323087
transform -1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1665323087
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1665323087
transform 1 0 12880 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1665323087
transform 1 0 12236 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1665323087
transform 1 0 12144 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1665323087
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1665323087
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1665323087
transform 1 0 12604 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1665323087
transform 1 0 12696 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1665323087
transform 1 0 12604 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1665323087
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6256 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1665323087
transform -1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1665323087
transform 1 0 1380 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1665323087
transform 1 0 11408 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1665323087
transform -1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1665323087
transform 1 0 11776 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1665323087
transform 1 0 12420 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1665323087
transform 1 0 11868 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1665323087
transform 1 0 12328 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1665323087
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12420 0 -1 7616
box -38 -48 498 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8210 13940 8530 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4210 13940 4530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12210 13940 12530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 3974 14200 4030 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 5170 14200 5226 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 6274 14200 6330 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 7470 14200 7526 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 8574 14200 8630 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 9770 14200 9826 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 10874 14200 10930 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 12070 14200 12126 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 13174 14200 13230 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 14200 13608 15000 13728 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 14200 11160 15000 11280 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 14200 8712 15000 8832 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 14200 6128 15000 6248 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 14200 3680 15000 3800 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 14200 1232 15000 1352 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 570 14200 626 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 1674 14200 1730 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 2870 14200 2926 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
