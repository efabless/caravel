magic
tech sky130A
magscale 1 2
timestamp 1665972027
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 113818 1007400 113824 1007412
rect 113146 1007372 113824 1007400
rect 106826 1007292 106832 1007344
rect 106884 1007332 106890 1007344
rect 113146 1007332 113174 1007372
rect 113818 1007360 113824 1007372
rect 113876 1007360 113882 1007412
rect 106884 1007304 113174 1007332
rect 106884 1007292 106890 1007304
rect 425514 1007088 425520 1007140
rect 425572 1007128 425578 1007140
rect 425572 1007100 441614 1007128
rect 425572 1007088 425578 1007100
rect 359734 1006952 359740 1007004
rect 359792 1006992 359798 1007004
rect 371234 1006992 371240 1007004
rect 359792 1006964 371240 1006992
rect 359792 1006952 359798 1006964
rect 371234 1006952 371240 1006964
rect 371292 1006952 371298 1007004
rect 428366 1006884 428372 1006936
rect 428424 1006924 428430 1006936
rect 428424 1006896 437474 1006924
rect 428424 1006884 428430 1006896
rect 359366 1006816 359372 1006868
rect 359424 1006856 359430 1006868
rect 367370 1006856 367376 1006868
rect 359424 1006828 367376 1006856
rect 359424 1006816 359430 1006828
rect 367370 1006816 367376 1006828
rect 367428 1006816 367434 1006868
rect 429194 1006748 429200 1006800
rect 429252 1006788 429258 1006800
rect 431862 1006788 431868 1006800
rect 429252 1006760 431868 1006788
rect 429252 1006748 429258 1006760
rect 431862 1006748 431868 1006760
rect 431920 1006748 431926 1006800
rect 437446 1006788 437474 1006896
rect 440234 1006788 440240 1006800
rect 437446 1006760 440240 1006788
rect 440234 1006748 440240 1006760
rect 440292 1006748 440298 1006800
rect 161750 1006680 161756 1006732
rect 161808 1006720 161814 1006732
rect 164878 1006720 164884 1006732
rect 161808 1006692 164884 1006720
rect 161808 1006680 161814 1006692
rect 164878 1006680 164884 1006692
rect 164936 1006680 164942 1006732
rect 361390 1006680 361396 1006732
rect 361448 1006720 361454 1006732
rect 376018 1006720 376024 1006732
rect 361448 1006692 376024 1006720
rect 361448 1006680 361454 1006692
rect 376018 1006680 376024 1006692
rect 376076 1006680 376082 1006732
rect 431678 1006652 431684 1006664
rect 412606 1006624 431684 1006652
rect 94498 1006544 94504 1006596
rect 94556 1006584 94562 1006596
rect 101950 1006584 101956 1006596
rect 94556 1006556 101956 1006584
rect 94556 1006544 94562 1006556
rect 101950 1006544 101956 1006556
rect 102008 1006544 102014 1006596
rect 145558 1006544 145564 1006596
rect 145616 1006584 145622 1006596
rect 153746 1006584 153752 1006596
rect 145616 1006556 153752 1006584
rect 145616 1006544 145622 1006556
rect 153746 1006544 153752 1006556
rect 153804 1006544 153810 1006596
rect 157426 1006544 157432 1006596
rect 157484 1006584 157490 1006596
rect 162302 1006584 162308 1006596
rect 157484 1006556 162308 1006584
rect 157484 1006544 157490 1006556
rect 162302 1006544 162308 1006556
rect 162360 1006544 162366 1006596
rect 162486 1006544 162492 1006596
rect 162544 1006584 162550 1006596
rect 173158 1006584 173164 1006596
rect 162544 1006556 173164 1006584
rect 162544 1006544 162550 1006556
rect 173158 1006544 173164 1006556
rect 173216 1006544 173222 1006596
rect 101582 1006408 101588 1006460
rect 101640 1006448 101646 1006460
rect 104802 1006448 104808 1006460
rect 101640 1006420 104808 1006448
rect 101640 1006408 101646 1006420
rect 104802 1006408 104808 1006420
rect 104860 1006408 104866 1006460
rect 145742 1006408 145748 1006460
rect 145800 1006448 145806 1006460
rect 152918 1006448 152924 1006460
rect 145800 1006420 152924 1006448
rect 145800 1006408 145806 1006420
rect 152918 1006408 152924 1006420
rect 152976 1006408 152982 1006460
rect 158254 1006408 158260 1006460
rect 158312 1006448 158318 1006460
rect 171778 1006448 171784 1006460
rect 158312 1006420 171784 1006448
rect 158312 1006408 158318 1006420
rect 171778 1006408 171784 1006420
rect 171836 1006408 171842 1006460
rect 247862 1006408 247868 1006460
rect 247920 1006448 247926 1006460
rect 256142 1006448 256148 1006460
rect 247920 1006420 256148 1006448
rect 247920 1006408 247926 1006420
rect 256142 1006408 256148 1006420
rect 256200 1006408 256206 1006460
rect 301498 1006408 301504 1006460
rect 301556 1006448 301562 1006460
rect 307754 1006448 307760 1006460
rect 301556 1006420 307760 1006448
rect 301556 1006408 301562 1006420
rect 307754 1006408 307760 1006420
rect 307812 1006408 307818 1006460
rect 360562 1006408 360568 1006460
rect 360620 1006448 360626 1006460
rect 367002 1006448 367008 1006460
rect 360620 1006420 367008 1006448
rect 360620 1006408 360626 1006420
rect 367002 1006408 367008 1006420
rect 367060 1006408 367066 1006460
rect 402238 1006408 402244 1006460
rect 402296 1006448 402302 1006460
rect 412606 1006448 412634 1006624
rect 431678 1006612 431684 1006624
rect 431736 1006612 431742 1006664
rect 441586 1006584 441614 1007100
rect 507854 1006884 507860 1006936
rect 507912 1006924 507918 1006936
rect 507912 1006896 509234 1006924
rect 507912 1006884 507918 1006896
rect 509206 1006856 509234 1006896
rect 520918 1006856 520924 1006868
rect 509206 1006828 520924 1006856
rect 520918 1006816 520924 1006828
rect 520976 1006816 520982 1006868
rect 505002 1006680 505008 1006732
rect 505060 1006720 505066 1006732
rect 518158 1006720 518164 1006732
rect 505060 1006692 518164 1006720
rect 505060 1006680 505066 1006692
rect 518158 1006680 518164 1006692
rect 518216 1006680 518222 1006732
rect 555970 1006680 555976 1006732
rect 556028 1006720 556034 1006732
rect 558822 1006720 558828 1006732
rect 556028 1006692 558828 1006720
rect 556028 1006680 556034 1006692
rect 558822 1006680 558828 1006692
rect 558880 1006680 558886 1006732
rect 467098 1006584 467104 1006596
rect 441586 1006556 467104 1006584
rect 467098 1006544 467104 1006556
rect 467156 1006544 467162 1006596
rect 501322 1006544 501328 1006596
rect 501380 1006584 501386 1006596
rect 514754 1006584 514760 1006596
rect 501380 1006556 514760 1006584
rect 501380 1006544 501386 1006556
rect 514754 1006544 514760 1006556
rect 514812 1006544 514818 1006596
rect 556798 1006544 556804 1006596
rect 556856 1006584 556862 1006596
rect 567838 1006584 567844 1006596
rect 556856 1006556 567844 1006584
rect 556856 1006544 556862 1006556
rect 567838 1006544 567844 1006556
rect 567896 1006544 567902 1006596
rect 402296 1006420 412634 1006448
rect 402296 1006408 402302 1006420
rect 429194 1006408 429200 1006460
rect 429252 1006448 429258 1006460
rect 429252 1006420 429424 1006448
rect 429252 1006408 429258 1006420
rect 93118 1006272 93124 1006324
rect 93176 1006312 93182 1006324
rect 100294 1006312 100300 1006324
rect 93176 1006284 100300 1006312
rect 93176 1006272 93182 1006284
rect 100294 1006272 100300 1006284
rect 100352 1006272 100358 1006324
rect 144270 1006272 144276 1006324
rect 144328 1006312 144334 1006324
rect 144328 1006284 151814 1006312
rect 144328 1006272 144334 1006284
rect 93302 1006136 93308 1006188
rect 93360 1006176 93366 1006188
rect 93360 1006148 98500 1006176
rect 93360 1006136 93366 1006148
rect 94682 1006000 94688 1006052
rect 94740 1006040 94746 1006052
rect 98270 1006040 98276 1006052
rect 94740 1006012 98276 1006040
rect 94740 1006000 94746 1006012
rect 98270 1006000 98276 1006012
rect 98328 1006000 98334 1006052
rect 98472 1006040 98500 1006148
rect 101398 1006136 101404 1006188
rect 101456 1006176 101462 1006188
rect 103974 1006176 103980 1006188
rect 101456 1006148 103980 1006176
rect 101456 1006136 101462 1006148
rect 103974 1006136 103980 1006148
rect 104032 1006136 104038 1006188
rect 105998 1006136 106004 1006188
rect 106056 1006176 106062 1006188
rect 124858 1006176 124864 1006188
rect 106056 1006148 124864 1006176
rect 106056 1006136 106062 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 144730 1006136 144736 1006188
rect 144788 1006176 144794 1006188
rect 151262 1006176 151268 1006188
rect 144788 1006148 151268 1006176
rect 144788 1006136 144794 1006148
rect 151262 1006136 151268 1006148
rect 151320 1006136 151326 1006188
rect 151786 1006176 151814 1006284
rect 158622 1006272 158628 1006324
rect 158680 1006312 158686 1006324
rect 162486 1006312 162492 1006324
rect 158680 1006284 162492 1006312
rect 158680 1006272 158686 1006284
rect 162486 1006272 162492 1006284
rect 162544 1006272 162550 1006324
rect 255958 1006272 255964 1006324
rect 256016 1006312 256022 1006324
rect 258994 1006312 259000 1006324
rect 256016 1006284 259000 1006312
rect 256016 1006272 256022 1006284
rect 258994 1006272 259000 1006284
rect 259052 1006272 259058 1006324
rect 300486 1006272 300492 1006324
rect 300544 1006312 300550 1006324
rect 306926 1006312 306932 1006324
rect 300544 1006284 306932 1006312
rect 300544 1006272 300550 1006284
rect 306926 1006272 306932 1006284
rect 306984 1006272 306990 1006324
rect 314654 1006272 314660 1006324
rect 314712 1006312 314718 1006324
rect 319438 1006312 319444 1006324
rect 314712 1006284 319444 1006312
rect 314712 1006272 314718 1006284
rect 319438 1006272 319444 1006284
rect 319496 1006272 319502 1006324
rect 354858 1006272 354864 1006324
rect 354916 1006312 354922 1006324
rect 360838 1006312 360844 1006324
rect 354916 1006284 360844 1006312
rect 354916 1006272 354922 1006284
rect 360838 1006272 360844 1006284
rect 360896 1006272 360902 1006324
rect 367370 1006272 367376 1006324
rect 367428 1006312 367434 1006324
rect 380158 1006312 380164 1006324
rect 367428 1006284 380164 1006312
rect 367428 1006272 367434 1006284
rect 380158 1006272 380164 1006284
rect 380216 1006272 380222 1006324
rect 423490 1006272 423496 1006324
rect 423548 1006312 423554 1006324
rect 429102 1006312 429108 1006324
rect 423548 1006284 429108 1006312
rect 423548 1006272 423554 1006284
rect 429102 1006272 429108 1006284
rect 429160 1006272 429166 1006324
rect 152090 1006176 152096 1006188
rect 151786 1006148 152096 1006176
rect 152090 1006136 152096 1006148
rect 152148 1006136 152154 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 161750 1006176 161756 1006188
rect 160336 1006148 161756 1006176
rect 160336 1006136 160342 1006148
rect 161750 1006136 161756 1006148
rect 161808 1006136 161814 1006188
rect 162302 1006136 162308 1006188
rect 162360 1006176 162366 1006188
rect 175918 1006176 175924 1006188
rect 162360 1006148 175924 1006176
rect 162360 1006136 162366 1006148
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 210418 1006136 210424 1006188
rect 210476 1006176 210482 1006188
rect 228358 1006176 228364 1006188
rect 210476 1006148 228364 1006176
rect 210476 1006136 210482 1006148
rect 228358 1006136 228364 1006148
rect 228416 1006136 228422 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 269758 1006176 269764 1006188
rect 262732 1006148 269764 1006176
rect 262732 1006136 262738 1006148
rect 269758 1006136 269764 1006148
rect 269816 1006136 269822 1006188
rect 298738 1006136 298744 1006188
rect 298796 1006176 298802 1006188
rect 304902 1006176 304908 1006188
rect 298796 1006148 304908 1006176
rect 298796 1006136 298802 1006148
rect 304902 1006136 304908 1006148
rect 304960 1006136 304966 1006188
rect 357710 1006136 357716 1006188
rect 357768 1006176 357774 1006188
rect 362218 1006176 362224 1006188
rect 357768 1006148 362224 1006176
rect 357768 1006136 357774 1006148
rect 362218 1006136 362224 1006148
rect 362276 1006136 362282 1006188
rect 365070 1006136 365076 1006188
rect 365128 1006176 365134 1006188
rect 367738 1006176 367744 1006188
rect 365128 1006148 367744 1006176
rect 365128 1006136 365134 1006148
rect 367738 1006136 367744 1006148
rect 367796 1006136 367802 1006188
rect 429396 1006176 429424 1006420
rect 553118 1006408 553124 1006460
rect 553176 1006448 553182 1006460
rect 553176 1006420 563054 1006448
rect 553176 1006408 553182 1006420
rect 431862 1006340 431868 1006392
rect 431920 1006380 431926 1006392
rect 431920 1006352 441614 1006380
rect 431920 1006340 431926 1006352
rect 412606 1006148 429424 1006176
rect 441586 1006176 441614 1006352
rect 505370 1006272 505376 1006324
rect 505428 1006312 505434 1006324
rect 505428 1006284 518894 1006312
rect 505428 1006272 505434 1006284
rect 469858 1006176 469864 1006188
rect 441586 1006148 469864 1006176
rect 102318 1006040 102324 1006052
rect 98472 1006012 102324 1006040
rect 102318 1006000 102324 1006012
rect 102376 1006000 102382 1006052
rect 108482 1006000 108488 1006052
rect 108540 1006040 108546 1006052
rect 126238 1006040 126244 1006052
rect 108540 1006012 126244 1006040
rect 108540 1006000 108546 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 148870 1006000 148876 1006052
rect 148928 1006040 148934 1006052
rect 150066 1006040 150072 1006052
rect 148928 1006012 150072 1006040
rect 148928 1006000 148934 1006012
rect 150066 1006000 150072 1006012
rect 150124 1006000 150130 1006052
rect 153930 1006000 153936 1006052
rect 153988 1006040 153994 1006052
rect 158254 1006040 158260 1006052
rect 153988 1006012 158260 1006040
rect 153988 1006000 153994 1006012
rect 158254 1006000 158260 1006012
rect 158312 1006000 158318 1006052
rect 159450 1006000 159456 1006052
rect 159508 1006040 159514 1006052
rect 177298 1006040 177304 1006052
rect 159508 1006012 177304 1006040
rect 159508 1006000 159514 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 198182 1006000 198188 1006052
rect 198240 1006040 198246 1006052
rect 201034 1006040 201040 1006052
rect 198240 1006012 201040 1006040
rect 198240 1006000 198246 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 208394 1006000 208400 1006052
rect 208452 1006040 208458 1006052
rect 229738 1006040 229744 1006052
rect 208452 1006012 229744 1006040
rect 208452 1006000 208458 1006012
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 249058 1006000 249064 1006052
rect 249116 1006040 249122 1006052
rect 257338 1006040 257344 1006052
rect 249116 1006012 257344 1006040
rect 249116 1006000 249122 1006012
rect 257338 1006000 257344 1006012
rect 257396 1006000 257402 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 279418 1006040 279424 1006052
rect 261904 1006012 279424 1006040
rect 261904 1006000 261910 1006012
rect 279418 1006000 279424 1006012
rect 279476 1006000 279482 1006052
rect 298922 1006000 298928 1006052
rect 298980 1006040 298986 1006052
rect 298980 1006012 303108 1006040
rect 298980 1006000 298986 1006012
rect 303080 1005904 303108 1006012
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 311802 1006040 311808 1006052
rect 304276 1006012 311808 1006040
rect 304276 1005904 304304 1006012
rect 311802 1006000 311808 1006012
rect 311860 1006000 311866 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 320818 1006040 320824 1006052
rect 314712 1006012 320824 1006040
rect 314712 1006000 314718 1006012
rect 320818 1006000 320824 1006012
rect 320876 1006000 320882 1006052
rect 355686 1006000 355692 1006052
rect 355744 1006040 355750 1006052
rect 359458 1006040 359464 1006052
rect 355744 1006012 359464 1006040
rect 355744 1006000 355750 1006012
rect 359458 1006000 359464 1006012
rect 359516 1006000 359522 1006052
rect 363414 1006000 363420 1006052
rect 363472 1006040 363478 1006052
rect 382918 1006040 382924 1006052
rect 363472 1006012 382924 1006040
rect 363472 1006000 363478 1006012
rect 382918 1006000 382924 1006012
rect 382976 1006000 382982 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 412606 1006040 412634 1006148
rect 469858 1006136 469864 1006148
rect 469916 1006136 469922 1006188
rect 507026 1006136 507032 1006188
rect 507084 1006176 507090 1006188
rect 509694 1006176 509700 1006188
rect 507084 1006148 509700 1006176
rect 507084 1006136 507090 1006148
rect 509694 1006136 509700 1006148
rect 509752 1006136 509758 1006188
rect 518866 1006176 518894 1006284
rect 552290 1006272 552296 1006324
rect 552348 1006312 552354 1006324
rect 558178 1006312 558184 1006324
rect 552348 1006284 558184 1006312
rect 552348 1006272 552354 1006284
rect 558178 1006272 558184 1006284
rect 558236 1006272 558242 1006324
rect 563026 1006312 563054 1006420
rect 570598 1006312 570604 1006324
rect 563026 1006284 570604 1006312
rect 570598 1006272 570604 1006284
rect 570656 1006272 570662 1006324
rect 519538 1006176 519544 1006188
rect 518866 1006148 519544 1006176
rect 519538 1006136 519544 1006148
rect 519596 1006136 519602 1006188
rect 551462 1006136 551468 1006188
rect 551520 1006176 551526 1006188
rect 557442 1006176 557448 1006188
rect 551520 1006148 557448 1006176
rect 551520 1006136 551526 1006148
rect 557442 1006136 557448 1006148
rect 557500 1006136 557506 1006188
rect 558822 1006136 558828 1006188
rect 558880 1006176 558886 1006188
rect 571978 1006176 571984 1006188
rect 558880 1006148 571984 1006176
rect 558880 1006136 558886 1006148
rect 571978 1006136 571984 1006148
rect 572036 1006136 572042 1006188
rect 400916 1006012 412634 1006040
rect 400916 1006000 400922 1006012
rect 423490 1006000 423496 1006052
rect 423548 1006040 423554 1006052
rect 430298 1006040 430304 1006052
rect 423548 1006012 430304 1006040
rect 423548 1006000 423554 1006012
rect 430298 1006000 430304 1006012
rect 430356 1006000 430362 1006052
rect 431678 1006000 431684 1006052
rect 431736 1006040 431742 1006052
rect 471238 1006040 471244 1006052
rect 431736 1006012 471244 1006040
rect 431736 1006000 431742 1006012
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 496722 1006000 496728 1006052
rect 496780 1006040 496786 1006052
rect 498838 1006040 498844 1006052
rect 496780 1006012 498844 1006040
rect 496780 1006000 496786 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 502518 1006000 502524 1006052
rect 502576 1006040 502582 1006052
rect 505738 1006040 505744 1006052
rect 502576 1006012 505744 1006040
rect 502576 1006000 502582 1006012
rect 505738 1006000 505744 1006012
rect 505796 1006000 505802 1006052
rect 506198 1006000 506204 1006052
rect 506256 1006040 506262 1006052
rect 506256 1006012 508912 1006040
rect 506256 1006000 506262 1006012
rect 303080 1005876 304304 1005904
rect 508884 1005904 508912 1006012
rect 509050 1006000 509056 1006052
rect 509108 1006040 509114 1006052
rect 509234 1006040 509240 1006052
rect 509108 1006012 509240 1006040
rect 509108 1006000 509114 1006012
rect 509234 1006000 509240 1006012
rect 509292 1006000 509298 1006052
rect 522298 1006040 522304 1006052
rect 509528 1006012 522304 1006040
rect 509528 1005904 509556 1006012
rect 522298 1006000 522304 1006012
rect 522356 1006000 522362 1006052
rect 555970 1006000 555976 1006052
rect 556028 1006040 556034 1006052
rect 573358 1006040 573364 1006052
rect 556028 1006012 573364 1006040
rect 556028 1006000 556034 1006012
rect 573358 1006000 573364 1006012
rect 573416 1006000 573422 1006052
rect 508884 1005876 509556 1005904
rect 429470 1005796 429476 1005848
rect 429528 1005836 429534 1005848
rect 429528 1005808 431724 1005836
rect 429528 1005796 429534 1005808
rect 426342 1005660 426348 1005712
rect 426400 1005700 426406 1005712
rect 431696 1005700 431724 1005808
rect 431862 1005796 431868 1005848
rect 431920 1005836 431926 1005848
rect 453298 1005836 453304 1005848
rect 431920 1005808 453304 1005836
rect 431920 1005796 431926 1005808
rect 453298 1005796 453304 1005808
rect 453356 1005796 453362 1005848
rect 509234 1005728 509240 1005780
rect 509292 1005768 509298 1005780
rect 514018 1005768 514024 1005780
rect 509292 1005740 514024 1005768
rect 509292 1005728 509298 1005740
rect 514018 1005728 514024 1005740
rect 514076 1005728 514082 1005780
rect 445018 1005700 445024 1005712
rect 426400 1005672 431632 1005700
rect 431696 1005672 445024 1005700
rect 426400 1005660 426406 1005672
rect 367002 1005524 367008 1005576
rect 367060 1005564 367066 1005576
rect 377398 1005564 377404 1005576
rect 367060 1005536 377404 1005564
rect 367060 1005524 367066 1005536
rect 377398 1005524 377404 1005536
rect 377456 1005524 377462 1005576
rect 425514 1005524 425520 1005576
rect 425572 1005564 425578 1005576
rect 431604 1005564 431632 1005672
rect 445018 1005660 445024 1005672
rect 445076 1005660 445082 1005712
rect 457438 1005564 457444 1005576
rect 425572 1005536 429700 1005564
rect 431604 1005536 457444 1005564
rect 425572 1005524 425578 1005536
rect 360562 1005388 360568 1005440
rect 360620 1005428 360626 1005440
rect 378778 1005428 378784 1005440
rect 360620 1005400 378784 1005428
rect 360620 1005388 360626 1005400
rect 378778 1005388 378784 1005400
rect 378836 1005388 378842 1005440
rect 424318 1005388 424324 1005440
rect 424376 1005428 424382 1005440
rect 429470 1005428 429476 1005440
rect 424376 1005400 429476 1005428
rect 424376 1005388 424382 1005400
rect 429470 1005388 429476 1005400
rect 429528 1005388 429534 1005440
rect 429672 1005428 429700 1005536
rect 457438 1005524 457444 1005536
rect 457496 1005524 457502 1005576
rect 462958 1005428 462964 1005440
rect 429672 1005400 462964 1005428
rect 462958 1005388 462964 1005400
rect 463016 1005388 463022 1005440
rect 552290 1005388 552296 1005440
rect 552348 1005428 552354 1005440
rect 566642 1005428 566648 1005440
rect 552348 1005400 566648 1005428
rect 552348 1005388 552354 1005400
rect 566642 1005388 566648 1005400
rect 566700 1005388 566706 1005440
rect 102778 1005252 102784 1005304
rect 102836 1005292 102842 1005304
rect 108850 1005292 108856 1005304
rect 102836 1005264 108856 1005292
rect 102836 1005252 102842 1005264
rect 108850 1005252 108856 1005264
rect 108908 1005252 108914 1005304
rect 204898 1005252 204904 1005304
rect 204956 1005292 204962 1005304
rect 212074 1005292 212080 1005304
rect 204956 1005264 212080 1005292
rect 204956 1005252 204962 1005264
rect 212074 1005252 212080 1005264
rect 212132 1005252 212138 1005304
rect 356514 1005252 356520 1005304
rect 356572 1005292 356578 1005304
rect 373258 1005292 373264 1005304
rect 356572 1005264 373264 1005292
rect 356572 1005252 356578 1005264
rect 373258 1005252 373264 1005264
rect 373316 1005252 373322 1005304
rect 425146 1005252 425152 1005304
rect 425204 1005292 425210 1005304
rect 468478 1005292 468484 1005304
rect 425204 1005264 468484 1005292
rect 425204 1005252 425210 1005264
rect 468478 1005252 468484 1005264
rect 468536 1005252 468542 1005304
rect 498838 1005252 498844 1005304
rect 498896 1005292 498902 1005304
rect 516778 1005292 516784 1005304
rect 498896 1005264 516784 1005292
rect 498896 1005252 498902 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 551462 1005252 551468 1005304
rect 551520 1005292 551526 1005304
rect 569218 1005292 569224 1005304
rect 551520 1005264 569224 1005292
rect 551520 1005252 551526 1005264
rect 569218 1005252 569224 1005264
rect 569276 1005252 569282 1005304
rect 304258 1005184 304264 1005236
rect 304316 1005224 304322 1005236
rect 307294 1005224 307300 1005236
rect 304316 1005196 307300 1005224
rect 304316 1005184 304322 1005196
rect 307294 1005184 307300 1005196
rect 307352 1005184 307358 1005236
rect 429102 1005116 429108 1005168
rect 429160 1005156 429166 1005168
rect 447778 1005156 447784 1005168
rect 429160 1005128 447784 1005156
rect 429160 1005116 429166 1005128
rect 447778 1005116 447784 1005128
rect 447836 1005116 447842 1005168
rect 149882 1005048 149888 1005100
rect 149940 1005088 149946 1005100
rect 152918 1005088 152924 1005100
rect 149940 1005060 152924 1005088
rect 149940 1005048 149946 1005060
rect 152918 1005048 152924 1005060
rect 152976 1005048 152982 1005100
rect 305822 1005048 305828 1005100
rect 305880 1005088 305886 1005100
rect 308950 1005088 308956 1005100
rect 305880 1005060 308956 1005088
rect 305880 1005048 305886 1005060
rect 308950 1005048 308956 1005060
rect 309008 1005048 309014 1005100
rect 365070 1005048 365076 1005100
rect 365128 1005088 365134 1005100
rect 370498 1005088 370504 1005100
rect 365128 1005060 370504 1005088
rect 365128 1005048 365134 1005060
rect 370498 1005048 370504 1005060
rect 370556 1005048 370562 1005100
rect 508222 1005048 508228 1005100
rect 508280 1005088 508286 1005100
rect 511258 1005088 511264 1005100
rect 508280 1005060 511264 1005088
rect 508280 1005048 508286 1005060
rect 511258 1005048 511264 1005060
rect 511316 1005048 511322 1005100
rect 427998 1004980 428004 1005032
rect 428056 1005020 428062 1005032
rect 431862 1005020 431868 1005032
rect 428056 1004992 431868 1005020
rect 428056 1004980 428062 1004992
rect 431862 1004980 431868 1004992
rect 431920 1004980 431926 1005032
rect 151078 1004912 151084 1004964
rect 151136 1004952 151142 1004964
rect 153746 1004952 153752 1004964
rect 151136 1004924 153752 1004952
rect 151136 1004912 151142 1004924
rect 153746 1004912 153752 1004924
rect 153804 1004912 153810 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 263042 1004912 263048 1004964
rect 263100 1004952 263106 1004964
rect 268378 1004952 268384 1004964
rect 263100 1004924 268384 1004952
rect 263100 1004912 263106 1004924
rect 268378 1004912 268384 1004924
rect 268436 1004912 268442 1004964
rect 353202 1004912 353208 1004964
rect 353260 1004952 353266 1004964
rect 355686 1004952 355692 1004964
rect 353260 1004924 355692 1004952
rect 353260 1004912 353266 1004924
rect 355686 1004912 355692 1004924
rect 355744 1004912 355750 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 364978 1004952 364984 1004964
rect 361448 1004924 364984 1004952
rect 361448 1004912 361454 1004924
rect 364978 1004912 364984 1004924
rect 365036 1004912 365042 1004964
rect 497918 1004912 497924 1004964
rect 497976 1004952 497982 1004964
rect 500494 1004952 500500 1004964
rect 497976 1004924 500500 1004952
rect 497976 1004912 497982 1004924
rect 500494 1004912 500500 1004924
rect 500552 1004912 500558 1004964
rect 149698 1004776 149704 1004828
rect 149756 1004816 149762 1004828
rect 151722 1004816 151728 1004828
rect 149756 1004788 151728 1004816
rect 149756 1004776 149762 1004788
rect 151722 1004776 151728 1004788
rect 151780 1004776 151786 1004828
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 211246 1004776 211252 1004828
rect 211304 1004816 211310 1004828
rect 215938 1004816 215944 1004828
rect 211304 1004788 215944 1004816
rect 211304 1004776 211310 1004788
rect 215938 1004776 215944 1004788
rect 215996 1004776 216002 1004828
rect 258166 1004776 258172 1004828
rect 258224 1004816 258230 1004828
rect 259454 1004816 259460 1004828
rect 258224 1004788 259460 1004816
rect 258224 1004776 258230 1004788
rect 259454 1004776 259460 1004788
rect 259512 1004776 259518 1004828
rect 305638 1004776 305644 1004828
rect 305696 1004816 305702 1004828
rect 308122 1004816 308128 1004828
rect 305696 1004788 308128 1004816
rect 305696 1004776 305702 1004788
rect 308122 1004776 308128 1004788
rect 308180 1004776 308186 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 354582 1004776 354588 1004828
rect 354640 1004816 354646 1004828
rect 356514 1004816 356520 1004828
rect 354640 1004788 356520 1004816
rect 354640 1004776 354646 1004788
rect 356514 1004776 356520 1004788
rect 356572 1004776 356578 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365162 1004816 365168 1004828
rect 362644 1004788 365168 1004816
rect 362644 1004776 362650 1004788
rect 365162 1004776 365168 1004788
rect 365220 1004776 365226 1004828
rect 420822 1004776 420828 1004828
rect 420880 1004816 420886 1004828
rect 422662 1004816 422668 1004828
rect 420880 1004788 422668 1004816
rect 420880 1004776 420886 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 498102 1004776 498108 1004828
rect 498160 1004816 498166 1004828
rect 499666 1004816 499672 1004828
rect 498160 1004788 499672 1004816
rect 498160 1004776 498166 1004788
rect 499666 1004776 499672 1004788
rect 499724 1004776 499730 1004828
rect 508222 1004776 508228 1004828
rect 508280 1004816 508286 1004828
rect 510798 1004816 510804 1004828
rect 508280 1004788 510804 1004816
rect 508280 1004776 508286 1004788
rect 510798 1004776 510804 1004788
rect 510856 1004776 510862 1004828
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 151262 1004640 151268 1004692
rect 151320 1004680 151326 1004692
rect 154114 1004680 154120 1004692
rect 151320 1004652 154120 1004680
rect 151320 1004640 151326 1004652
rect 154114 1004640 154120 1004652
rect 154172 1004640 154178 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 304902 1004640 304908 1004692
rect 304960 1004680 304966 1004692
rect 306926 1004680 306932 1004692
rect 304960 1004652 306932 1004680
rect 304960 1004640 304966 1004652
rect 306926 1004640 306932 1004652
rect 306984 1004640 306990 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 432874 1004640 432880 1004692
rect 432932 1004680 432938 1004692
rect 438118 1004680 438124 1004692
rect 432932 1004652 438124 1004680
rect 432932 1004640 432938 1004652
rect 438118 1004640 438124 1004652
rect 438176 1004640 438182 1004692
rect 499482 1004640 499488 1004692
rect 499540 1004680 499546 1004692
rect 500494 1004680 500500 1004692
rect 499540 1004652 500500 1004680
rect 499540 1004640 499546 1004652
rect 500494 1004640 500500 1004652
rect 500552 1004640 500558 1004692
rect 507394 1004640 507400 1004692
rect 507452 1004680 507458 1004692
rect 509234 1004680 509240 1004692
rect 507452 1004652 509240 1004680
rect 507452 1004640 507458 1004652
rect 509234 1004640 509240 1004652
rect 509292 1004640 509298 1004692
rect 560846 1004640 560852 1004692
rect 560904 1004680 560910 1004692
rect 566458 1004680 566464 1004692
rect 560904 1004652 566464 1004680
rect 560904 1004640 560910 1004652
rect 566458 1004640 566464 1004652
rect 566516 1004640 566522 1004692
rect 504542 1004368 504548 1004420
rect 504600 1004408 504606 1004420
rect 510982 1004408 510988 1004420
rect 504600 1004380 510988 1004408
rect 504600 1004368 504606 1004380
rect 510982 1004368 510988 1004380
rect 511040 1004368 511046 1004420
rect 426342 1004028 426348 1004080
rect 426400 1004068 426406 1004080
rect 455874 1004068 455880 1004080
rect 426400 1004040 455880 1004068
rect 426400 1004028 426406 1004040
rect 455874 1004028 455880 1004040
rect 455932 1004028 455938 1004080
rect 92290 1003892 92296 1003944
rect 92348 1003932 92354 1003944
rect 103146 1003932 103152 1003944
rect 92348 1003904 103152 1003932
rect 92348 1003892 92354 1003904
rect 103146 1003892 103152 1003904
rect 103204 1003892 103210 1003944
rect 247310 1003892 247316 1003944
rect 247368 1003932 247374 1003944
rect 255314 1003932 255320 1003944
rect 247368 1003904 255320 1003932
rect 247368 1003892 247374 1003904
rect 255314 1003892 255320 1003904
rect 255372 1003892 255378 1003944
rect 421834 1003892 421840 1003944
rect 421892 1003932 421898 1003944
rect 464338 1003932 464344 1003944
rect 421892 1003904 464344 1003932
rect 421892 1003892 421898 1003904
rect 464338 1003892 464344 1003904
rect 464396 1003892 464402 1003944
rect 557166 1003892 557172 1003944
rect 557224 1003932 557230 1003944
rect 571242 1003932 571248 1003944
rect 557224 1003904 571248 1003932
rect 557224 1003892 557230 1003904
rect 571242 1003892 571248 1003904
rect 571300 1003892 571306 1003944
rect 300302 1003280 300308 1003332
rect 300360 1003320 300366 1003332
rect 305270 1003320 305276 1003332
rect 300360 1003292 305276 1003320
rect 300360 1003280 300366 1003292
rect 305270 1003280 305276 1003292
rect 305328 1003280 305334 1003332
rect 501690 1003280 501696 1003332
rect 501748 1003320 501754 1003332
rect 504726 1003320 504732 1003332
rect 501748 1003292 504732 1003320
rect 501748 1003280 501754 1003292
rect 504726 1003280 504732 1003292
rect 504784 1003280 504790 1003332
rect 371234 1002940 371240 1002992
rect 371292 1002980 371298 1002992
rect 374362 1002980 374368 1002992
rect 371292 1002952 374368 1002980
rect 371292 1002940 371298 1002952
rect 374362 1002940 374368 1002952
rect 374420 1002940 374426 1002992
rect 253106 1002668 253112 1002720
rect 253164 1002708 253170 1002720
rect 256142 1002708 256148 1002720
rect 253164 1002680 256148 1002708
rect 253164 1002668 253170 1002680
rect 256142 1002668 256148 1002680
rect 256200 1002668 256206 1002720
rect 98638 1002600 98644 1002652
rect 98696 1002640 98702 1002652
rect 101950 1002640 101956 1002652
rect 98696 1002612 101956 1002640
rect 98696 1002600 98702 1002612
rect 101950 1002600 101956 1002612
rect 102008 1002600 102014 1002652
rect 302234 1002600 302240 1002652
rect 302292 1002640 302298 1002652
rect 304902 1002640 304908 1002652
rect 302292 1002612 304908 1002640
rect 302292 1002600 302298 1002612
rect 304902 1002600 304908 1002612
rect 304960 1002600 304966 1002652
rect 246574 1002532 246580 1002584
rect 246632 1002572 246638 1002584
rect 254118 1002572 254124 1002584
rect 246632 1002544 254124 1002572
rect 246632 1002532 246638 1002544
rect 254118 1002532 254124 1002544
rect 254176 1002532 254182 1002584
rect 440234 1002532 440240 1002584
rect 440292 1002572 440298 1002584
rect 466362 1002572 466368 1002584
rect 440292 1002544 466368 1002572
rect 440292 1002532 440298 1002544
rect 466362 1002532 466368 1002544
rect 466420 1002532 466426 1002584
rect 97442 1002464 97448 1002516
rect 97500 1002504 97506 1002516
rect 100294 1002504 100300 1002516
rect 97500 1002476 100300 1002504
rect 97500 1002464 97506 1002476
rect 100294 1002464 100300 1002476
rect 100352 1002464 100358 1002516
rect 261018 1002464 261024 1002516
rect 261076 1002504 261082 1002516
rect 264238 1002504 264244 1002516
rect 261076 1002476 264244 1002504
rect 261076 1002464 261082 1002476
rect 264238 1002464 264244 1002476
rect 264296 1002464 264302 1002516
rect 560846 1002464 560852 1002516
rect 560904 1002504 560910 1002516
rect 565078 1002504 565084 1002516
rect 560904 1002476 565084 1002504
rect 560904 1002464 560910 1002476
rect 565078 1002464 565084 1002476
rect 565136 1002464 565142 1002516
rect 96062 1002328 96068 1002380
rect 96120 1002368 96126 1002380
rect 99098 1002368 99104 1002380
rect 96120 1002340 99104 1002368
rect 96120 1002328 96126 1002340
rect 99098 1002328 99104 1002340
rect 99156 1002328 99162 1002380
rect 107654 1002328 107660 1002380
rect 107712 1002368 107718 1002380
rect 109494 1002368 109500 1002380
rect 107712 1002340 109500 1002368
rect 107712 1002328 107718 1002340
rect 109494 1002328 109500 1002340
rect 109552 1002328 109558 1002380
rect 148502 1002328 148508 1002380
rect 148560 1002368 148566 1002380
rect 150894 1002368 150900 1002380
rect 148560 1002340 150900 1002368
rect 148560 1002328 148566 1002340
rect 150894 1002328 150900 1002340
rect 150952 1002328 150958 1002380
rect 251818 1002328 251824 1002380
rect 251876 1002368 251882 1002380
rect 254486 1002368 254492 1002380
rect 251876 1002340 254492 1002368
rect 251876 1002328 251882 1002340
rect 254486 1002328 254492 1002340
rect 254544 1002328 254550 1002380
rect 260190 1002328 260196 1002380
rect 260248 1002368 260254 1002380
rect 262858 1002368 262864 1002380
rect 260248 1002340 262864 1002368
rect 260248 1002328 260254 1002340
rect 262858 1002328 262864 1002340
rect 262916 1002328 262922 1002380
rect 503346 1002328 503352 1002380
rect 503404 1002368 503410 1002380
rect 506474 1002368 506480 1002380
rect 503404 1002340 506480 1002368
rect 503404 1002328 503410 1002340
rect 506474 1002328 506480 1002340
rect 506532 1002328 506538 1002380
rect 551922 1002328 551928 1002380
rect 551980 1002368 551986 1002380
rect 553946 1002368 553952 1002380
rect 551980 1002340 553952 1002368
rect 551980 1002328 551986 1002340
rect 553946 1002328 553952 1002340
rect 554004 1002328 554010 1002380
rect 560478 1002328 560484 1002380
rect 560536 1002368 560542 1002380
rect 563054 1002368 563060 1002380
rect 560536 1002340 563060 1002368
rect 560536 1002328 560542 1002340
rect 563054 1002328 563060 1002340
rect 563112 1002328 563118 1002380
rect 98822 1002192 98828 1002244
rect 98880 1002232 98886 1002244
rect 101122 1002232 101128 1002244
rect 98880 1002204 101128 1002232
rect 98880 1002192 98886 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 105630 1002192 105636 1002244
rect 105688 1002232 105694 1002244
rect 107838 1002232 107844 1002244
rect 105688 1002204 107844 1002232
rect 105688 1002192 105694 1002204
rect 107838 1002192 107844 1002204
rect 107896 1002192 107902 1002244
rect 108022 1002192 108028 1002244
rect 108080 1002232 108086 1002244
rect 110414 1002232 110420 1002244
rect 108080 1002204 110420 1002232
rect 108080 1002192 108086 1002204
rect 110414 1002192 110420 1002204
rect 110472 1002192 110478 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 157334 1002232 157340 1002244
rect 155828 1002204 157340 1002232
rect 155828 1002192 155834 1002204
rect 157334 1002192 157340 1002204
rect 157392 1002192 157398 1002244
rect 203334 1002192 203340 1002244
rect 203392 1002232 203398 1002244
rect 206370 1002232 206376 1002244
rect 203392 1002204 206376 1002232
rect 203392 1002192 203398 1002204
rect 206370 1002192 206376 1002204
rect 206428 1002192 206434 1002244
rect 206738 1002192 206744 1002244
rect 206796 1002232 206802 1002244
rect 208578 1002232 208584 1002244
rect 206796 1002204 208584 1002232
rect 206796 1002192 206802 1002204
rect 208578 1002192 208584 1002204
rect 208636 1002192 208642 1002244
rect 254578 1002192 254584 1002244
rect 254636 1002232 254642 1002244
rect 256510 1002232 256516 1002244
rect 254636 1002204 256516 1002232
rect 254636 1002192 254642 1002204
rect 256510 1002192 256516 1002204
rect 256568 1002192 256574 1002244
rect 259822 1002192 259828 1002244
rect 259880 1002232 259886 1002244
rect 262214 1002232 262220 1002244
rect 259880 1002204 262220 1002232
rect 259880 1002192 259886 1002204
rect 262214 1002192 262220 1002204
rect 262272 1002192 262278 1002244
rect 303246 1002192 303252 1002244
rect 303304 1002232 303310 1002244
rect 306098 1002232 306104 1002244
rect 303304 1002204 306104 1002232
rect 303304 1002192 303310 1002204
rect 306098 1002192 306104 1002204
rect 306156 1002192 306162 1002244
rect 308398 1002192 308404 1002244
rect 308456 1002232 308462 1002244
rect 310606 1002232 310612 1002244
rect 308456 1002204 310612 1002232
rect 308456 1002192 308462 1002204
rect 310606 1002192 310612 1002204
rect 310664 1002192 310670 1002244
rect 355318 1002192 355324 1002244
rect 355376 1002232 355382 1002244
rect 358538 1002232 358544 1002244
rect 355376 1002204 358544 1002232
rect 355376 1002192 355382 1002204
rect 358538 1002192 358544 1002204
rect 358596 1002192 358602 1002244
rect 553302 1002192 553308 1002244
rect 553360 1002232 553366 1002244
rect 555142 1002232 555148 1002244
rect 553360 1002204 555148 1002232
rect 553360 1002192 553366 1002204
rect 555142 1002192 555148 1002204
rect 555200 1002192 555206 1002244
rect 97258 1002056 97264 1002108
rect 97316 1002096 97322 1002108
rect 99466 1002096 99472 1002108
rect 97316 1002068 99472 1002096
rect 97316 1002056 97322 1002068
rect 99466 1002056 99472 1002068
rect 99524 1002056 99530 1002108
rect 100018 1002056 100024 1002108
rect 100076 1002096 100082 1002108
rect 103146 1002096 103152 1002108
rect 100076 1002068 103152 1002096
rect 100076 1002056 100082 1002068
rect 103146 1002056 103152 1002068
rect 103204 1002056 103210 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111794 1002096 111800 1002108
rect 109736 1002068 111800 1002096
rect 109736 1002056 109742 1002068
rect 111794 1002056 111800 1002068
rect 111852 1002056 111858 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 152458 1002056 152464 1002108
rect 152516 1002096 152522 1002108
rect 154574 1002096 154580 1002108
rect 152516 1002068 154580 1002096
rect 152516 1002056 152522 1002068
rect 154574 1002056 154580 1002068
rect 154632 1002056 154638 1002108
rect 157794 1002056 157800 1002108
rect 157852 1002096 157858 1002108
rect 160094 1002096 160100 1002108
rect 157852 1002068 160100 1002096
rect 157852 1002056 157858 1002068
rect 160094 1002056 160100 1002068
rect 160152 1002056 160158 1002108
rect 205082 1002056 205088 1002108
rect 205140 1002096 205146 1002108
rect 207198 1002096 207204 1002108
rect 205140 1002068 207204 1002096
rect 205140 1002056 205146 1002068
rect 207198 1002056 207204 1002068
rect 207256 1002056 207262 1002108
rect 210878 1002056 210884 1002108
rect 210936 1002096 210942 1002108
rect 213178 1002096 213184 1002108
rect 210936 1002068 213184 1002096
rect 210936 1002056 210942 1002068
rect 213178 1002056 213184 1002068
rect 213236 1002056 213242 1002108
rect 253382 1002056 253388 1002108
rect 253440 1002096 253446 1002108
rect 255314 1002096 255320 1002108
rect 253440 1002068 255320 1002096
rect 253440 1002056 253446 1002068
rect 255314 1002056 255320 1002068
rect 255372 1002056 255378 1002108
rect 261018 1002056 261024 1002108
rect 261076 1002096 261082 1002108
rect 261076 1002068 263364 1002096
rect 261076 1002056 261082 1002068
rect 95878 1001920 95884 1001972
rect 95936 1001960 95942 1001972
rect 98270 1001960 98276 1001972
rect 95936 1001932 98276 1001960
rect 95936 1001920 95942 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 99006 1001920 99012 1001972
rect 99064 1001960 99070 1001972
rect 101122 1001960 101128 1001972
rect 99064 1001932 101128 1001960
rect 99064 1001920 99070 1001932
rect 101122 1001920 101128 1001932
rect 101180 1001920 101186 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 107746 1001960 107752 1001972
rect 106056 1001932 107752 1001960
rect 106056 1001920 106062 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 156598 1001920 156604 1001972
rect 156656 1001960 156662 1001972
rect 158714 1001960 158720 1001972
rect 156656 1001932 158720 1001960
rect 156656 1001920 156662 1001932
rect 158714 1001920 158720 1001932
rect 158772 1001920 158778 1001972
rect 195146 1001920 195152 1001972
rect 195204 1001960 195210 1001972
rect 202690 1001960 202696 1001972
rect 195204 1001932 202696 1001960
rect 195204 1001920 195210 1001932
rect 202690 1001920 202696 1001932
rect 202748 1001920 202754 1001972
rect 203702 1001920 203708 1001972
rect 203760 1001960 203766 1001972
rect 205542 1001960 205548 1001972
rect 203760 1001932 205548 1001960
rect 203760 1001920 203766 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 212534 1001920 212540 1001972
rect 212592 1001960 212598 1001972
rect 214558 1001960 214564 1001972
rect 212592 1001932 214564 1001960
rect 212592 1001920 212598 1001932
rect 214558 1001920 214564 1001932
rect 214616 1001920 214622 1001972
rect 254762 1001920 254768 1001972
rect 254820 1001960 254826 1001972
rect 256970 1001960 256976 1001972
rect 254820 1001932 256976 1001960
rect 254820 1001920 254826 1001932
rect 256970 1001920 256976 1001932
rect 257028 1001920 257034 1001972
rect 260190 1001920 260196 1001972
rect 260248 1001960 260254 1001972
rect 260926 1001960 260932 1001972
rect 260248 1001932 260932 1001960
rect 260248 1001920 260254 1001932
rect 260926 1001920 260932 1001932
rect 260984 1001920 260990 1001972
rect 263336 1001960 263364 1002068
rect 263502 1002056 263508 1002108
rect 263560 1002096 263566 1002108
rect 265618 1002096 265624 1002108
rect 263560 1002068 265624 1002096
rect 263560 1002056 263566 1002068
rect 265618 1002056 265624 1002068
rect 265676 1002056 265682 1002108
rect 300118 1002056 300124 1002108
rect 300176 1002096 300182 1002108
rect 304074 1002096 304080 1002108
rect 300176 1002068 304080 1002096
rect 300176 1002056 300182 1002068
rect 304074 1002056 304080 1002068
rect 304132 1002056 304138 1002108
rect 355778 1002056 355784 1002108
rect 355836 1002096 355842 1002108
rect 357710 1002096 357716 1002108
rect 355836 1002068 357716 1002096
rect 355836 1002056 355842 1002068
rect 357710 1002056 357716 1002068
rect 357768 1002056 357774 1002108
rect 503346 1002056 503352 1002108
rect 503404 1002096 503410 1002108
rect 506290 1002096 506296 1002108
rect 503404 1002068 506296 1002096
rect 503404 1002056 503410 1002068
rect 506290 1002056 506296 1002068
rect 506348 1002056 506354 1002108
rect 509878 1002056 509884 1002108
rect 509936 1002096 509942 1002108
rect 515398 1002096 515404 1002108
rect 509936 1002068 515404 1002096
rect 509936 1002056 509942 1002068
rect 515398 1002056 515404 1002068
rect 515456 1002056 515462 1002108
rect 427538 1001988 427544 1002040
rect 427596 1002028 427602 1002040
rect 431862 1002028 431868 1002040
rect 427596 1002000 431868 1002028
rect 427596 1001988 427602 1002000
rect 431862 1001988 431868 1002000
rect 431920 1001988 431926 1002040
rect 263594 1001960 263600 1001972
rect 263336 1001932 263600 1001960
rect 263594 1001920 263600 1001932
rect 263652 1001920 263658 1001972
rect 263870 1001920 263876 1001972
rect 263928 1001960 263934 1001972
rect 266998 1001960 267004 1001972
rect 263928 1001932 267004 1001960
rect 263928 1001920 263934 1001932
rect 266998 1001920 267004 1001932
rect 267056 1001920 267062 1001972
rect 302878 1001920 302884 1001972
rect 302936 1001960 302942 1001972
rect 306098 1001960 306104 1001972
rect 302936 1001932 306104 1001960
rect 302936 1001920 302942 1001932
rect 306098 1001920 306104 1001932
rect 306156 1001920 306162 1001972
rect 307018 1001920 307024 1001972
rect 307076 1001960 307082 1001972
rect 308950 1001960 308956 1001972
rect 307076 1001932 308956 1001960
rect 307076 1001920 307082 1001932
rect 308950 1001920 308956 1001932
rect 309008 1001920 309014 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 360194 1001920 360200 1001972
rect 360252 1001960 360258 1001972
rect 363598 1001960 363604 1001972
rect 360252 1001932 363604 1001960
rect 360252 1001920 360258 1001932
rect 363598 1001920 363604 1001932
rect 363656 1001920 363662 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 423582 1001920 423588 1001972
rect 423640 1001960 423646 1001972
rect 424318 1001960 424324 1001972
rect 423640 1001932 424324 1001960
rect 423640 1001920 423646 1001932
rect 424318 1001920 424324 1001932
rect 424376 1001920 424382 1001972
rect 500862 1001920 500868 1001972
rect 500920 1001960 500926 1001972
rect 501690 1001960 501696 1001972
rect 500920 1001932 501696 1001960
rect 500920 1001920 500926 1001932
rect 501690 1001920 501696 1001932
rect 501748 1001920 501754 1001972
rect 502150 1001920 502156 1001972
rect 502208 1001960 502214 1001972
rect 504174 1001960 504180 1001972
rect 502208 1001932 504180 1001960
rect 502208 1001920 502214 1001932
rect 504174 1001920 504180 1001932
rect 504232 1001920 504238 1001972
rect 505370 1001920 505376 1001972
rect 505428 1001960 505434 1001972
rect 508498 1001960 508504 1001972
rect 505428 1001932 508504 1001960
rect 505428 1001920 505434 1001932
rect 508498 1001920 508504 1001932
rect 508556 1001920 508562 1001972
rect 510338 1001920 510344 1001972
rect 510396 1001960 510402 1001972
rect 512638 1001960 512644 1001972
rect 510396 1001932 512644 1001960
rect 510396 1001920 510402 1001932
rect 512638 1001920 512644 1001932
rect 512696 1001920 512702 1001972
rect 552658 1001920 552664 1001972
rect 552716 1001960 552722 1001972
rect 554314 1001960 554320 1001972
rect 552716 1001932 554320 1001960
rect 552716 1001920 552722 1001932
rect 554314 1001920 554320 1001932
rect 554372 1001920 554378 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 563698 1001960 563704 1001972
rect 561732 1001932 563704 1001960
rect 561732 1001920 561738 1001932
rect 563698 1001920 563704 1001932
rect 563756 1001920 563762 1001972
rect 551094 1001308 551100 1001360
rect 551152 1001348 551158 1001360
rect 568482 1001348 568488 1001360
rect 551152 1001320 568488 1001348
rect 551152 1001308 551158 1001320
rect 568482 1001308 568488 1001320
rect 568540 1001308 568546 1001360
rect 195514 1001172 195520 1001224
rect 195572 1001212 195578 1001224
rect 203886 1001212 203892 1001224
rect 195572 1001184 203892 1001212
rect 195572 1001172 195578 1001184
rect 203886 1001172 203892 1001184
rect 203944 1001172 203950 1001224
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 423582 1001172 423588 1001224
rect 423640 1001212 423646 1001224
rect 440234 1001212 440240 1001224
rect 423640 1001184 440240 1001212
rect 423640 1001172 423646 1001184
rect 440234 1001172 440240 1001184
rect 440292 1001172 440298 1001224
rect 498102 1001172 498108 1001224
rect 498160 1001212 498166 1001224
rect 521286 1001212 521292 1001224
rect 498160 1001184 521292 1001212
rect 498160 1001172 498166 1001184
rect 521286 1001172 521292 1001184
rect 521344 1001172 521350 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 298278 1000492 298284 1000544
rect 298336 1000532 298342 1000544
rect 305822 1000532 305828 1000544
rect 298336 1000504 305828 1000532
rect 298336 1000492 298342 1000504
rect 305822 1000492 305828 1000504
rect 305880 1000492 305886 1000544
rect 427170 1000492 427176 1000544
rect 427228 1000532 427234 1000544
rect 430482 1000532 430488 1000544
rect 427228 1000504 430488 1000532
rect 427228 1000492 427234 1000504
rect 430482 1000492 430488 1000504
rect 430540 1000492 430546 1000544
rect 247126 999744 247132 999796
rect 247184 999784 247190 999796
rect 254762 999784 254768 999796
rect 247184 999756 254768 999784
rect 247184 999744 247190 999756
rect 254762 999744 254768 999756
rect 254820 999744 254826 999796
rect 430298 999744 430304 999796
rect 430356 999784 430362 999796
rect 443638 999784 443644 999796
rect 430356 999756 443644 999784
rect 430356 999744 430362 999756
rect 443638 999744 443644 999756
rect 443696 999744 443702 999796
rect 514754 999268 514760 999320
rect 514812 999308 514818 999320
rect 514812 999280 518894 999308
rect 514812 999268 514818 999280
rect 95142 999132 95148 999184
rect 95200 999172 95206 999184
rect 99006 999172 99012 999184
rect 95200 999144 99012 999172
rect 95200 999132 95206 999144
rect 99006 999132 99012 999144
rect 99064 999132 99070 999184
rect 506474 999132 506480 999184
rect 506532 999172 506538 999184
rect 517422 999172 517428 999184
rect 506532 999144 517428 999172
rect 506532 999132 506538 999144
rect 517422 999132 517428 999144
rect 517480 999132 517486 999184
rect 518866 999104 518894 999280
rect 555142 999132 555148 999184
rect 555200 999172 555206 999184
rect 556154 999172 556160 999184
rect 555200 999144 556160 999172
rect 555200 999132 555206 999144
rect 556154 999132 556160 999144
rect 556212 999132 556218 999184
rect 618162 999132 618168 999184
rect 618220 999172 618226 999184
rect 625246 999172 625252 999184
rect 618220 999144 625252 999172
rect 618220 999132 618226 999144
rect 625246 999132 625252 999144
rect 625304 999132 625310 999184
rect 523494 999104 523500 999116
rect 518866 999076 523500 999104
rect 523494 999064 523500 999076
rect 523552 999064 523558 999116
rect 457438 998928 457444 998980
rect 457496 998968 457502 998980
rect 472618 998968 472624 998980
rect 457496 998940 472624 998968
rect 457496 998928 457502 998940
rect 472618 998928 472624 998940
rect 472676 998928 472682 998980
rect 504726 998928 504732 998980
rect 504784 998968 504790 998980
rect 517698 998968 517704 998980
rect 504784 998940 517704 998968
rect 504784 998928 504790 998940
rect 517698 998928 517704 998940
rect 517756 998928 517762 998980
rect 92290 998792 92296 998844
rect 92348 998832 92354 998844
rect 92934 998832 92940 998844
rect 92348 998804 92940 998832
rect 92348 998792 92354 998804
rect 92934 998792 92940 998804
rect 92992 998792 92998 998844
rect 428366 998792 428372 998844
rect 428424 998832 428430 998844
rect 436094 998832 436100 998844
rect 428424 998804 436100 998832
rect 428424 998792 428430 998804
rect 436094 998792 436100 998804
rect 436152 998792 436158 998844
rect 453298 998792 453304 998844
rect 453356 998832 453362 998844
rect 472434 998832 472440 998844
rect 453356 998804 472440 998832
rect 453356 998792 453362 998804
rect 472434 998792 472440 998804
rect 472492 998792 472498 998844
rect 517238 998792 517244 998844
rect 517296 998832 517302 998844
rect 522114 998832 522120 998844
rect 517296 998804 522120 998832
rect 517296 998792 517302 998804
rect 522114 998792 522120 998804
rect 522172 998792 522178 998844
rect 383286 998764 383292 998776
rect 373966 998736 383292 998764
rect 196802 998656 196808 998708
rect 196860 998696 196866 998708
rect 204346 998696 204352 998708
rect 196860 998668 204352 998696
rect 196860 998656 196866 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 357434 998656 357440 998708
rect 357492 998696 357498 998708
rect 373966 998696 373994 998736
rect 383286 998724 383292 998736
rect 383344 998724 383350 998776
rect 502150 998724 502156 998776
rect 502208 998764 502214 998776
rect 516870 998764 516876 998776
rect 502208 998736 516876 998764
rect 502208 998724 502214 998736
rect 516870 998724 516876 998736
rect 516928 998724 516934 998776
rect 357492 998668 373994 998696
rect 357492 998656 357498 998668
rect 430482 998656 430488 998708
rect 430540 998696 430546 998708
rect 456794 998696 456800 998708
rect 430540 998668 456800 998696
rect 430540 998656 430546 998668
rect 456794 998656 456800 998668
rect 456852 998656 456858 998708
rect 467098 998656 467104 998708
rect 467156 998696 467162 998708
rect 471974 998696 471980 998708
rect 467156 998668 471980 998696
rect 467156 998656 467162 998668
rect 471974 998656 471980 998668
rect 472032 998656 472038 998708
rect 517422 998656 517428 998708
rect 517480 998696 517486 998708
rect 523678 998696 523684 998708
rect 517480 998668 523684 998696
rect 517480 998656 517486 998668
rect 523678 998656 523684 998668
rect 523736 998656 523742 998708
rect 378778 998588 378784 998640
rect 378836 998628 378842 998640
rect 383562 998628 383568 998640
rect 378836 998600 383568 998628
rect 378836 998588 378842 998600
rect 383562 998588 383568 998600
rect 383620 998588 383626 998640
rect 196618 998520 196624 998572
rect 196676 998560 196682 998572
rect 203518 998560 203524 998572
rect 196676 998532 203524 998560
rect 196676 998520 196682 998532
rect 203518 998520 203524 998532
rect 203576 998520 203582 998572
rect 351822 998520 351828 998572
rect 351880 998560 351886 998572
rect 378594 998560 378600 998572
rect 351880 998532 378600 998560
rect 351880 998520 351886 998532
rect 378594 998520 378600 998532
rect 378652 998520 378658 998572
rect 430850 998520 430856 998572
rect 430908 998560 430914 998572
rect 433978 998560 433984 998572
rect 430908 998532 433984 998560
rect 430908 998520 430914 998532
rect 433978 998520 433984 998532
rect 434036 998520 434042 998572
rect 436094 998520 436100 998572
rect 436152 998560 436158 998572
rect 472434 998560 472440 998572
rect 436152 998532 472440 998560
rect 436152 998520 436158 998532
rect 472434 998520 472440 998532
rect 472492 998520 472498 998572
rect 500862 998520 500868 998572
rect 500920 998560 500926 998572
rect 517514 998560 517520 998572
rect 500920 998532 517520 998560
rect 500920 998520 500926 998532
rect 517514 998520 517520 998532
rect 517572 998520 517578 998572
rect 557442 998520 557448 998572
rect 557500 998560 557506 998572
rect 557500 998532 563054 998560
rect 557500 998520 557506 998532
rect 92382 998384 92388 998436
rect 92440 998424 92446 998436
rect 100018 998424 100024 998436
rect 92440 998396 100024 998424
rect 92440 998384 92446 998396
rect 100018 998384 100024 998396
rect 100076 998384 100082 998436
rect 143994 998384 144000 998436
rect 144052 998424 144058 998436
rect 155954 998424 155960 998436
rect 144052 998396 155960 998424
rect 144052 998384 144058 998396
rect 155954 998384 155960 998396
rect 156012 998384 156018 998436
rect 247494 998384 247500 998436
rect 247552 998424 247558 998436
rect 247552 998396 253934 998424
rect 247552 998384 247558 998396
rect 200850 998316 200856 998368
rect 200908 998356 200914 998368
rect 203518 998356 203524 998368
rect 200908 998328 203524 998356
rect 200908 998316 200914 998328
rect 203518 998316 203524 998328
rect 203576 998316 203582 998368
rect 246758 998248 246764 998300
rect 246816 998288 246822 998300
rect 252462 998288 252468 998300
rect 246816 998260 252468 998288
rect 246816 998248 246822 998260
rect 252462 998248 252468 998260
rect 252520 998248 252526 998300
rect 200022 998180 200028 998232
rect 200080 998220 200086 998232
rect 202690 998220 202696 998232
rect 200080 998192 202696 998220
rect 200080 998180 200086 998192
rect 202690 998180 202696 998192
rect 202748 998180 202754 998232
rect 250622 998112 250628 998164
rect 250680 998152 250686 998164
rect 253658 998152 253664 998164
rect 250680 998124 253664 998152
rect 250680 998112 250686 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 197354 998044 197360 998096
rect 197412 998084 197418 998096
rect 201862 998084 201868 998096
rect 197412 998056 201868 998084
rect 197412 998044 197418 998056
rect 201862 998044 201868 998056
rect 201920 998044 201926 998096
rect 202322 998044 202328 998096
rect 202380 998084 202386 998096
rect 205542 998084 205548 998096
rect 202380 998056 205548 998084
rect 202380 998044 202386 998056
rect 205542 998044 205548 998056
rect 205600 998044 205606 998096
rect 92750 997976 92756 998028
rect 92808 998016 92814 998028
rect 92808 997988 103514 998016
rect 92808 997976 92814 997988
rect 93486 997840 93492 997892
rect 93544 997880 93550 997892
rect 94682 997880 94688 997892
rect 93544 997852 94688 997880
rect 93544 997840 93550 997852
rect 94682 997840 94688 997852
rect 94740 997840 94746 997892
rect 103486 997880 103514 997988
rect 197998 997908 198004 997960
rect 198056 997948 198062 997960
rect 200666 997948 200672 997960
rect 198056 997920 200672 997948
rect 198056 997908 198062 997920
rect 200666 997908 200672 997920
rect 200724 997908 200730 997960
rect 202138 997908 202144 997960
rect 202196 997948 202202 997960
rect 204714 997948 204720 997960
rect 202196 997920 204720 997948
rect 202196 997908 202202 997920
rect 204714 997908 204720 997920
rect 204772 997908 204778 997960
rect 250438 997908 250444 997960
rect 250496 997948 250502 997960
rect 253658 997948 253664 997960
rect 250496 997920 253664 997948
rect 250496 997908 250502 997920
rect 253658 997908 253664 997920
rect 253716 997908 253722 997960
rect 121730 997880 121736 997892
rect 103486 997852 121736 997880
rect 121730 997840 121736 997852
rect 121788 997840 121794 997892
rect 195698 997772 195704 997824
rect 195756 997812 195762 997824
rect 226334 997812 226340 997824
rect 195756 997784 226340 997812
rect 195756 997772 195762 997784
rect 226334 997772 226340 997784
rect 226392 997772 226398 997824
rect 247678 997772 247684 997824
rect 247736 997812 247742 997824
rect 252462 997812 252468 997824
rect 247736 997784 252468 997812
rect 247736 997772 247742 997784
rect 252462 997772 252468 997784
rect 252520 997772 252526 997824
rect 253906 997812 253934 998396
rect 355318 998384 355324 998436
rect 355376 998424 355382 998436
rect 383470 998424 383476 998436
rect 355376 998396 383476 998424
rect 355376 998384 355382 998396
rect 383470 998384 383476 998396
rect 383528 998384 383534 998436
rect 431862 998384 431868 998436
rect 431920 998424 431926 998436
rect 471790 998424 471796 998436
rect 431920 998396 471796 998424
rect 431920 998384 431926 998396
rect 471790 998384 471796 998396
rect 471848 998384 471854 998436
rect 497918 998384 497924 998436
rect 497976 998424 497982 998436
rect 524046 998424 524052 998436
rect 497976 998396 524052 998424
rect 497976 998384 497982 998396
rect 524046 998384 524052 998396
rect 524104 998384 524110 998436
rect 555418 998384 555424 998436
rect 555476 998424 555482 998436
rect 558822 998424 558828 998436
rect 555476 998396 558828 998424
rect 555476 998384 555482 998396
rect 558822 998384 558828 998396
rect 558880 998384 558886 998436
rect 563026 998424 563054 998532
rect 572714 998424 572720 998436
rect 563026 998396 572720 998424
rect 572714 998384 572720 998396
rect 572772 998384 572778 998436
rect 378594 998248 378600 998300
rect 378652 998288 378658 998300
rect 382274 998288 382280 998300
rect 378652 998260 382280 998288
rect 378652 998248 378658 998260
rect 382274 998248 382280 998260
rect 382332 998248 382338 998300
rect 430022 998248 430028 998300
rect 430080 998288 430086 998300
rect 432598 998288 432604 998300
rect 430080 998260 432604 998288
rect 430080 998248 430086 998260
rect 432598 998248 432604 998260
rect 432656 998248 432662 998300
rect 506290 998248 506296 998300
rect 506348 998288 506354 998300
rect 517238 998288 517244 998300
rect 506348 998260 517244 998288
rect 506348 998248 506354 998260
rect 517238 998248 517244 998260
rect 517296 998248 517302 998300
rect 518158 998248 518164 998300
rect 518216 998288 518222 998300
rect 523862 998288 523868 998300
rect 518216 998260 523868 998288
rect 518216 998248 518222 998260
rect 523862 998248 523868 998260
rect 523920 998248 523926 998300
rect 557994 998248 558000 998300
rect 558052 998288 558058 998300
rect 560938 998288 560944 998300
rect 558052 998260 560944 998288
rect 558052 998248 558058 998260
rect 560938 998248 560944 998260
rect 560996 998248 561002 998300
rect 431218 998112 431224 998164
rect 431276 998152 431282 998164
rect 433518 998152 433524 998164
rect 431276 998124 433524 998152
rect 431276 998112 431282 998124
rect 433518 998112 433524 998124
rect 433576 998112 433582 998164
rect 558822 998112 558828 998164
rect 558880 998152 558886 998164
rect 562502 998152 562508 998164
rect 558880 998124 562508 998152
rect 558880 998112 558886 998124
rect 562502 998112 562508 998124
rect 562560 998112 562566 998164
rect 489270 998044 489276 998096
rect 489328 998084 489334 998096
rect 493962 998084 493968 998096
rect 489328 998056 493968 998084
rect 489328 998044 489334 998056
rect 493962 998044 493968 998056
rect 494020 998044 494026 998096
rect 591298 998044 591304 998096
rect 591356 998084 591362 998096
rect 625614 998084 625620 998096
rect 591356 998056 625620 998084
rect 591356 998044 591362 998056
rect 625614 998044 625620 998056
rect 625672 998044 625678 998096
rect 432046 997976 432052 998028
rect 432104 998016 432110 998028
rect 436738 998016 436744 998028
rect 432104 997988 436744 998016
rect 432104 997976 432110 997988
rect 436738 997976 436744 997988
rect 436796 997976 436802 998028
rect 557994 997976 558000 998028
rect 558052 998016 558058 998028
rect 560294 998016 560300 998028
rect 558052 997988 560300 998016
rect 558052 997976 558058 997988
rect 560294 997976 560300 997988
rect 560352 997976 560358 998028
rect 591114 997908 591120 997960
rect 591172 997948 591178 997960
rect 625798 997948 625804 997960
rect 591172 997920 625804 997948
rect 591172 997908 591178 997920
rect 625798 997908 625804 997920
rect 625856 997908 625862 997960
rect 557626 997840 557632 997892
rect 557684 997880 557690 997892
rect 559558 997880 559564 997892
rect 557684 997852 559564 997880
rect 557684 997840 557690 997852
rect 559558 997840 559564 997852
rect 559616 997840 559622 997892
rect 560018 997840 560024 997892
rect 560076 997880 560082 997892
rect 562318 997880 562324 997892
rect 560076 997852 562324 997880
rect 560076 997840 560082 997852
rect 562318 997840 562324 997852
rect 562376 997840 562382 997892
rect 253906 997784 277394 997812
rect 113818 997704 113824 997756
rect 113876 997744 113882 997756
rect 117130 997744 117136 997756
rect 113876 997716 117136 997744
rect 113876 997704 113882 997716
rect 117130 997704 117136 997716
rect 117188 997704 117194 997756
rect 143810 997704 143816 997756
rect 143868 997744 143874 997756
rect 160094 997744 160100 997756
rect 143868 997716 160100 997744
rect 143868 997704 143874 997716
rect 160094 997704 160100 997716
rect 160152 997704 160158 997756
rect 277366 997744 277394 997784
rect 430022 997772 430028 997824
rect 430080 997812 430086 997824
rect 432046 997812 432052 997824
rect 430080 997784 432052 997812
rect 430080 997772 430086 997784
rect 432046 997772 432052 997784
rect 432104 997772 432110 997824
rect 553946 997772 553952 997824
rect 554004 997812 554010 997824
rect 555602 997812 555608 997824
rect 554004 997784 555608 997812
rect 554004 997772 554010 997784
rect 555602 997772 555608 997784
rect 555660 997772 555666 997824
rect 592034 997772 592040 997824
rect 592092 997812 592098 997824
rect 625430 997812 625436 997824
rect 592092 997784 625436 997812
rect 592092 997772 592098 997784
rect 625430 997772 625436 997784
rect 625488 997772 625494 997824
rect 279234 997744 279240 997756
rect 277366 997716 279240 997744
rect 279234 997704 279240 997716
rect 279292 997704 279298 997756
rect 298462 997704 298468 997756
rect 298520 997744 298526 997756
rect 311894 997744 311900 997756
rect 298520 997716 311900 997744
rect 298520 997704 298526 997716
rect 311894 997704 311900 997716
rect 311952 997704 311958 997756
rect 355778 997704 355784 997756
rect 355836 997744 355842 997756
rect 372338 997744 372344 997756
rect 355836 997716 372344 997744
rect 355836 997704 355842 997716
rect 372338 997704 372344 997716
rect 372396 997704 372402 997756
rect 433978 997704 433984 997756
rect 434036 997744 434042 997756
rect 439682 997744 439688 997756
rect 434036 997716 439688 997744
rect 434036 997704 434042 997716
rect 439682 997704 439688 997716
rect 439740 997704 439746 997756
rect 489086 997704 489092 997756
rect 489144 997744 489150 997756
rect 509234 997744 509240 997756
rect 489144 997716 509240 997744
rect 489144 997704 489150 997716
rect 509234 997704 509240 997716
rect 509292 997704 509298 997756
rect 509694 997704 509700 997756
rect 509752 997744 509758 997756
rect 517054 997744 517060 997756
rect 509752 997716 517060 997744
rect 509752 997704 509758 997716
rect 517054 997704 517060 997716
rect 517112 997704 517118 997756
rect 558178 997704 558184 997756
rect 558236 997744 558242 997756
rect 562686 997744 562692 997756
rect 558236 997716 562692 997744
rect 558236 997704 558242 997716
rect 562686 997704 562692 997716
rect 562744 997704 562750 997756
rect 566642 997704 566648 997756
rect 566700 997744 566706 997756
rect 566700 997716 576854 997744
rect 566700 997704 566706 997716
rect 92566 997636 92572 997688
rect 92624 997676 92630 997688
rect 101582 997676 101588 997688
rect 92624 997648 101588 997676
rect 92624 997636 92630 997648
rect 101582 997636 101588 997648
rect 101640 997636 101646 997688
rect 248046 997636 248052 997688
rect 248104 997676 248110 997688
rect 259454 997676 259460 997688
rect 248104 997648 259460 997676
rect 248104 997636 248110 997648
rect 259454 997636 259460 997648
rect 259512 997636 259518 997688
rect 399938 997636 399944 997688
rect 399996 997676 400002 997688
rect 432046 997676 432052 997688
rect 399996 997648 432052 997676
rect 399996 997636 400002 997648
rect 432046 997636 432052 997648
rect 432104 997636 432110 997688
rect 552658 997636 552664 997688
rect 552716 997676 552722 997688
rect 576826 997676 576854 997716
rect 618162 997676 618168 997688
rect 552716 997648 557534 997676
rect 576826 997648 618168 997676
rect 552716 997636 552722 997648
rect 109494 997568 109500 997620
rect 109552 997608 109558 997620
rect 116118 997608 116124 997620
rect 109552 997580 116124 997608
rect 109552 997568 109558 997580
rect 116118 997568 116124 997580
rect 116176 997568 116182 997620
rect 144822 997568 144828 997620
rect 144880 997608 144886 997620
rect 153930 997608 153936 997620
rect 144880 997580 153936 997608
rect 144880 997568 144886 997580
rect 153930 997568 153936 997580
rect 153988 997568 153994 997620
rect 299198 997568 299204 997620
rect 299256 997608 299262 997620
rect 310514 997608 310520 997620
rect 299256 997580 310520 997608
rect 299256 997568 299262 997580
rect 310514 997568 310520 997580
rect 310572 997568 310578 997620
rect 365162 997568 365168 997620
rect 365220 997608 365226 997620
rect 372522 997608 372528 997620
rect 365220 997580 372528 997608
rect 365220 997568 365226 997580
rect 372522 997568 372528 997580
rect 372580 997568 372586 997620
rect 432598 997568 432604 997620
rect 432656 997608 432662 997620
rect 439866 997608 439872 997620
rect 432656 997580 439872 997608
rect 432656 997568 432662 997580
rect 439866 997568 439872 997580
rect 439924 997568 439930 997620
rect 488902 997568 488908 997620
rect 488960 997608 488966 997620
rect 510798 997608 510804 997620
rect 488960 997580 510804 997608
rect 488960 997568 488966 997580
rect 510798 997568 510804 997580
rect 510856 997568 510862 997620
rect 557506 997608 557534 997648
rect 618162 997636 618168 997648
rect 618220 997636 618226 997688
rect 562134 997608 562140 997620
rect 557506 997580 562140 997608
rect 562134 997568 562140 997580
rect 562192 997568 562198 997620
rect 571794 997608 571800 997620
rect 562520 997580 571800 997608
rect 246942 997500 246948 997552
rect 247000 997540 247006 997552
rect 255958 997540 255964 997552
rect 247000 997512 255964 997540
rect 247000 997500 247006 997512
rect 255958 997500 255964 997512
rect 256016 997500 256022 997552
rect 540882 997500 540888 997552
rect 540940 997540 540946 997552
rect 555418 997540 555424 997552
rect 540940 997512 555424 997540
rect 540940 997500 540946 997512
rect 555418 997500 555424 997512
rect 555476 997500 555482 997552
rect 508498 997432 508504 997484
rect 508556 997472 508562 997484
rect 516686 997472 516692 997484
rect 508556 997444 516692 997472
rect 508556 997432 508562 997444
rect 516686 997432 516692 997444
rect 516744 997432 516750 997484
rect 562520 997472 562548 997580
rect 571794 997568 571800 997580
rect 571852 997568 571858 997620
rect 557506 997444 562548 997472
rect 553302 997364 553308 997416
rect 553360 997404 553366 997416
rect 557506 997404 557534 997444
rect 562686 997432 562692 997484
rect 562744 997472 562750 997484
rect 571610 997472 571616 997484
rect 562744 997444 571616 997472
rect 562744 997432 562750 997444
rect 571610 997432 571616 997444
rect 571668 997432 571674 997484
rect 571978 997432 571984 997484
rect 572036 997472 572042 997484
rect 592034 997472 592040 997484
rect 572036 997444 592040 997472
rect 572036 997432 572042 997444
rect 592034 997432 592040 997444
rect 592092 997432 592098 997484
rect 553360 997376 557534 997404
rect 553360 997364 553366 997376
rect 562134 997296 562140 997348
rect 562192 997336 562198 997348
rect 591298 997336 591304 997348
rect 562192 997308 591304 997336
rect 562192 997296 562198 997308
rect 591298 997296 591304 997308
rect 591356 997296 591362 997348
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 440234 997160 440240 997212
rect 440292 997200 440298 997212
rect 445662 997200 445668 997212
rect 440292 997172 445668 997200
rect 440292 997160 440298 997172
rect 445662 997160 445668 997172
rect 445720 997160 445726 997212
rect 555602 997160 555608 997212
rect 555660 997200 555666 997212
rect 570414 997200 570420 997212
rect 555660 997172 570420 997200
rect 555660 997160 555666 997172
rect 570414 997160 570420 997172
rect 570472 997160 570478 997212
rect 571794 997160 571800 997212
rect 571852 997200 571858 997212
rect 590562 997200 590568 997212
rect 571852 997172 590568 997200
rect 571852 997160 571858 997172
rect 590562 997160 590568 997172
rect 590620 997160 590626 997212
rect 320818 997024 320824 997076
rect 320876 997064 320882 997076
rect 332594 997064 332600 997076
rect 320876 997036 332600 997064
rect 320876 997024 320882 997036
rect 332594 997024 332600 997036
rect 332652 997024 332658 997076
rect 356054 997024 356060 997076
rect 356112 997064 356118 997076
rect 372706 997064 372712 997076
rect 356112 997036 372712 997064
rect 356112 997024 356118 997036
rect 372706 997024 372712 997036
rect 372764 997024 372770 997076
rect 443638 997024 443644 997076
rect 443696 997064 443702 997076
rect 453850 997064 453856 997076
rect 443696 997036 453856 997064
rect 443696 997024 443702 997036
rect 453850 997024 453856 997036
rect 453908 997024 453914 997076
rect 502978 997024 502984 997076
rect 503036 997064 503042 997076
rect 516870 997064 516876 997076
rect 503036 997036 516876 997064
rect 503036 997024 503042 997036
rect 516870 997024 516876 997036
rect 516928 997024 516934 997076
rect 551922 997024 551928 997076
rect 551980 997064 551986 997076
rect 623682 997064 623688 997076
rect 551980 997036 623688 997064
rect 551980 997024 551986 997036
rect 623682 997024 623688 997036
rect 623740 997024 623746 997076
rect 143718 996888 143724 996940
rect 143776 996928 143782 996940
rect 151262 996928 151268 996940
rect 143776 996900 151268 996928
rect 143776 996888 143782 996900
rect 151262 996888 151268 996900
rect 151320 996888 151326 996940
rect 568482 996888 568488 996940
rect 568540 996928 568546 996940
rect 571058 996928 571064 996940
rect 568540 996900 571064 996928
rect 568540 996888 568546 996900
rect 571058 996888 571064 996900
rect 571116 996888 571122 996940
rect 571610 996888 571616 996940
rect 571668 996928 571674 996940
rect 572898 996928 572904 996940
rect 571668 996900 572904 996928
rect 571668 996888 571674 996900
rect 572898 996888 572904 996900
rect 572956 996888 572962 996940
rect 573358 996888 573364 996940
rect 573416 996928 573422 996940
rect 591114 996928 591120 996940
rect 573416 996900 591120 996928
rect 573416 996888 573422 996900
rect 591114 996888 591120 996900
rect 591172 996888 591178 996940
rect 153010 996820 153016 996872
rect 153068 996860 153074 996872
rect 158714 996860 158720 996872
rect 153068 996832 158720 996860
rect 153068 996820 153074 996832
rect 158714 996820 158720 996832
rect 158772 996820 158778 996872
rect 200206 996820 200212 996872
rect 200264 996860 200270 996872
rect 203702 996860 203708 996872
rect 200264 996832 203708 996860
rect 200264 996820 200270 996832
rect 203702 996820 203708 996832
rect 203760 996820 203766 996872
rect 571242 996752 571248 996804
rect 571300 996792 571306 996804
rect 590378 996792 590384 996804
rect 571300 996764 590384 996792
rect 571300 996752 571306 996764
rect 590378 996752 590384 996764
rect 590436 996752 590442 996804
rect 143810 996616 143816 996668
rect 143868 996656 143874 996668
rect 149882 996656 149888 996668
rect 143868 996628 149888 996656
rect 143868 996616 143874 996628
rect 149882 996616 149888 996628
rect 149940 996616 149946 996668
rect 570598 996616 570604 996668
rect 570656 996656 570662 996668
rect 570656 996628 586514 996656
rect 570656 996616 570662 996628
rect 144546 996480 144552 996532
rect 144604 996520 144610 996532
rect 149054 996520 149060 996532
rect 144604 996492 149060 996520
rect 144604 996480 144610 996492
rect 149054 996480 149060 996492
rect 149112 996480 149118 996532
rect 586486 996452 586514 996628
rect 590562 996452 590568 996464
rect 586486 996424 590568 996452
rect 590562 996412 590568 996424
rect 590620 996412 590626 996464
rect 195238 996344 195244 996396
rect 195296 996384 195302 996396
rect 197998 996384 198004 996396
rect 195296 996356 198004 996384
rect 195296 996344 195302 996356
rect 197998 996344 198004 996356
rect 198056 996344 198062 996396
rect 549438 996344 549444 996396
rect 549496 996384 549502 996396
rect 550634 996384 550640 996396
rect 549496 996356 550640 996384
rect 549496 996344 549502 996356
rect 550634 996344 550640 996356
rect 550692 996344 550698 996396
rect 262858 996276 262864 996328
rect 262916 996316 262922 996328
rect 270402 996316 270408 996328
rect 262916 996288 270408 996316
rect 262916 996276 262922 996288
rect 270402 996276 270408 996288
rect 270460 996276 270466 996328
rect 556154 996276 556160 996328
rect 556212 996316 556218 996328
rect 556212 996288 586514 996316
rect 556212 996276 556218 996288
rect 586486 996248 586514 996288
rect 590562 996248 590568 996260
rect 586486 996220 590568 996248
rect 590562 996208 590568 996220
rect 590620 996208 590626 996260
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 211154 996112 211160 996124
rect 171836 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 228358 996072 228364 996124
rect 228416 996112 228422 996124
rect 263594 996112 263600 996124
rect 228416 996084 263600 996112
rect 228416 996072 228422 996084
rect 263594 996072 263600 996084
rect 263652 996072 263658 996124
rect 264238 996072 264244 996124
rect 264296 996112 264302 996124
rect 299014 996112 299020 996124
rect 264296 996084 299020 996112
rect 264296 996072 264302 996084
rect 299014 996072 299020 996084
rect 299072 996072 299078 996124
rect 433518 996112 433524 996124
rect 385236 996084 433524 996112
rect 382918 996004 382924 996056
rect 382976 996044 382982 996056
rect 382976 996016 384804 996044
rect 382976 996004 382982 996016
rect 169386 995936 169392 995988
rect 169444 995976 169450 995988
rect 171686 995976 171692 995988
rect 169444 995948 171692 995976
rect 169444 995936 169450 995948
rect 171686 995936 171692 995948
rect 171744 995936 171750 995988
rect 213178 995936 213184 995988
rect 213236 995976 213242 995988
rect 261110 995976 261116 995988
rect 213236 995948 261116 995976
rect 213236 995936 213242 995948
rect 261110 995936 261116 995948
rect 261168 995936 261174 995988
rect 269758 995936 269764 995988
rect 269816 995976 269822 995988
rect 316034 995976 316040 995988
rect 269816 995948 316040 995976
rect 269816 995936 269822 995948
rect 316034 995936 316040 995948
rect 316092 995936 316098 995988
rect 354582 995936 354588 995988
rect 354640 995976 354646 995988
rect 381538 995976 381544 995988
rect 354640 995948 381544 995976
rect 354640 995936 354646 995948
rect 381538 995936 381544 995948
rect 381596 995936 381602 995988
rect 384776 995976 384804 996016
rect 385236 995976 385264 996084
rect 433518 996072 433524 996084
rect 433576 996072 433582 996124
rect 511258 996072 511264 996124
rect 511316 996112 511322 996124
rect 563054 996112 563060 996124
rect 511316 996084 563060 996112
rect 511316 996072 511322 996084
rect 563054 996072 563060 996084
rect 563112 996072 563118 996124
rect 384776 995948 385264 995976
rect 522298 995936 522304 995988
rect 522356 995976 522362 995988
rect 560294 995976 560300 995988
rect 522356 995948 560300 995976
rect 522356 995936 522362 995948
rect 560294 995936 560300 995948
rect 560352 995936 560358 995988
rect 202966 995868 202972 995920
rect 203024 995908 203030 995920
rect 205082 995908 205088 995920
rect 203024 995880 205088 995908
rect 203024 995868 203030 995880
rect 205082 995868 205088 995880
rect 205140 995868 205146 995920
rect 386386 995880 389174 995908
rect 140774 995800 140780 995852
rect 140832 995840 140838 995852
rect 143994 995840 144000 995852
rect 140832 995812 144000 995840
rect 140832 995800 140838 995812
rect 143994 995800 144000 995812
rect 144052 995800 144058 995852
rect 170674 995800 170680 995852
rect 170732 995840 170738 995852
rect 171226 995840 171232 995852
rect 170732 995812 171232 995840
rect 170732 995800 170738 995812
rect 171226 995800 171232 995812
rect 171284 995800 171290 995852
rect 229738 995800 229744 995852
rect 229796 995840 229802 995852
rect 262214 995840 262220 995852
rect 229796 995812 262220 995840
rect 229796 995800 229802 995812
rect 262214 995800 262220 995812
rect 262272 995800 262278 995852
rect 364978 995800 364984 995852
rect 365036 995840 365042 995852
rect 386386 995840 386414 995880
rect 365036 995812 386414 995840
rect 389146 995840 389174 995880
rect 400858 995840 400864 995852
rect 389146 995812 400864 995840
rect 365036 995800 365042 995812
rect 400858 995800 400864 995812
rect 400916 995800 400922 995852
rect 170858 995528 170864 995580
rect 170916 995568 170922 995580
rect 170916 995540 171916 995568
rect 170916 995528 170922 995540
rect 171888 995415 171916 995540
rect 246206 995528 246212 995580
rect 246264 995568 246270 995580
rect 247126 995568 247132 995580
rect 246264 995540 247132 995568
rect 246264 995528 246270 995540
rect 247126 995528 247132 995540
rect 247184 995528 247190 995580
rect 297818 995528 297824 995580
rect 297876 995568 297882 995580
rect 299382 995568 299388 995580
rect 297876 995540 299388 995568
rect 297876 995528 297882 995540
rect 299382 995528 299388 995540
rect 299440 995528 299446 995580
rect 380158 995528 380164 995580
rect 380216 995568 380222 995580
rect 383102 995568 383108 995580
rect 380216 995540 383108 995568
rect 380216 995528 380222 995540
rect 383102 995528 383108 995540
rect 383160 995528 383166 995580
rect 383286 995528 383292 995580
rect 383344 995568 383350 995580
rect 384758 995568 384764 995580
rect 383344 995540 384764 995568
rect 383344 995528 383350 995540
rect 384758 995528 384764 995540
rect 384816 995528 384822 995580
rect 385402 995528 385408 995580
rect 385460 995568 385466 995580
rect 386966 995568 386972 995580
rect 385460 995540 386972 995568
rect 385460 995528 385466 995540
rect 386966 995528 386972 995540
rect 387024 995528 387030 995580
rect 472710 995528 472716 995580
rect 472768 995568 472774 995580
rect 473998 995568 474004 995580
rect 472768 995540 474004 995568
rect 472768 995528 472774 995540
rect 473998 995528 474004 995540
rect 474056 995528 474062 995580
rect 493962 995528 493968 995580
rect 494020 995568 494026 995580
rect 511074 995568 511080 995580
rect 494020 995540 511080 995568
rect 494020 995528 494026 995540
rect 511074 995528 511080 995540
rect 511132 995528 511138 995580
rect 524046 995528 524052 995580
rect 524104 995568 524110 995580
rect 526070 995568 526076 995580
rect 524104 995540 526076 995568
rect 524104 995528 524110 995540
rect 526070 995528 526076 995540
rect 526128 995528 526134 995580
rect 625798 995528 625804 995580
rect 625856 995568 625862 995580
rect 626534 995568 626540 995580
rect 625856 995540 626540 995568
rect 625856 995528 625862 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 194870 995460 194876 995512
rect 194928 995500 194934 995512
rect 195514 995500 195520 995512
rect 194928 995472 195520 995500
rect 194928 995460 194934 995472
rect 195514 995460 195520 995472
rect 195572 995460 195578 995512
rect 475930 995460 475936 995512
rect 475988 995500 475994 995512
rect 476390 995500 476396 995512
rect 475988 995472 476396 995500
rect 475988 995460 475994 995472
rect 476390 995460 476396 995472
rect 476448 995460 476454 995512
rect 476942 995460 476948 995512
rect 477000 995500 477006 995512
rect 478966 995500 478972 995512
rect 477000 995472 478972 995500
rect 477000 995460 477006 995472
rect 478966 995460 478972 995472
rect 479024 995460 479030 995512
rect 211798 995392 211804 995444
rect 211856 995432 211862 995444
rect 260926 995432 260932 995444
rect 211856 995404 260932 995432
rect 211856 995392 211862 995404
rect 260926 995392 260932 995404
rect 260984 995392 260990 995444
rect 292546 995404 306374 995432
rect 171686 995277 171692 995329
rect 171744 995277 171750 995329
rect 180702 995324 180708 995376
rect 180760 995364 180766 995376
rect 202322 995364 202328 995376
rect 180760 995336 202328 995364
rect 180760 995324 180766 995336
rect 202322 995324 202328 995336
rect 202380 995324 202386 995376
rect 290642 995324 290648 995376
rect 290700 995364 290706 995376
rect 292546 995364 292574 995404
rect 290700 995336 292574 995364
rect 290700 995324 290706 995336
rect 296162 995256 296168 995308
rect 296220 995296 296226 995308
rect 298646 995296 298652 995308
rect 296220 995268 298652 995296
rect 296220 995256 296226 995268
rect 298646 995256 298652 995268
rect 298704 995256 298710 995308
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 182956 995188 182962 995240
rect 183014 995228 183020 995240
rect 208578 995228 208584 995240
rect 183014 995200 208584 995228
rect 183014 995188 183020 995200
rect 208578 995188 208584 995200
rect 208636 995188 208642 995240
rect 236224 995188 236230 995240
rect 236282 995228 236288 995240
rect 251818 995228 251824 995240
rect 236282 995200 251824 995228
rect 236282 995188 236288 995200
rect 251818 995188 251824 995200
rect 251876 995188 251882 995240
rect 290826 995188 290832 995240
rect 290884 995228 290890 995240
rect 295518 995228 295524 995240
rect 290884 995200 295524 995228
rect 290884 995188 290890 995200
rect 295518 995188 295524 995200
rect 295576 995188 295582 995240
rect 306346 995228 306374 995404
rect 366358 995392 366364 995444
rect 366416 995432 366422 995444
rect 402238 995432 402244 995444
rect 366416 995404 402244 995432
rect 366416 995392 366422 995404
rect 402238 995392 402244 995404
rect 402296 995392 402302 995444
rect 415394 995392 415400 995444
rect 415452 995432 415458 995444
rect 415452 995404 415716 995432
rect 415452 995392 415458 995404
rect 415688 995387 415716 995404
rect 402790 995324 402796 995376
rect 402848 995364 402854 995376
rect 402974 995364 402980 995376
rect 402848 995336 402980 995364
rect 402848 995324 402854 995336
rect 402974 995324 402980 995336
rect 403032 995324 403038 995376
rect 415688 995359 415978 995387
rect 362218 995256 362224 995308
rect 362276 995296 362282 995308
rect 394602 995296 394608 995308
rect 362276 995268 394608 995296
rect 362276 995256 362282 995268
rect 394602 995256 394608 995268
rect 394660 995256 394666 995308
rect 307018 995228 307024 995240
rect 306346 995200 307024 995228
rect 307018 995188 307024 995200
rect 307076 995188 307082 995240
rect 416130 995235 416136 995287
rect 416188 995235 416194 995287
rect 384298 995160 384304 995172
rect 373966 995132 384304 995160
rect 171232 995105 171284 995111
rect 171232 995047 171284 995053
rect 180150 995052 180156 995104
rect 180208 995092 180214 995104
rect 206278 995092 206284 995104
rect 180208 995064 206284 995092
rect 180208 995052 180214 995064
rect 206278 995052 206284 995064
rect 206336 995052 206342 995104
rect 231578 995052 231584 995104
rect 231636 995092 231642 995104
rect 257338 995092 257344 995104
rect 231636 995064 257344 995092
rect 231636 995052 231642 995064
rect 257338 995052 257344 995064
rect 257396 995052 257402 995104
rect 283466 995052 283472 995104
rect 283524 995092 283530 995104
rect 305638 995092 305644 995104
rect 283524 995064 305644 995092
rect 283524 995052 283530 995064
rect 305638 995052 305644 995064
rect 305696 995052 305702 995104
rect 363598 994984 363604 995036
rect 363656 995024 363662 995036
rect 373966 995024 373994 995132
rect 384298 995120 384304 995132
rect 384356 995120 384362 995172
rect 392118 995160 392124 995172
rect 384500 995132 392124 995160
rect 363656 994996 373994 995024
rect 363656 994984 363662 994996
rect 374362 994984 374368 995036
rect 374420 995024 374426 995036
rect 384500 995024 384528 995132
rect 392118 995120 392124 995132
rect 392176 995120 392182 995172
rect 537754 995120 537760 995172
rect 537812 995160 537818 995172
rect 538398 995160 538404 995172
rect 537812 995132 538404 995160
rect 537812 995120 537818 995132
rect 538398 995120 538404 995132
rect 538456 995120 538462 995172
rect 660304 995147 660356 995153
rect 455874 995052 455880 995104
rect 455932 995092 455938 995104
rect 487798 995092 487804 995104
rect 455932 995064 487804 995092
rect 455932 995052 455938 995064
rect 487798 995052 487804 995064
rect 487856 995052 487862 995104
rect 517698 995052 517704 995104
rect 517756 995092 517762 995104
rect 533706 995092 533712 995104
rect 517756 995064 533712 995092
rect 517756 995052 517762 995064
rect 533706 995052 533712 995064
rect 533764 995052 533770 995104
rect 572714 995052 572720 995104
rect 572772 995092 572778 995104
rect 635826 995092 635832 995104
rect 572772 995064 635832 995092
rect 572772 995052 572778 995064
rect 635826 995052 635832 995064
rect 635884 995052 635890 995104
rect 638862 995052 638868 995104
rect 638920 995092 638926 995104
rect 640794 995092 640800 995104
rect 638920 995064 640800 995092
rect 638920 995052 638926 995064
rect 640794 995052 640800 995064
rect 640852 995052 640858 995104
rect 660304 995089 660356 995095
rect 374420 994996 384528 995024
rect 374420 994984 374426 994996
rect 384666 994984 384672 995036
rect 384724 995024 384730 995036
rect 387794 995024 387800 995036
rect 384724 994996 387800 995024
rect 384724 994984 384730 994996
rect 387794 994984 387800 994996
rect 387852 994984 387858 995036
rect 387978 994984 387984 995036
rect 388036 995024 388042 995036
rect 389358 995024 389364 995036
rect 388036 994996 389364 995024
rect 388036 994984 388042 994996
rect 389358 994984 389364 994996
rect 389416 994984 389422 995036
rect 389542 994984 389548 995036
rect 389600 995024 389606 995036
rect 398834 995024 398840 995036
rect 389600 994996 398840 995024
rect 389600 994984 389606 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 641732 995023 660252 995024
rect 641732 994996 660606 995023
rect 171244 994881 171272 994967
rect 183830 994916 183836 994968
rect 183888 994956 183894 994968
rect 202138 994956 202144 994968
rect 183888 994928 202144 994956
rect 183888 994916 183894 994928
rect 202138 994916 202144 994928
rect 202196 994916 202202 994968
rect 232222 994916 232228 994968
rect 232280 994956 232286 994968
rect 254578 994956 254584 994968
rect 232280 994928 254584 994956
rect 232280 994916 232286 994928
rect 254578 994916 254584 994928
rect 254636 994916 254642 994968
rect 284110 994916 284116 994968
rect 284168 994956 284174 994968
rect 308398 994956 308404 994968
rect 284168 994928 308404 994956
rect 284168 994916 284174 994928
rect 308398 994916 308404 994928
rect 308456 994916 308462 994968
rect 420822 994916 420828 994968
rect 420880 994956 420886 994968
rect 641732 994956 641760 994996
rect 660224 994995 660606 994996
rect 420880 994928 641760 994956
rect 420880 994916 420886 994928
rect 78306 994780 78312 994832
rect 78364 994820 78370 994832
rect 104158 994820 104164 994832
rect 78364 994792 104164 994820
rect 78364 994780 78370 994792
rect 104158 994780 104164 994792
rect 104216 994780 104222 994832
rect 128446 994780 128452 994832
rect 128504 994820 128510 994832
rect 157334 994820 157340 994832
rect 128504 994792 157340 994820
rect 128504 994780 128510 994792
rect 157334 994780 157340 994792
rect 157392 994780 157398 994832
rect 170490 994712 170496 994764
rect 170548 994752 170554 994764
rect 170876 994752 170904 994855
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 360838 994848 360844 994900
rect 360896 994888 360902 994900
rect 402974 994888 402980 994900
rect 360896 994860 402980 994888
rect 360896 994848 360902 994860
rect 402974 994848 402980 994860
rect 403032 994848 403038 994900
rect 243262 994780 243268 994832
rect 243320 994820 243326 994832
rect 246666 994820 246672 994832
rect 243320 994792 246672 994820
rect 243320 994780 243326 994792
rect 246666 994780 246672 994792
rect 246724 994780 246730 994832
rect 293218 994780 293224 994832
rect 293276 994820 293282 994832
rect 298462 994820 298468 994832
rect 293276 994792 298468 994820
rect 293276 994780 293282 994792
rect 298462 994780 298468 994792
rect 298520 994780 298526 994832
rect 453850 994780 453856 994832
rect 453908 994820 453914 994832
rect 489914 994820 489920 994832
rect 453908 994792 489920 994820
rect 453908 994780 453914 994792
rect 489914 994780 489920 994792
rect 489972 994780 489978 994832
rect 496722 994780 496728 994832
rect 496780 994820 496786 994832
rect 538214 994820 538220 994832
rect 496780 994792 538220 994820
rect 496780 994780 496786 994792
rect 538214 994780 538220 994792
rect 538272 994780 538278 994832
rect 567838 994780 567844 994832
rect 567896 994820 567902 994832
rect 639046 994820 639052 994832
rect 567896 994792 639052 994820
rect 567896 994780 567902 994792
rect 639046 994780 639052 994792
rect 639104 994780 639110 994832
rect 170548 994724 170904 994752
rect 170548 994712 170554 994724
rect 171042 994712 171048 994764
rect 171100 994752 171106 994764
rect 243078 994752 243084 994764
rect 171100 994724 243084 994752
rect 171100 994712 171106 994724
rect 243078 994712 243084 994724
rect 243136 994712 243142 994764
rect 372706 994712 372712 994764
rect 372764 994752 372770 994764
rect 393314 994752 393320 994764
rect 372764 994724 393320 994752
rect 372764 994712 372770 994724
rect 393314 994712 393320 994724
rect 393372 994712 393378 994764
rect 397638 994712 397644 994764
rect 397696 994752 397702 994764
rect 402790 994752 402796 994764
rect 397696 994724 402796 994752
rect 397696 994712 397702 994724
rect 402790 994712 402796 994724
rect 402848 994712 402854 994764
rect 81342 994644 81348 994696
rect 81400 994684 81406 994696
rect 98638 994684 98644 994696
rect 81400 994656 98644 994684
rect 81400 994644 81406 994656
rect 98638 994644 98644 994656
rect 98696 994644 98702 994696
rect 129090 994644 129096 994696
rect 129148 994684 129154 994696
rect 142108 994684 142114 994696
rect 129148 994656 142114 994684
rect 129148 994644 129154 994656
rect 142108 994644 142114 994656
rect 142166 994644 142172 994696
rect 419442 994644 419448 994696
rect 419500 994684 419506 994696
rect 660298 994684 660304 994696
rect 419500 994656 660304 994684
rect 419500 994644 419506 994656
rect 660298 994644 660304 994656
rect 660356 994644 660362 994696
rect 660776 994628 660804 994897
rect 149698 994616 149704 994628
rect 142264 994588 149704 994616
rect 77662 994508 77668 994560
rect 77720 994548 77726 994560
rect 93302 994548 93308 994560
rect 77720 994520 93308 994548
rect 77720 994508 77726 994520
rect 93302 994508 93308 994520
rect 93360 994508 93366 994560
rect 129734 994508 129740 994560
rect 129792 994548 129798 994560
rect 134886 994548 134892 994560
rect 129792 994520 134892 994548
rect 129792 994508 129798 994520
rect 134886 994508 134892 994520
rect 134944 994508 134950 994560
rect 135088 994520 142154 994548
rect 132402 994372 132408 994424
rect 132460 994412 132466 994424
rect 135088 994412 135116 994520
rect 142126 994480 142154 994520
rect 142264 994480 142292 994588
rect 149698 994576 149704 994588
rect 149756 994576 149762 994628
rect 170858 994576 170864 994628
rect 170916 994616 170922 994628
rect 300118 994616 300124 994628
rect 170916 994588 300124 994616
rect 170916 994576 170922 994588
rect 300118 994576 300124 994588
rect 300176 994576 300182 994628
rect 377398 994576 377404 994628
rect 377456 994616 377462 994628
rect 396994 994616 397000 994628
rect 377456 994588 397000 994616
rect 377456 994576 377462 994588
rect 396994 994576 397000 994588
rect 397052 994576 397058 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 472250 994508 472256 994560
rect 472308 994548 472314 994560
rect 474918 994548 474924 994560
rect 472308 994520 474924 994548
rect 472308 994508 472314 994520
rect 474918 994508 474924 994520
rect 474976 994508 474982 994560
rect 481634 994508 481640 994560
rect 481692 994548 481698 994560
rect 489730 994548 489736 994560
rect 481692 994520 489736 994548
rect 481692 994508 481698 994520
rect 489730 994508 489736 994520
rect 489788 994508 489794 994560
rect 499482 994508 499488 994560
rect 499540 994548 499546 994560
rect 538582 994548 538588 994560
rect 499540 994520 538588 994548
rect 499540 994508 499546 994520
rect 538582 994508 538588 994520
rect 538640 994508 538646 994560
rect 571058 994508 571064 994560
rect 571116 994548 571122 994560
rect 639506 994548 639512 994560
rect 571116 994520 639512 994548
rect 571116 994508 571122 994520
rect 639506 994508 639512 994520
rect 639564 994508 639570 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 153010 994480 153016 994492
rect 142126 994452 142292 994480
rect 146956 994452 153016 994480
rect 132460 994384 135116 994412
rect 132460 994372 132466 994384
rect 134886 994236 134892 994288
rect 134944 994276 134950 994288
rect 146956 994276 146984 994452
rect 153010 994440 153016 994452
rect 153068 994440 153074 994492
rect 170674 994440 170680 994492
rect 170732 994480 170738 994492
rect 250438 994480 250444 994492
rect 170732 994452 250444 994480
rect 170732 994440 170738 994452
rect 250438 994440 250444 994452
rect 250496 994440 250502 994492
rect 383102 994440 383108 994492
rect 383160 994480 383166 994492
rect 389542 994480 389548 994492
rect 383160 994452 389548 994480
rect 383160 994440 383166 994452
rect 389542 994440 389548 994452
rect 389600 994440 389606 994492
rect 279234 994372 279240 994424
rect 279292 994412 279298 994424
rect 316402 994412 316408 994424
rect 279292 994384 316408 994412
rect 279292 994372 279298 994384
rect 316402 994372 316408 994384
rect 316460 994372 316466 994424
rect 468478 994372 468484 994424
rect 468536 994412 468542 994424
rect 484118 994412 484124 994424
rect 468536 994384 484124 994412
rect 468536 994372 468542 994384
rect 484118 994372 484124 994384
rect 484176 994372 484182 994424
rect 505738 994372 505744 994424
rect 505796 994412 505802 994424
rect 505796 994384 509234 994412
rect 505796 994372 505802 994384
rect 149054 994304 149060 994356
rect 149112 994344 149118 994356
rect 186130 994344 186136 994356
rect 149112 994316 186136 994344
rect 149112 994304 149118 994316
rect 186130 994304 186136 994316
rect 186188 994304 186194 994356
rect 186268 994304 186274 994356
rect 186326 994344 186332 994356
rect 195790 994344 195796 994356
rect 186326 994316 195796 994344
rect 186326 994304 186332 994316
rect 195790 994304 195796 994316
rect 195848 994304 195854 994356
rect 134944 994248 146984 994276
rect 134944 994236 134950 994248
rect 226334 994236 226340 994288
rect 226392 994276 226398 994288
rect 251450 994276 251456 994288
rect 226392 994248 251456 994276
rect 226392 994236 226398 994248
rect 251450 994236 251456 994248
rect 251508 994236 251514 994288
rect 294506 994236 294512 994288
rect 294564 994276 294570 994288
rect 381170 994276 381176 994288
rect 294564 994248 381176 994276
rect 294564 994236 294570 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 414474 994236 414480 994288
rect 414532 994276 414538 994288
rect 446122 994276 446128 994288
rect 414532 994248 446128 994276
rect 414532 994236 414538 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 471606 994236 471612 994288
rect 471664 994276 471670 994288
rect 476298 994276 476304 994288
rect 471664 994248 476304 994276
rect 471664 994236 471670 994248
rect 476298 994236 476304 994248
rect 476356 994236 476362 994288
rect 509206 994276 509234 994384
rect 519538 994372 519544 994424
rect 519596 994412 519602 994424
rect 538398 994412 538404 994424
rect 519596 994384 538404 994412
rect 519596 994372 519602 994384
rect 538398 994372 538404 994384
rect 538456 994372 538462 994424
rect 572898 994372 572904 994424
rect 572956 994412 572962 994424
rect 590562 994412 590568 994424
rect 572956 994384 590568 994412
rect 572956 994372 572962 994384
rect 590562 994372 590568 994384
rect 590620 994372 590626 994424
rect 625246 994372 625252 994424
rect 625304 994412 625310 994424
rect 631502 994412 631508 994424
rect 625304 994384 631508 994412
rect 625304 994372 625310 994384
rect 631502 994372 631508 994384
rect 631560 994372 631566 994424
rect 528738 994276 528744 994288
rect 509206 994248 528744 994276
rect 528738 994236 528744 994248
rect 528796 994236 528802 994288
rect 539226 994276 539232 994288
rect 538186 994248 539232 994276
rect 169386 994168 169392 994220
rect 169444 994208 169450 994220
rect 169444 994180 176654 994208
rect 169444 994168 169450 994180
rect 142338 994100 142344 994152
rect 142396 994140 142402 994152
rect 151078 994140 151084 994152
rect 142396 994112 151084 994140
rect 142396 994100 142402 994112
rect 151078 994100 151084 994112
rect 151136 994100 151142 994152
rect 176626 994140 176654 994180
rect 298830 994140 298836 994152
rect 176626 994112 298836 994140
rect 298830 994100 298836 994112
rect 298888 994100 298894 994152
rect 471790 994100 471796 994152
rect 471848 994140 471854 994152
rect 475930 994140 475936 994152
rect 471848 994112 475936 994140
rect 471848 994100 471854 994112
rect 475930 994100 475936 994112
rect 475988 994100 475994 994152
rect 522114 994100 522120 994152
rect 522172 994140 522178 994152
rect 538186 994140 538214 994248
rect 539226 994236 539232 994248
rect 539284 994236 539290 994288
rect 550634 994236 550640 994288
rect 550692 994276 550698 994288
rect 572714 994276 572720 994288
rect 550692 994248 572720 994276
rect 550692 994236 550698 994248
rect 572714 994236 572720 994248
rect 572772 994236 572778 994288
rect 522172 994112 538214 994140
rect 522172 994100 522178 994112
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 141970 993964 141976 994016
rect 142028 994004 142034 994016
rect 142338 994004 142344 994016
rect 142028 993976 142344 994004
rect 142028 993964 142034 993976
rect 142338 993964 142344 993976
rect 142396 993964 142402 994016
rect 181438 993964 181444 994016
rect 181496 994004 181502 994016
rect 184290 994004 184296 994016
rect 181496 993976 184296 994004
rect 181496 993964 181502 993976
rect 184290 993964 184296 993976
rect 184348 993964 184354 994016
rect 184474 993964 184480 994016
rect 184532 994004 184538 994016
rect 186130 994004 186136 994016
rect 184532 993976 186136 994004
rect 184532 993964 184538 993976
rect 186130 993964 186136 993976
rect 186188 993964 186194 994016
rect 186268 993964 186274 994016
rect 186326 994004 186332 994016
rect 186326 993976 190960 994004
rect 186326 993964 186332 993976
rect 137554 993828 137560 993880
rect 137612 993868 137618 993880
rect 141786 993868 141792 993880
rect 137612 993840 141792 993868
rect 137612 993828 137618 993840
rect 141786 993828 141792 993840
rect 141844 993828 141850 993880
rect 187602 993828 187608 993880
rect 187660 993868 187666 993880
rect 190730 993868 190736 993880
rect 187660 993840 190736 993868
rect 187660 993828 187666 993840
rect 190730 993828 190736 993840
rect 190788 993828 190794 993880
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 187418 993800 187424 993812
rect 171284 993772 187424 993800
rect 171284 993760 171290 993772
rect 187418 993760 187424 993772
rect 187476 993760 187482 993812
rect 190932 993800 190960 993976
rect 191098 993964 191104 994016
rect 191156 994004 191162 994016
rect 203518 994004 203524 994016
rect 191156 993976 203524 994004
rect 191156 993964 191162 993976
rect 203518 993964 203524 993976
rect 203576 993964 203582 994016
rect 232866 993964 232872 994016
rect 232924 994004 232930 994016
rect 258074 994004 258080 994016
rect 232924 993976 258080 994004
rect 232924 993964 232930 993976
rect 258074 993964 258080 993976
rect 258132 993964 258138 994016
rect 471974 993964 471980 994016
rect 472032 994004 472038 994016
rect 477310 994004 477316 994016
rect 472032 993976 477316 994004
rect 472032 993964 472038 993976
rect 477310 993964 477316 993976
rect 477368 993964 477374 994016
rect 569218 993896 569224 993948
rect 569276 993936 569282 993948
rect 661328 993936 661356 994561
rect 569276 993908 661356 993936
rect 569276 993896 569282 993908
rect 207014 993868 207020 993880
rect 191116 993840 207020 993868
rect 191116 993800 191144 993840
rect 207014 993828 207020 993840
rect 207072 993828 207078 993880
rect 243078 993828 243084 993880
rect 243136 993868 243142 993880
rect 247678 993868 247684 993880
rect 243136 993840 247684 993868
rect 243136 993828 243142 993840
rect 247678 993828 247684 993840
rect 247736 993828 247742 993880
rect 190932 993772 191144 993800
rect 521286 993760 521292 993812
rect 521344 993800 521350 993812
rect 660942 993800 660948 993812
rect 521344 993772 660948 993800
rect 521344 993760 521350 993772
rect 660942 993760 660948 993772
rect 661000 993760 661006 993812
rect 195928 993692 195934 993744
rect 195986 993732 195992 993744
rect 196802 993732 196808 993744
rect 195986 993704 196808 993732
rect 195986 993692 195992 993704
rect 196802 993692 196808 993704
rect 196860 993692 196866 993744
rect 170490 993624 170496 993676
rect 170548 993664 170554 993676
rect 197354 993664 197360 993676
rect 170548 993636 195836 993664
rect 170548 993624 170554 993636
rect 195808 993596 195836 993636
rect 197004 993636 197360 993664
rect 195808 993568 195974 993596
rect 190546 993488 190552 993540
rect 190604 993528 190610 993540
rect 194870 993528 194876 993540
rect 190604 993500 194876 993528
rect 190604 993488 190610 993500
rect 194870 993488 194876 993500
rect 194928 993488 194934 993540
rect 195946 993460 195974 993568
rect 197004 993460 197032 993636
rect 197354 993624 197360 993636
rect 197412 993624 197418 993676
rect 517238 993624 517244 993676
rect 517296 993664 517302 993676
rect 660758 993664 660764 993676
rect 517296 993636 660764 993664
rect 517296 993624 517302 993636
rect 660758 993624 660764 993636
rect 660816 993624 660822 993676
rect 195946 993432 197032 993460
rect 50338 993148 50344 993200
rect 50396 993188 50402 993200
rect 107746 993188 107752 993200
rect 50396 993160 107752 993188
rect 50396 993148 50402 993160
rect 107746 993148 107752 993160
rect 107804 993148 107810 993200
rect 44818 993012 44824 993064
rect 44876 993052 44882 993064
rect 109034 993052 109040 993064
rect 44876 993024 109040 993052
rect 44876 993012 44882 993024
rect 109034 993012 109040 993024
rect 109092 993012 109098 993064
rect 318058 993012 318064 993064
rect 318116 993052 318122 993064
rect 349154 993052 349160 993064
rect 318116 993024 349160 993052
rect 318116 993012 318122 993024
rect 349154 993012 349160 993024
rect 349212 993012 349218 993064
rect 562502 993012 562508 993064
rect 562560 993052 562566 993064
rect 660298 993052 660304 993064
rect 562560 993024 660304 993052
rect 562560 993012 562566 993024
rect 660298 993012 660304 993024
rect 660356 993012 660362 993064
rect 54478 992876 54484 992928
rect 54536 992916 54542 992928
rect 148318 992916 148324 992928
rect 54536 992888 148324 992916
rect 54536 992876 54542 992888
rect 148318 992876 148324 992888
rect 148376 992876 148382 992928
rect 319438 992876 319444 992928
rect 319496 992916 319502 992928
rect 364978 992916 364984 992928
rect 319496 992888 364984 992916
rect 319496 992876 319502 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 560938 992876 560944 992928
rect 560996 992916 561002 992928
rect 667198 992916 667204 992928
rect 560996 992888 667204 992916
rect 560996 992876 561002 992888
rect 667198 992876 667204 992888
rect 667256 992876 667262 992928
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 51718 991584 51724 991636
rect 51776 991624 51782 991636
rect 110414 991624 110420 991636
rect 51776 991596 110420 991624
rect 51776 991584 51782 991596
rect 110414 991584 110420 991596
rect 110472 991584 110478 991636
rect 138290 991584 138296 991636
rect 138348 991624 138354 991636
rect 163130 991624 163136 991636
rect 138348 991596 163136 991624
rect 138348 991584 138354 991596
rect 163130 991584 163136 991596
rect 163188 991584 163194 991636
rect 369118 991584 369124 991636
rect 369176 991624 369182 991636
rect 414106 991624 414112 991636
rect 369176 991596 414112 991624
rect 369176 991584 369182 991596
rect 414106 991584 414112 991596
rect 414164 991584 414170 991636
rect 55858 991448 55864 991500
rect 55916 991488 55922 991500
rect 146938 991488 146944 991500
rect 55916 991460 146944 991488
rect 55916 991448 55922 991460
rect 146938 991448 146944 991460
rect 146996 991448 147002 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 430298 991488 430304 991500
rect 367796 991460 430304 991488
rect 367796 991448 367802 991460
rect 430298 991448 430304 991460
rect 430356 991448 430362 991500
rect 435358 991448 435364 991500
rect 435416 991488 435422 991500
rect 478966 991488 478972 991500
rect 435416 991460 478972 991488
rect 435416 991448 435422 991460
rect 478966 991448 478972 991460
rect 479024 991448 479030 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 214558 991176 214564 991228
rect 214616 991216 214622 991228
rect 219434 991216 219440 991228
rect 214616 991188 219440 991216
rect 214616 991176 214622 991188
rect 219434 991176 219440 991188
rect 219492 991176 219498 991228
rect 164878 990836 164884 990888
rect 164936 990876 164942 990888
rect 170766 990876 170772 990888
rect 164936 990848 170772 990876
rect 164936 990836 164942 990848
rect 170766 990836 170772 990848
rect 170824 990836 170830 990888
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 572714 990836 572720 990888
rect 572772 990876 572778 990888
rect 576302 990876 576308 990888
rect 572772 990848 576308 990876
rect 572772 990836 572778 990848
rect 576302 990836 576308 990848
rect 576360 990836 576366 990888
rect 53282 990224 53288 990276
rect 53340 990264 53346 990276
rect 95878 990264 95884 990276
rect 53340 990236 95884 990264
rect 53340 990224 53346 990236
rect 95878 990224 95884 990236
rect 95936 990224 95942 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 108114 990128 108120 990140
rect 49016 990100 108120 990128
rect 49016 990088 49022 990100
rect 108114 990088 108120 990100
rect 108172 990088 108178 990140
rect 512638 990088 512644 990140
rect 512696 990128 512702 990140
rect 543826 990128 543832 990140
rect 512696 990100 543832 990128
rect 512696 990088 512702 990100
rect 543826 990088 543832 990100
rect 543884 990088 543890 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 668578 990128 668584 990140
rect 562376 990100 668584 990128
rect 562376 990088 562382 990100
rect 668578 990088 668584 990100
rect 668636 990088 668642 990140
rect 563698 987368 563704 987420
rect 563756 987408 563762 987420
rect 608778 987408 608784 987420
rect 563756 987380 608784 987408
rect 563756 987368 563762 987380
rect 608778 987368 608784 987380
rect 608836 987368 608842 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 204898 986660 204904 986672
rect 203208 986632 204904 986660
rect 203208 986620 203214 986632
rect 204898 986620 204904 986632
rect 204956 986620 204962 986672
rect 89622 986076 89628 986128
rect 89680 986116 89686 986128
rect 111794 986116 111800 986128
rect 89680 986088 111800 986116
rect 89680 986076 89686 986088
rect 111794 986076 111800 986088
rect 111852 986076 111858 986128
rect 438118 986076 438124 986128
rect 438176 986116 438182 986128
rect 462774 986116 462780 986128
rect 438176 986088 462780 986116
rect 438176 986076 438182 986088
rect 462774 986076 462780 986088
rect 462832 986076 462838 986128
rect 515398 986076 515404 986128
rect 515456 986116 515462 986128
rect 527634 986116 527640 986128
rect 515456 986088 527640 986116
rect 515456 986076 515462 986088
rect 527634 986076 527640 986088
rect 527692 986076 527698 986128
rect 566458 986076 566464 986128
rect 566516 986116 566522 986128
rect 592494 986116 592500 986128
rect 566516 986088 592500 986116
rect 566516 986076 566522 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 370498 985940 370504 985992
rect 370556 985980 370562 985992
rect 397822 985980 397828 985992
rect 370556 985952 397828 985980
rect 370556 985940 370562 985952
rect 397822 985940 397828 985952
rect 397880 985940 397886 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 495158 985980 495164 985992
rect 436796 985952 495164 985980
rect 436796 985940 436802 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 664438 975712 664444 975724
rect 651708 975684 664444 975712
rect 651708 975672 651714 975684
rect 664438 975672 664444 975684
rect 664496 975672 664502 975724
rect 46198 961868 46204 961920
rect 46256 961908 46262 961920
rect 62114 961908 62120 961920
rect 46256 961880 62120 961908
rect 46256 961868 46262 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952348 36544 952400
rect 36596 952388 36602 952400
rect 41690 952388 41696 952400
rect 36596 952360 41696 952388
rect 36596 952348 36602 952360
rect 41690 952348 41696 952360
rect 41748 952348 41754 952400
rect 33778 951464 33784 951516
rect 33836 951504 33842 951516
rect 41506 951504 41512 951516
rect 33836 951476 41512 951504
rect 33836 951464 33842 951476
rect 41506 951464 41512 951476
rect 41564 951464 41570 951516
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 663058 948104 663064 948116
rect 652260 948076 663064 948104
rect 652260 948064 652266 948076
rect 663058 948064 663064 948076
rect 663116 948064 663122 948116
rect 676030 947996 676036 948048
rect 676088 948036 676094 948048
rect 680998 948036 681004 948048
rect 676088 948008 681004 948036
rect 676088 947996 676094 948008
rect 680998 947996 681004 948008
rect 681056 947996 681062 948048
rect 45554 945956 45560 946008
rect 45612 945996 45618 946008
rect 62114 945996 62120 946008
rect 45612 945968 62120 945996
rect 45612 945956 45618 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 28718 945276 28724 945328
rect 28776 945316 28782 945328
rect 31754 945316 31760 945328
rect 28776 945288 31760 945316
rect 28776 945276 28782 945288
rect 31754 945276 31760 945288
rect 31812 945276 31818 945328
rect 35802 942556 35808 942608
rect 35860 942596 35866 942608
rect 41690 942596 41696 942608
rect 35860 942568 41696 942596
rect 35860 942556 35866 942568
rect 41690 942556 41696 942568
rect 41748 942556 41754 942608
rect 35802 941196 35808 941248
rect 35860 941236 35866 941248
rect 35860 941208 37274 941236
rect 35860 941196 35866 941208
rect 37246 941168 37274 941208
rect 41690 941168 41696 941180
rect 37246 941140 41696 941168
rect 41690 941128 41696 941140
rect 41748 941128 41754 941180
rect 35802 939768 35808 939820
rect 35860 939808 35866 939820
rect 41506 939808 41512 939820
rect 35860 939780 41512 939808
rect 35860 939768 35866 939780
rect 41506 939768 41512 939780
rect 41564 939768 41570 939820
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 661678 921856 661684 921868
rect 651524 921828 661684 921856
rect 651524 921816 651530 921828
rect 661678 921816 661684 921828
rect 661736 921816 661742 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 663058 909480 663064 909492
rect 652444 909452 663064 909480
rect 652444 909440 652450 909452
rect 663058 909440 663064 909452
rect 663116 909440 663122 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 671338 895676 671344 895688
rect 651524 895648 671344 895676
rect 651524 895636 651530 895648
rect 671338 895636 671344 895648
rect 671396 895636 671402 895688
rect 44082 892752 44088 892764
rect 42858 892724 44088 892752
rect 42858 892466 42886 892724
rect 44082 892712 44088 892724
rect 44140 892712 44146 892764
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43070 892202 43076 892254
rect 43128 892202 43134 892254
rect 43088 892058 43116 892202
rect 44082 891936 44088 891948
rect 43180 891908 44088 891936
rect 43180 891854 43208 891908
rect 44082 891896 44088 891908
rect 44140 891896 44146 891948
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 652386 855584 652392 855636
rect 652444 855624 652450 855636
rect 664438 855624 664444 855636
rect 652444 855596 664444 855624
rect 652444 855584 652450 855596
rect 664438 855584 664444 855596
rect 664496 855584 664502 855636
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817028 35808 817080
rect 35860 817068 35866 817080
rect 41690 817068 41696 817080
rect 35860 817040 41696 817068
rect 35860 817028 35866 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 41598 815640 41604 815652
rect 35860 815612 41604 815640
rect 35860 815600 35866 815612
rect 41598 815600 41604 815612
rect 41656 815600 41662 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 669958 815640 669964 815652
rect 651524 815612 669964 815640
rect 651524 815600 651530 815612
rect 669958 815600 669964 815612
rect 670016 815600 670022 815652
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 41414 814280 41420 814292
rect 35860 814252 41420 814280
rect 35860 814240 35866 814252
rect 41414 814240 41420 814252
rect 41472 814240 41478 814292
rect 41322 811588 41328 811640
rect 41380 811628 41386 811640
rect 41690 811628 41696 811640
rect 41380 811600 41696 811628
rect 41380 811588 41386 811600
rect 41690 811588 41696 811600
rect 41748 811588 41754 811640
rect 40770 808936 40776 808988
rect 40828 808976 40834 808988
rect 41598 808976 41604 808988
rect 40828 808948 41604 808976
rect 40828 808936 40834 808948
rect 41598 808936 41604 808948
rect 41656 808936 41662 808988
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 35158 802408 35164 802460
rect 35216 802448 35222 802460
rect 41690 802448 41696 802460
rect 35216 802420 41696 802448
rect 35216 802408 35222 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 35894 802272 35900 802324
rect 35952 802312 35958 802324
rect 41690 802312 41696 802324
rect 35952 802284 41696 802312
rect 35952 802272 35958 802284
rect 41690 802272 41696 802284
rect 41748 802272 41754 802324
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 668762 775588 668768 775600
rect 651524 775560 668768 775588
rect 651524 775548 651530 775560
rect 668762 775548 668768 775560
rect 668820 775548 668826 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 41322 768992 41328 769004
rect 35860 768964 41328 768992
rect 35860 768952 35866 768964
rect 41322 768952 41328 768964
rect 41380 768952 41386 769004
rect 35618 768816 35624 768868
rect 35676 768856 35682 768868
rect 41690 768856 41696 768868
rect 35676 768828 41696 768856
rect 35676 768816 35682 768828
rect 41690 768816 41696 768828
rect 41748 768816 41754 768868
rect 35434 768680 35440 768732
rect 35492 768720 35498 768732
rect 40034 768720 40040 768732
rect 35492 768692 40040 768720
rect 35492 768680 35498 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 35526 767320 35532 767372
rect 35584 767360 35590 767372
rect 37918 767360 37924 767372
rect 35584 767332 37924 767360
rect 35584 767320 35590 767332
rect 37918 767320 37924 767332
rect 37976 767320 37982 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 37090 763240 37096 763292
rect 37148 763280 37154 763292
rect 39298 763280 39304 763292
rect 37148 763252 39304 763280
rect 37148 763240 37154 763252
rect 39298 763240 39304 763252
rect 39356 763240 39362 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 37918 759024 37924 759076
rect 37976 759064 37982 759076
rect 39482 759064 39488 759076
rect 37976 759036 39488 759064
rect 37976 759024 37982 759036
rect 39482 759024 39488 759036
rect 39540 759024 39546 759076
rect 35158 758412 35164 758464
rect 35216 758452 35222 758464
rect 41690 758452 41696 758464
rect 35216 758424 41696 758452
rect 35216 758412 35222 758424
rect 41690 758412 41696 758424
rect 41748 758412 41754 758464
rect 42058 758344 42064 758396
rect 42116 758344 42122 758396
rect 31018 758208 31024 758260
rect 31076 758248 31082 758260
rect 31076 758220 38654 758248
rect 31076 758208 31082 758220
rect 38626 758180 38654 758220
rect 40678 758180 40684 758192
rect 38626 758152 40684 758180
rect 40678 758140 40684 758152
rect 40736 758140 40742 758192
rect 42076 758056 42104 758344
rect 42058 758004 42064 758056
rect 42116 758004 42122 758056
rect 39298 757596 39304 757648
rect 39356 757636 39362 757648
rect 41690 757636 41696 757648
rect 39356 757608 41696 757636
rect 39356 757596 39362 757608
rect 41690 757596 41696 757608
rect 41748 757596 41754 757648
rect 676030 757120 676036 757172
rect 676088 757160 676094 757172
rect 683114 757160 683120 757172
rect 676088 757132 683120 757160
rect 676088 757120 676094 757132
rect 683114 757120 683120 757132
rect 683172 757120 683178 757172
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 652570 735564 652576 735616
rect 652628 735604 652634 735616
rect 671338 735604 671344 735616
rect 652628 735576 671344 735604
rect 652628 735564 652634 735576
rect 671338 735564 671344 735576
rect 671396 735564 671402 735616
rect 673546 732096 673552 732148
rect 673604 732136 673610 732148
rect 674006 732136 674012 732148
rect 673604 732108 674012 732136
rect 673604 732096 673610 732108
rect 674006 732096 674012 732108
rect 674064 732096 674070 732148
rect 35802 730192 35808 730244
rect 35860 730232 35866 730244
rect 41690 730232 41696 730244
rect 35860 730204 41696 730232
rect 35860 730192 35866 730204
rect 41690 730192 41696 730204
rect 41748 730192 41754 730244
rect 35618 730056 35624 730108
rect 35676 730096 35682 730108
rect 41690 730096 41696 730108
rect 35676 730068 41696 730096
rect 35676 730056 35682 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 674208 728640 674406 728668
rect 673822 728560 673828 728612
rect 673880 728600 673886 728612
rect 674208 728600 674236 728640
rect 673880 728572 674236 728600
rect 673880 728560 673886 728572
rect 673362 728424 673368 728476
rect 673420 728464 673426 728476
rect 673420 728436 674268 728464
rect 673420 728424 673426 728436
rect 674150 728136 674202 728142
rect 672994 728084 673000 728136
rect 673052 728124 673058 728136
rect 673052 728096 674058 728124
rect 673052 728084 673058 728096
rect 674150 728078 674202 728084
rect 41322 725908 41328 725960
rect 41380 725948 41386 725960
rect 41690 725948 41696 725960
rect 41380 725920 41696 725948
rect 41380 725908 41386 725920
rect 41690 725908 41696 725920
rect 41748 725908 41754 725960
rect 41322 724480 41328 724532
rect 41380 724520 41386 724532
rect 41690 724520 41696 724532
rect 41380 724492 41696 724520
rect 41380 724480 41386 724492
rect 41690 724480 41696 724492
rect 41748 724480 41754 724532
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 31018 716796 31024 716848
rect 31076 716836 31082 716848
rect 41598 716836 41604 716848
rect 31076 716808 41604 716836
rect 31076 716796 31082 716808
rect 41598 716796 41604 716808
rect 41656 716796 41662 716848
rect 33778 715640 33784 715692
rect 33836 715680 33842 715692
rect 41506 715680 41512 715692
rect 33836 715652 41512 715680
rect 33836 715640 33842 715652
rect 41506 715640 41512 715652
rect 41564 715640 41570 715692
rect 33042 715504 33048 715556
rect 33100 715544 33106 715556
rect 41690 715544 41696 715556
rect 33100 715516 41696 715544
rect 33100 715504 33106 715516
rect 41690 715504 41696 715516
rect 41748 715504 41754 715556
rect 36538 715368 36544 715420
rect 36596 715408 36602 715420
rect 36596 715380 41414 715408
rect 36596 715368 36602 715380
rect 41386 715068 41414 715380
rect 41598 715068 41604 715080
rect 41386 715040 41604 715068
rect 41598 715028 41604 715040
rect 41656 715028 41662 715080
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 652570 709316 652576 709368
rect 652628 709356 652634 709368
rect 664438 709356 664444 709368
rect 652628 709328 664444 709356
rect 652628 709316 652634 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 672442 707208 672448 707260
rect 672500 707248 672506 707260
rect 672994 707248 673000 707260
rect 672500 707220 673000 707248
rect 672500 707208 672506 707220
rect 672994 707208 673000 707220
rect 673052 707208 673058 707260
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 652386 696940 652392 696992
rect 652444 696980 652450 696992
rect 661678 696980 661684 696992
rect 652444 696952 661684 696980
rect 652444 696940 652450 696952
rect 661678 696940 661684 696952
rect 661736 696940 661742 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 35802 687216 35808 687268
rect 35860 687256 35866 687268
rect 41690 687256 41696 687268
rect 35860 687228 41696 687256
rect 35860 687216 35866 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 35802 683136 35808 683188
rect 35860 683176 35866 683188
rect 41506 683176 41512 683188
rect 35860 683148 41512 683176
rect 35860 683136 35866 683148
rect 41506 683136 41512 683148
rect 41564 683136 41570 683188
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35802 681708 35808 681760
rect 35860 681748 35866 681760
rect 41322 681748 41328 681760
rect 35860 681720 41328 681748
rect 35860 681708 35866 681720
rect 41322 681708 41328 681720
rect 41380 681708 41386 681760
rect 35434 681028 35440 681080
rect 35492 681068 35498 681080
rect 41598 681068 41604 681080
rect 35492 681040 41604 681068
rect 35492 681028 35498 681040
rect 41598 681028 41604 681040
rect 41656 681028 41662 681080
rect 35802 680620 35808 680672
rect 35860 680660 35866 680672
rect 37918 680660 37924 680672
rect 35860 680632 37924 680660
rect 35860 680620 35866 680632
rect 37918 680620 37924 680632
rect 37976 680620 37982 680672
rect 35618 680348 35624 680400
rect 35676 680388 35682 680400
rect 36538 680388 36544 680400
rect 35676 680360 36544 680388
rect 35676 680348 35682 680360
rect 36538 680348 36544 680360
rect 36596 680348 36602 680400
rect 51718 674840 51724 674892
rect 51776 674880 51782 674892
rect 62114 674880 62120 674892
rect 51776 674852 62120 674880
rect 51776 674840 51782 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 40494 672772 40500 672784
rect 35216 672744 40500 672772
rect 35216 672732 35222 672744
rect 40494 672732 40500 672744
rect 40552 672732 40558 672784
rect 36538 672052 36544 672104
rect 36596 672092 36602 672104
rect 41598 672092 41604 672104
rect 36596 672064 41604 672092
rect 36596 672052 36602 672064
rect 41598 672052 41604 672064
rect 41656 672052 41662 672104
rect 39942 671440 39948 671492
rect 40000 671480 40006 671492
rect 41690 671480 41696 671492
rect 40000 671452 41696 671480
rect 40000 671440 40006 671452
rect 41690 671440 41696 671452
rect 41748 671440 41754 671492
rect 651466 669332 651472 669384
rect 651524 669372 651530 669384
rect 661862 669372 661868 669384
rect 651524 669344 661868 669372
rect 651524 669332 651530 669344
rect 661862 669332 661868 669344
rect 661920 669332 661926 669384
rect 671062 666204 671068 666256
rect 671120 666244 671126 666256
rect 673362 666244 673368 666256
rect 671120 666216 673368 666244
rect 671120 666204 671126 666216
rect 673362 666204 673368 666216
rect 673420 666204 673426 666256
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651466 656888 651472 656940
rect 651524 656928 651530 656940
rect 670142 656928 670148 656940
rect 651524 656900 670148 656928
rect 651524 656888 651530 656900
rect 670142 656888 670148 656900
rect 670200 656888 670206 656940
rect 54478 647844 54484 647896
rect 54536 647884 54542 647896
rect 62114 647884 62120 647896
rect 54536 647856 62120 647884
rect 54536 647844 54542 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 41690 639112 41696 639124
rect 35866 639084 41696 639112
rect 41690 639072 41696 639084
rect 41748 639072 41754 639124
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 40034 638976 40040 638988
rect 35860 638948 40040 638976
rect 35860 638936 35866 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 41322 637616 41328 637628
rect 35860 637588 41328 637616
rect 35860 637576 35866 637588
rect 41322 637576 41328 637588
rect 41380 637576 41386 637628
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651466 629280 651472 629332
rect 651524 629320 651530 629332
rect 667198 629320 667204 629332
rect 651524 629292 667204 629320
rect 651524 629280 651530 629292
rect 667198 629280 667204 629292
rect 667256 629280 667262 629332
rect 675846 626560 675852 626612
rect 675904 626600 675910 626612
rect 676490 626600 676496 626612
rect 675904 626572 676496 626600
rect 675904 626560 675910 626572
rect 676490 626560 676496 626572
rect 676548 626560 676554 626612
rect 48958 623772 48964 623824
rect 49016 623812 49022 623824
rect 62114 623812 62120 623824
rect 49016 623784 62120 623812
rect 49016 623772 49022 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 43530 612932 43536 612944
rect 43286 612904 43536 612932
rect 43530 612892 43536 612904
rect 43588 612892 43594 612944
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43714 612524 43720 612536
rect 43516 612496 43720 612524
rect 43714 612484 43720 612496
rect 43772 612484 43778 612536
rect 46382 612388 46388 612400
rect 43732 612360 46388 612388
rect 43582 612332 43634 612338
rect 43582 612274 43634 612280
rect 43732 612102 43760 612360
rect 46382 612348 46388 612360
rect 46440 612348 46446 612400
rect 671890 612320 671896 612332
rect 671448 612292 671896 612320
rect 671448 612196 671476 612292
rect 671890 612280 671896 612292
rect 671948 612280 671954 612332
rect 671430 612144 671436 612196
rect 671488 612144 671494 612196
rect 45554 611912 45560 611924
rect 43838 611884 45560 611912
rect 45554 611872 45560 611884
rect 45612 611872 45618 611924
rect 46934 611708 46940 611720
rect 43957 611680 46940 611708
rect 46934 611668 46940 611680
rect 46992 611668 46998 611720
rect 44042 611516 44094 611522
rect 44042 611458 44094 611464
rect 45738 611300 45744 611312
rect 44181 611272 45744 611300
rect 45738 611260 45744 611272
rect 45796 611260 45802 611312
rect 47210 611096 47216 611108
rect 44298 611068 47216 611096
rect 47210 611056 47216 611068
rect 47268 611056 47274 611108
rect 44818 610920 44824 610972
rect 44876 610920 44882 610972
rect 44379 610904 44431 610910
rect 44379 610846 44431 610852
rect 44836 610688 44864 610920
rect 44528 610660 44864 610688
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 664622 603140 664628 603152
rect 651524 603112 664628 603140
rect 651524 603100 651530 603112
rect 664622 603100 664628 603112
rect 664680 603100 664686 603152
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 41230 594668 41236 594720
rect 41288 594708 41294 594720
rect 41506 594708 41512 594720
rect 41288 594680 41512 594708
rect 41288 594668 41294 594680
rect 41506 594668 41512 594680
rect 41564 594668 41570 594720
rect 41322 593376 41328 593428
rect 41380 593416 41386 593428
rect 41690 593416 41696 593428
rect 41380 593388 41696 593416
rect 41380 593376 41386 593388
rect 41690 593376 41696 593388
rect 41748 593376 41754 593428
rect 40494 592356 40500 592408
rect 40552 592396 40558 592408
rect 41690 592396 41696 592408
rect 40552 592368 41696 592396
rect 40552 592356 40558 592368
rect 41690 592356 41696 592368
rect 41748 592356 41754 592408
rect 41046 592016 41052 592068
rect 41104 592056 41110 592068
rect 41690 592056 41696 592068
rect 41104 592028 41696 592056
rect 41104 592016 41110 592028
rect 41690 592016 41696 592028
rect 41748 592016 41754 592068
rect 675938 591336 675944 591388
rect 675996 591376 676002 591388
rect 679618 591376 679624 591388
rect 675996 591348 679624 591376
rect 675996 591336 676002 591348
rect 679618 591336 679624 591348
rect 679676 591336 679682 591388
rect 676122 591200 676128 591252
rect 676180 591240 676186 591252
rect 682378 591240 682384 591252
rect 676180 591212 682384 591240
rect 676180 591200 676186 591212
rect 682378 591200 682384 591212
rect 682436 591200 682442 591252
rect 651466 590656 651472 590708
rect 651524 590696 651530 590708
rect 662046 590696 662052 590708
rect 651524 590668 662052 590696
rect 651524 590656 651530 590668
rect 662046 590656 662052 590668
rect 662104 590656 662110 590708
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 41690 585936 41696 585948
rect 35216 585908 41696 585936
rect 35216 585896 35222 585908
rect 41690 585896 41696 585908
rect 41748 585896 41754 585948
rect 32398 585760 32404 585812
rect 32456 585800 32462 585812
rect 41690 585800 41696 585812
rect 32456 585772 41696 585800
rect 32456 585760 32462 585772
rect 41690 585760 41696 585772
rect 41748 585760 41754 585812
rect 36538 585148 36544 585200
rect 36596 585188 36602 585200
rect 41414 585188 41420 585200
rect 36596 585160 41420 585188
rect 36596 585148 36602 585160
rect 41414 585148 41420 585160
rect 41472 585148 41478 585200
rect 51718 583720 51724 583772
rect 51776 583760 51782 583772
rect 62114 583760 62120 583772
rect 51776 583732 62120 583760
rect 51776 583720 51782 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 671062 578008 671068 578060
rect 671120 578048 671126 578060
rect 671706 578048 671712 578060
rect 671120 578020 671712 578048
rect 671120 578008 671126 578020
rect 671706 578008 671712 578020
rect 671764 578008 671770 578060
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 666002 576892 666008 576904
rect 651524 576864 666008 576892
rect 651524 576852 651530 576864
rect 666002 576852 666008 576864
rect 666060 576852 666066 576904
rect 672258 571956 672264 572008
rect 672316 571996 672322 572008
rect 672810 571996 672816 572008
rect 672316 571968 672816 571996
rect 672316 571956 672322 571968
rect 672810 571956 672816 571968
rect 672868 571956 672874 572008
rect 679618 571276 679624 571328
rect 679676 571316 679682 571328
rect 683114 571316 683120 571328
rect 679676 571288 683120 571316
rect 679676 571276 679682 571288
rect 683114 571276 683120 571288
rect 683172 571276 683178 571328
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 41506 557580 41512 557592
rect 35860 557552 41512 557580
rect 35860 557540 35866 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 41690 554792 41696 554804
rect 35860 554764 41696 554792
rect 35860 554752 35866 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 35802 553528 35808 553580
rect 35860 553568 35866 553580
rect 41690 553568 41696 553580
rect 35860 553540 41696 553568
rect 35860 553528 35866 553540
rect 41690 553528 41696 553540
rect 41748 553528 41754 553580
rect 35618 553392 35624 553444
rect 35676 553432 35682 553444
rect 41322 553432 41328 553444
rect 35676 553404 41328 553432
rect 35676 553392 35682 553404
rect 41322 553392 41328 553404
rect 41380 553392 41386 553444
rect 41322 552032 41328 552084
rect 41380 552072 41386 552084
rect 41598 552072 41604 552084
rect 41380 552044 41604 552072
rect 41380 552032 41386 552044
rect 41598 552032 41604 552044
rect 41656 552032 41662 552084
rect 41322 550740 41328 550792
rect 41380 550780 41386 550792
rect 41598 550780 41604 550792
rect 41380 550752 41604 550780
rect 41380 550740 41386 550752
rect 41598 550740 41604 550752
rect 41656 550740 41662 550792
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 675846 547544 675852 547596
rect 675904 547584 675910 547596
rect 678238 547584 678244 547596
rect 675904 547556 678244 547584
rect 675904 547544 675910 547556
rect 678238 547544 678244 547556
rect 678296 547544 678302 547596
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 37090 547448 37096 547460
rect 31812 547420 37096 547448
rect 31812 547408 31818 547420
rect 37090 547408 37096 547420
rect 37148 547408 37154 547460
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 41506 543028 41512 543040
rect 33836 543000 41512 543028
rect 33836 542988 33842 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 37090 542308 37096 542360
rect 37148 542348 37154 542360
rect 41690 542348 41696 542360
rect 37148 542320 41696 542348
rect 37148 542308 37154 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669958 536840 669964 536852
rect 651524 536812 669964 536840
rect 651524 536800 651530 536812
rect 669958 536800 669964 536812
rect 670016 536800 670022 536852
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 672258 531972 672264 532024
rect 672316 532012 672322 532024
rect 672626 532012 672632 532024
rect 672316 531984 672632 532012
rect 672316 531972 672322 531984
rect 672626 531972 672632 531984
rect 672684 531972 672690 532024
rect 673178 530408 673184 530460
rect 673236 530448 673242 530460
rect 673822 530448 673828 530460
rect 673236 530420 673828 530448
rect 673236 530408 673242 530420
rect 673822 530408 673828 530420
rect 673880 530408 673886 530460
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 675846 518780 675852 518832
rect 675904 518820 675910 518832
rect 677870 518820 677876 518832
rect 675904 518792 677876 518820
rect 675904 518780 675910 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675846 503616 675852 503668
rect 675904 503656 675910 503668
rect 679618 503656 679624 503668
rect 675904 503628 679624 503656
rect 675904 503616 675910 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 676030 503480 676036 503532
rect 676088 503520 676094 503532
rect 682378 503520 682384 503532
rect 676088 503492 682384 503520
rect 676088 503480 676094 503492
rect 682378 503480 682384 503492
rect 682436 503480 682442 503532
rect 675846 502324 675852 502376
rect 675904 502364 675910 502376
rect 676858 502364 676864 502376
rect 675904 502336 676864 502364
rect 675904 502324 675910 502336
rect 676858 502324 676864 502336
rect 676916 502324 676922 502376
rect 676030 500896 676036 500948
rect 676088 500936 676094 500948
rect 680998 500936 681004 500948
rect 676088 500908 681004 500936
rect 676088 500896 676094 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 652570 494708 652576 494760
rect 652628 494748 652634 494760
rect 665818 494748 665824 494760
rect 652628 494720 665824 494748
rect 652628 494708 652634 494720
rect 665818 494708 665824 494720
rect 665876 494708 665882 494760
rect 676030 492668 676036 492720
rect 676088 492708 676094 492720
rect 683390 492708 683396 492720
rect 676088 492680 683396 492708
rect 676088 492668 676094 492680
rect 683390 492668 683396 492680
rect 683448 492668 683454 492720
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 673362 488656 673368 488708
rect 673420 488656 673426 488708
rect 673380 488300 673408 488656
rect 673362 488248 673368 488300
rect 673420 488248 673426 488300
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 668762 484412 668768 484424
rect 654106 484384 668768 484412
rect 668762 484372 668768 484384
rect 668820 484372 668826 484424
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 663058 470608 663064 470620
rect 651524 470580 663064 470608
rect 651524 470568 651530 470580
rect 663058 470568 663064 470580
rect 663116 470568 663122 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 667198 456804 667204 456816
rect 652444 456776 667204 456804
rect 652444 456764 652450 456776
rect 667198 456764 667204 456776
rect 667256 456764 667262 456816
rect 673948 456204 674000 456210
rect 673948 456146 674000 456152
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673454 455812 673460 455864
rect 673512 455852 673518 455864
rect 673512 455824 673762 455852
rect 673512 455812 673518 455824
rect 673598 455660 673650 455666
rect 673598 455602 673650 455608
rect 673506 455388 673558 455394
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673388 455126 673440 455132
rect 671982 455064 671988 455116
rect 672040 455104 672046 455116
rect 672040 455076 673316 455104
rect 672040 455064 672046 455076
rect 673288 455022 673316 455076
rect 673164 454844 673216 454850
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673046 454582 673098 454588
rect 672954 454368 673006 454374
rect 672954 454310 673006 454316
rect 672816 454096 672868 454102
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672816 454038 672868 454044
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 671338 430624 671344 430636
rect 651524 430596 671344 430624
rect 651524 430584 651530 430596
rect 671338 430584 671344 430596
rect 671396 430584 671402 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41322 423648 41328 423700
rect 41380 423688 41386 423700
rect 41690 423688 41696 423700
rect 41380 423660 41696 423688
rect 41380 423648 41386 423660
rect 41690 423648 41696 423660
rect 41748 423648 41754 423700
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 661678 416820 661684 416832
rect 651892 416792 661684 416820
rect 651892 416780 651898 416792
rect 661678 416780 661684 416792
rect 661736 416780 661742 416832
rect 49142 415420 49148 415472
rect 49200 415460 49206 415472
rect 62114 415460 62120 415472
rect 49200 415432 62120 415460
rect 49200 415420 49206 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 36538 415352 36544 415404
rect 36596 415392 36602 415404
rect 41690 415392 41696 415404
rect 36596 415364 41696 415392
rect 36596 415352 36602 415364
rect 41690 415352 41696 415364
rect 41748 415352 41754 415404
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 41138 387064 41144 387116
rect 41196 387104 41202 387116
rect 41690 387104 41696 387116
rect 41196 387076 41696 387104
rect 41196 387064 41202 387076
rect 41690 387064 41696 387076
rect 41748 387064 41754 387116
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41506 382412 41512 382424
rect 41380 382384 41512 382412
rect 41380 382372 41386 382384
rect 41506 382372 41512 382384
rect 41564 382372 41570 382424
rect 35802 379652 35808 379704
rect 35860 379692 35866 379704
rect 41690 379692 41696 379704
rect 35860 379664 41696 379692
rect 35860 379652 35866 379664
rect 41690 379652 41696 379664
rect 41748 379652 41754 379704
rect 40218 378496 40224 378548
rect 40276 378536 40282 378548
rect 41690 378536 41696 378548
rect 40276 378508 41696 378536
rect 40276 378496 40282 378508
rect 41690 378496 41696 378508
rect 41748 378496 41754 378548
rect 35802 375368 35808 375420
rect 35860 375408 35866 375420
rect 41690 375408 41696 375420
rect 35860 375380 41696 375408
rect 35860 375368 35866 375380
rect 41690 375368 41696 375380
rect 41748 375368 41754 375420
rect 51718 375368 51724 375420
rect 51776 375408 51782 375420
rect 62114 375408 62120 375420
rect 51776 375380 62120 375408
rect 51776 375368 51782 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 37918 373260 37924 373312
rect 37976 373300 37982 373312
rect 41690 373300 41696 373312
rect 37976 373272 41696 373300
rect 37976 373260 37982 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 651650 364352 651656 364404
rect 651708 364392 651714 364404
rect 663242 364392 663248 364404
rect 651708 364364 663248 364392
rect 651708 364352 651714 364364
rect 663242 364352 663248 364364
rect 663300 364352 663306 364404
rect 46382 362924 46388 362976
rect 46440 362964 46446 362976
rect 62114 362964 62120 362976
rect 46440 362936 62120 362964
rect 46440 362924 46446 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 45002 355784 45008 355836
rect 45060 355824 45066 355836
rect 45646 355824 45652 355836
rect 45060 355796 45652 355824
rect 45060 355784 45066 355796
rect 45646 355784 45652 355796
rect 45704 355784 45710 355836
rect 44634 355648 44640 355700
rect 44692 355688 44698 355700
rect 44692 355660 45048 355688
rect 44692 355648 44698 355660
rect 44569 354832 44575 354884
rect 44627 354872 44633 354884
rect 44627 354844 44839 354872
rect 44627 354832 44633 354844
rect 44575 354680 44627 354686
rect 44575 354622 44627 354628
rect 44811 354600 44839 354844
rect 45020 354600 45048 355660
rect 44811 354572 44956 354600
rect 45020 354572 45063 354600
rect 44793 354424 44799 354476
rect 44851 354424 44857 354476
rect 44686 354340 44738 354346
rect 44811 354314 44839 354424
rect 44686 354282 44738 354288
rect 44928 354110 44956 354572
rect 45035 353906 45063 354572
rect 45646 354056 45652 354068
rect 45158 354028 45652 354056
rect 45158 353702 45186 354028
rect 45646 354016 45652 354028
rect 45704 354016 45710 354068
rect 45922 353784 45928 353796
rect 45250 353756 45928 353784
rect 45250 353498 45278 353756
rect 45922 353744 45928 353756
rect 45980 353744 45986 353796
rect 45554 353240 45560 353252
rect 45385 353212 45560 353240
rect 45554 353200 45560 353212
rect 45612 353200 45618 353252
rect 651466 350548 651472 350600
rect 651524 350588 651530 350600
rect 667382 350588 667388 350600
rect 651524 350560 667388 350588
rect 651524 350548 651530 350560
rect 667382 350548 667388 350560
rect 667440 350548 667446 350600
rect 28902 345040 28908 345092
rect 28960 345080 28966 345092
rect 38286 345080 38292 345092
rect 28960 345052 38292 345080
rect 28960 345040 28966 345052
rect 38286 345040 38292 345052
rect 38344 345040 38350 345092
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 37918 339504 37924 339516
rect 35860 339476 37924 339504
rect 35860 339464 35866 339476
rect 37918 339464 37924 339476
rect 37976 339464 37982 339516
rect 35802 338104 35808 338156
rect 35860 338144 35866 338156
rect 36538 338144 36544 338156
rect 35860 338116 36544 338144
rect 35860 338104 35866 338116
rect 36538 338104 36544 338116
rect 36596 338104 36602 338156
rect 651466 338104 651472 338156
rect 651524 338144 651530 338156
rect 666186 338144 666192 338156
rect 651524 338116 666192 338144
rect 651524 338104 651530 338116
rect 666186 338104 666192 338116
rect 666244 338104 666250 338156
rect 50338 336744 50344 336796
rect 50396 336784 50402 336796
rect 62114 336784 62120 336796
rect 50396 336756 62120 336784
rect 50396 336744 50402 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 667750 324340 667756 324352
rect 651524 324312 667756 324340
rect 651524 324300 651530 324312
rect 667750 324300 667756 324312
rect 667808 324300 667814 324352
rect 54478 310496 54484 310548
rect 54536 310536 54542 310548
rect 62114 310536 62120 310548
rect 54536 310508 62120 310536
rect 54536 310496 54542 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667198 310536 667204 310548
rect 651524 310508 667204 310536
rect 651524 310496 651530 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675938 298052 675944 298104
rect 675996 298092 676002 298104
rect 678974 298092 678980 298104
rect 675996 298064 678980 298092
rect 675996 298052 676002 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676122 297848 676128 297900
rect 676180 297888 676186 297900
rect 680998 297888 681004 297900
rect 676180 297860 681004 297888
rect 676180 297848 676186 297860
rect 680998 297848 681004 297860
rect 681056 297848 681062 297900
rect 41322 285064 41328 285116
rect 41380 285104 41386 285116
rect 41690 285104 41696 285116
rect 41380 285076 41696 285104
rect 41380 285064 41386 285076
rect 41690 285064 41696 285076
rect 41748 285064 41754 285116
rect 32398 284928 32404 284980
rect 32456 284968 32462 284980
rect 41690 284968 41696 284980
rect 32456 284940 41696 284968
rect 32456 284928 32462 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667566 284356 667572 284368
rect 651524 284328 667572 284356
rect 651524 284316 651530 284328
rect 667566 284316 667572 284328
rect 667624 284316 667630 284368
rect 522942 276224 522948 276276
rect 523000 276264 523006 276276
rect 526898 276264 526904 276276
rect 523000 276236 526904 276264
rect 523000 276224 523006 276236
rect 526898 276224 526904 276236
rect 526956 276224 526962 276276
rect 524874 276128 524880 276140
rect 524156 276100 524880 276128
rect 524156 276060 524184 276100
rect 524874 276088 524880 276100
rect 524932 276088 524938 276140
rect 524064 276032 524184 276060
rect 88334 275952 88340 276004
rect 88392 275992 88398 276004
rect 143350 275992 143356 276004
rect 88392 275964 143356 275992
rect 88392 275952 88398 275964
rect 143350 275952 143356 275964
rect 143408 275952 143414 276004
rect 156874 275952 156880 276004
rect 156932 275992 156938 276004
rect 193858 275992 193864 276004
rect 156932 275964 193864 275992
rect 156932 275952 156938 275964
rect 193858 275952 193864 275964
rect 193916 275952 193922 276004
rect 201770 275952 201776 276004
rect 201828 275992 201834 276004
rect 222102 275992 222108 276004
rect 201828 275964 222108 275992
rect 201828 275952 201834 275964
rect 222102 275952 222108 275964
rect 222160 275952 222166 276004
rect 389174 275952 389180 276004
rect 389232 275992 389238 276004
rect 393314 275992 393320 276004
rect 389232 275964 393320 275992
rect 389232 275952 389238 275964
rect 393314 275952 393320 275964
rect 393372 275952 393378 276004
rect 400582 275952 400588 276004
rect 400640 275992 400646 276004
rect 415762 275992 415768 276004
rect 400640 275964 415768 275992
rect 400640 275952 400646 275964
rect 415762 275952 415768 275964
rect 415820 275952 415826 276004
rect 427814 275952 427820 276004
rect 427872 275992 427878 276004
rect 442994 275992 443000 276004
rect 427872 275964 443000 275992
rect 427872 275952 427878 275964
rect 442994 275952 443000 275964
rect 443052 275952 443058 276004
rect 443730 275952 443736 276004
rect 443788 275992 443794 276004
rect 453574 275992 453580 276004
rect 443788 275964 453580 275992
rect 443788 275952 443794 275964
rect 453574 275952 453580 275964
rect 453632 275952 453638 276004
rect 456978 275952 456984 276004
rect 457036 275992 457042 276004
rect 486694 275992 486700 276004
rect 457036 275964 486700 275992
rect 457036 275952 457042 275964
rect 486694 275952 486700 275964
rect 486752 275952 486758 276004
rect 486878 275952 486884 276004
rect 486936 275992 486942 276004
rect 494698 275992 494704 276004
rect 486936 275964 494704 275992
rect 486936 275952 486942 275964
rect 494698 275952 494704 275964
rect 494756 275952 494762 276004
rect 495434 275952 495440 276004
rect 495492 275992 495498 276004
rect 504358 275992 504364 276004
rect 495492 275964 504364 275992
rect 495492 275952 495498 275964
rect 504358 275952 504364 275964
rect 504416 275952 504422 276004
rect 504910 275952 504916 276004
rect 504968 275992 504974 276004
rect 507026 275992 507032 276004
rect 504968 275964 507032 275992
rect 504968 275952 504974 275964
rect 507026 275952 507032 275964
rect 507084 275952 507090 276004
rect 508038 275952 508044 276004
rect 508096 275992 508102 276004
rect 514018 275992 514024 276004
rect 508096 275964 514024 275992
rect 508096 275952 508102 275964
rect 514018 275952 514024 275964
rect 514076 275952 514082 276004
rect 519814 275992 519820 276004
rect 514220 275964 519820 275992
rect 95418 275816 95424 275868
rect 95476 275856 95482 275868
rect 104802 275856 104808 275868
rect 95476 275828 104808 275856
rect 95476 275816 95482 275828
rect 104802 275816 104808 275828
rect 104860 275816 104866 275868
rect 113174 275816 113180 275868
rect 113232 275856 113238 275868
rect 169938 275856 169944 275868
rect 113232 275828 169944 275856
rect 113232 275816 113238 275828
rect 169938 275816 169944 275828
rect 169996 275816 170002 275868
rect 181714 275816 181720 275868
rect 181772 275856 181778 275868
rect 218882 275856 218888 275868
rect 181772 275828 218888 275856
rect 181772 275816 181778 275828
rect 218882 275816 218888 275828
rect 218940 275816 218946 275868
rect 393590 275816 393596 275868
rect 393648 275856 393654 275868
rect 412266 275856 412272 275868
rect 393648 275828 412272 275856
rect 393648 275816 393654 275828
rect 412266 275816 412272 275828
rect 412324 275816 412330 275868
rect 415302 275816 415308 275868
rect 415360 275856 415366 275868
rect 425238 275856 425244 275868
rect 415360 275828 425244 275856
rect 415360 275816 415366 275828
rect 425238 275816 425244 275828
rect 425296 275816 425302 275868
rect 432966 275816 432972 275868
rect 433024 275856 433030 275868
rect 487890 275856 487896 275868
rect 433024 275828 487896 275856
rect 433024 275816 433030 275828
rect 487890 275816 487896 275828
rect 487948 275816 487954 275868
rect 498194 275816 498200 275868
rect 498252 275856 498258 275868
rect 505646 275856 505652 275868
rect 498252 275828 505652 275856
rect 498252 275816 498258 275828
rect 505646 275816 505652 275828
rect 505704 275816 505710 275868
rect 507210 275816 507216 275868
rect 507268 275856 507274 275868
rect 512730 275856 512736 275868
rect 507268 275828 512736 275856
rect 507268 275816 507274 275828
rect 512730 275816 512736 275828
rect 512788 275816 512794 275868
rect 512914 275816 512920 275868
rect 512972 275856 512978 275868
rect 514220 275856 514248 275964
rect 519814 275952 519820 275964
rect 519872 275952 519878 276004
rect 519998 275952 520004 276004
rect 520056 275992 520062 276004
rect 524064 275992 524092 276032
rect 604914 275992 604920 276004
rect 520056 275964 524092 275992
rect 524248 275964 604920 275992
rect 520056 275952 520062 275964
rect 512972 275828 514248 275856
rect 512972 275816 512978 275828
rect 515490 275816 515496 275868
rect 515548 275856 515554 275868
rect 515548 275828 516456 275856
rect 515548 275816 515554 275828
rect 81250 275680 81256 275732
rect 81308 275720 81314 275732
rect 88978 275720 88984 275732
rect 81308 275692 88984 275720
rect 81308 275680 81314 275692
rect 88978 275680 88984 275692
rect 89036 275680 89042 275732
rect 103698 275680 103704 275732
rect 103756 275720 103762 275732
rect 160094 275720 160100 275732
rect 103756 275692 160100 275720
rect 103756 275680 103762 275692
rect 160094 275680 160100 275692
rect 160152 275680 160158 275732
rect 178126 275680 178132 275732
rect 178184 275720 178190 275732
rect 216858 275720 216864 275732
rect 178184 275692 216864 275720
rect 178184 275680 178190 275692
rect 216858 275680 216864 275692
rect 216916 275680 216922 275732
rect 299934 275680 299940 275732
rect 299992 275720 299998 275732
rect 300762 275720 300768 275732
rect 299992 275692 300768 275720
rect 299992 275680 299998 275692
rect 300762 275680 300768 275692
rect 300820 275680 300826 275732
rect 370498 275680 370504 275732
rect 370556 275720 370562 275732
rect 388622 275720 388628 275732
rect 370556 275692 388628 275720
rect 370556 275680 370562 275692
rect 388622 275680 388628 275692
rect 388680 275680 388686 275732
rect 410058 275680 410064 275732
rect 410116 275720 410122 275732
rect 428826 275720 428832 275732
rect 410116 275692 428832 275720
rect 410116 275680 410122 275692
rect 428826 275680 428832 275692
rect 428884 275680 428890 275732
rect 429194 275680 429200 275732
rect 429252 275720 429258 275732
rect 446490 275720 446496 275732
rect 429252 275692 446496 275720
rect 429252 275680 429258 275692
rect 446490 275680 446496 275692
rect 446548 275680 446554 275732
rect 502058 275720 502064 275732
rect 446692 275692 502064 275720
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86862 275584 86868 275596
rect 76524 275556 86868 275584
rect 76524 275544 76530 275556
rect 86862 275544 86868 275556
rect 86920 275544 86926 275596
rect 96614 275544 96620 275596
rect 96672 275584 96678 275596
rect 156598 275584 156604 275596
rect 96672 275556 156604 275584
rect 96672 275544 96678 275556
rect 156598 275544 156604 275556
rect 156656 275544 156662 275596
rect 163958 275544 163964 275596
rect 164016 275584 164022 275596
rect 202138 275584 202144 275596
rect 164016 275556 202144 275584
rect 164016 275544 164022 275556
rect 202138 275544 202144 275556
rect 202196 275544 202202 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 233878 275584 233884 275596
rect 221976 275556 233884 275584
rect 221976 275544 221982 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 236086 275544 236092 275596
rect 236144 275584 236150 275596
rect 251082 275584 251088 275596
rect 236144 275556 251088 275584
rect 236144 275544 236150 275556
rect 251082 275544 251088 275556
rect 251140 275544 251146 275596
rect 350718 275544 350724 275596
rect 350776 275584 350782 275596
rect 361390 275584 361396 275596
rect 350776 275556 361396 275584
rect 350776 275544 350782 275556
rect 361390 275544 361396 275556
rect 361448 275544 361454 275596
rect 362218 275544 362224 275596
rect 362276 275584 362282 275596
rect 385034 275584 385040 275596
rect 362276 275556 385040 275584
rect 362276 275544 362282 275556
rect 385034 275544 385040 275556
rect 385092 275544 385098 275596
rect 388162 275544 388168 275596
rect 388220 275584 388226 275596
rect 418154 275584 418160 275596
rect 388220 275556 418160 275584
rect 388220 275544 388226 275556
rect 418154 275544 418160 275556
rect 418212 275544 418218 275596
rect 418338 275544 418344 275596
rect 418396 275584 418402 275596
rect 435910 275584 435916 275596
rect 418396 275556 435916 275584
rect 418396 275544 418402 275556
rect 435910 275544 435916 275556
rect 435968 275544 435974 275596
rect 445754 275544 445760 275596
rect 445812 275584 445818 275596
rect 446692 275584 446720 275692
rect 502058 275680 502064 275692
rect 502116 275680 502122 275732
rect 502242 275680 502248 275732
rect 502300 275720 502306 275732
rect 509142 275720 509148 275732
rect 502300 275692 509148 275720
rect 502300 275680 502306 275692
rect 509142 275680 509148 275692
rect 509200 275680 509206 275732
rect 512178 275680 512184 275732
rect 512236 275720 512242 275732
rect 516226 275720 516232 275732
rect 512236 275692 516232 275720
rect 512236 275680 512242 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 516428 275720 516456 275828
rect 516778 275816 516784 275868
rect 516836 275856 516842 275868
rect 524248 275856 524276 275964
rect 604914 275952 604920 275964
rect 604972 275952 604978 276004
rect 516836 275828 524276 275856
rect 516836 275816 516842 275828
rect 524874 275816 524880 275868
rect 524932 275856 524938 275868
rect 611998 275856 612004 275868
rect 524932 275828 612004 275856
rect 524932 275816 524938 275828
rect 611998 275816 612004 275828
rect 612056 275816 612062 275868
rect 519170 275720 519176 275732
rect 516428 275692 519176 275720
rect 519170 275680 519176 275692
rect 519228 275680 519234 275732
rect 519354 275680 519360 275732
rect 519412 275720 519418 275732
rect 519412 275692 524276 275720
rect 519412 275680 519418 275692
rect 445812 275556 446720 275584
rect 445812 275544 445818 275556
rect 449158 275544 449164 275596
rect 449216 275584 449222 275596
rect 501782 275584 501788 275596
rect 449216 275556 501788 275584
rect 449216 275544 449222 275556
rect 501782 275544 501788 275556
rect 501840 275544 501846 275596
rect 519538 275584 519544 275596
rect 501984 275556 519544 275584
rect 85942 275408 85948 275460
rect 86000 275448 86006 275460
rect 146662 275448 146668 275460
rect 86000 275420 146668 275448
rect 86000 275408 86006 275420
rect 146662 275408 146668 275420
rect 146720 275408 146726 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 167730 275448 167736 275460
rect 160520 275420 167736 275448
rect 160520 275408 160526 275420
rect 167730 275408 167736 275420
rect 167788 275408 167794 275460
rect 171042 275408 171048 275460
rect 171100 275448 171106 275460
rect 210786 275448 210792 275460
rect 171100 275420 210792 275448
rect 171100 275408 171106 275420
rect 210786 275408 210792 275420
rect 210844 275408 210850 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 237466 275448 237472 275460
rect 218388 275420 237472 275448
rect 218388 275408 218394 275420
rect 237466 275408 237472 275420
rect 237524 275408 237530 275460
rect 244366 275408 244372 275460
rect 244424 275448 244430 275460
rect 254578 275448 254584 275460
rect 244424 275420 254584 275448
rect 244424 275408 244430 275420
rect 254578 275408 254584 275420
rect 254636 275408 254642 275460
rect 260926 275408 260932 275460
rect 260984 275448 260990 275460
rect 273530 275448 273536 275460
rect 260984 275420 273536 275448
rect 260984 275408 260990 275420
rect 273530 275408 273536 275420
rect 273588 275408 273594 275460
rect 273898 275408 273904 275460
rect 273956 275448 273962 275460
rect 282914 275448 282920 275460
rect 273956 275420 282920 275448
rect 273956 275408 273962 275420
rect 282914 275408 282920 275420
rect 282972 275408 282978 275460
rect 326430 275408 326436 275460
rect 326488 275448 326494 275460
rect 335354 275448 335360 275460
rect 326488 275420 335360 275448
rect 326488 275408 326494 275420
rect 335354 275408 335360 275420
rect 335412 275408 335418 275460
rect 341518 275408 341524 275460
rect 341576 275448 341582 275460
rect 354306 275448 354312 275460
rect 341576 275420 354312 275448
rect 341576 275408 341582 275420
rect 354306 275408 354312 275420
rect 354364 275408 354370 275460
rect 360194 275448 360200 275460
rect 354646 275420 360200 275448
rect 298738 275340 298744 275392
rect 298796 275380 298802 275392
rect 300026 275380 300032 275392
rect 298796 275352 300032 275380
rect 298796 275340 298802 275352
rect 300026 275340 300032 275352
rect 300084 275340 300090 275392
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 142706 275272 142712 275324
rect 142764 275312 142770 275324
rect 183462 275312 183468 275324
rect 142764 275284 183468 275312
rect 142764 275272 142770 275284
rect 183462 275272 183468 275284
rect 183520 275272 183526 275324
rect 186406 275272 186412 275324
rect 186464 275312 186470 275324
rect 187786 275312 187792 275324
rect 186464 275284 187792 275312
rect 186464 275272 186470 275284
rect 187786 275272 187792 275284
rect 187844 275272 187850 275324
rect 188798 275272 188804 275324
rect 188856 275312 188862 275324
rect 222838 275312 222844 275324
rect 188856 275284 222844 275312
rect 188856 275272 188862 275284
rect 222838 275272 222844 275284
rect 222896 275272 222902 275324
rect 225414 275272 225420 275324
rect 225472 275312 225478 275324
rect 245102 275312 245108 275324
rect 225472 275284 245108 275312
rect 225472 275272 225478 275284
rect 245102 275272 245108 275284
rect 245160 275272 245166 275324
rect 250254 275272 250260 275324
rect 250312 275312 250318 275324
rect 266354 275312 266360 275324
rect 250312 275284 266360 275312
rect 250312 275272 250318 275284
rect 266354 275272 266360 275284
rect 266412 275272 266418 275324
rect 266814 275272 266820 275324
rect 266872 275312 266878 275324
rect 276658 275312 276664 275324
rect 266872 275284 276664 275312
rect 266872 275272 266878 275284
rect 276658 275272 276664 275284
rect 276716 275272 276722 275324
rect 284570 275272 284576 275324
rect 284628 275312 284634 275324
rect 290090 275312 290096 275324
rect 284628 275284 290096 275312
rect 284628 275272 284634 275284
rect 290090 275272 290096 275284
rect 290148 275272 290154 275324
rect 329466 275272 329472 275324
rect 329524 275312 329530 275324
rect 338942 275312 338948 275324
rect 329524 275284 338948 275312
rect 329524 275272 329530 275284
rect 338942 275272 338948 275284
rect 339000 275272 339006 275324
rect 353110 275312 353116 275324
rect 344986 275284 353116 275312
rect 74074 275136 74080 275188
rect 74132 275176 74138 275188
rect 77202 275176 77208 275188
rect 74132 275148 77208 275176
rect 74132 275136 74138 275148
rect 77202 275136 77208 275148
rect 77260 275136 77266 275188
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 162118 275176 162124 275188
rect 110840 275148 162124 275176
rect 110840 275136 110846 275148
rect 162118 275136 162124 275148
rect 162176 275136 162182 275188
rect 338942 275136 338948 275188
rect 339000 275176 339006 275188
rect 344986 275176 345014 275284
rect 353110 275272 353116 275284
rect 353168 275272 353174 275324
rect 353938 275272 353944 275324
rect 353996 275312 354002 275324
rect 354646 275312 354674 275420
rect 360194 275408 360200 275420
rect 360252 275408 360258 275460
rect 363046 275408 363052 275460
rect 363104 275448 363110 275460
rect 367278 275448 367284 275460
rect 363104 275420 367284 275448
rect 363104 275408 363110 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 369118 275408 369124 275460
rect 369176 275448 369182 275460
rect 377950 275448 377956 275460
rect 369176 275420 377956 275448
rect 369176 275408 369182 275420
rect 377950 275408 377956 275420
rect 378008 275408 378014 275460
rect 381998 275408 382004 275460
rect 382056 275448 382062 275460
rect 414566 275448 414572 275460
rect 382056 275420 414572 275448
rect 382056 275408 382062 275420
rect 414566 275408 414572 275420
rect 414624 275408 414630 275460
rect 416406 275408 416412 275460
rect 416464 275448 416470 275460
rect 463050 275448 463056 275460
rect 416464 275420 463056 275448
rect 416464 275408 416470 275420
rect 463050 275408 463056 275420
rect 463108 275408 463114 275460
rect 467650 275408 467656 275460
rect 467708 275448 467714 275460
rect 501984 275448 502012 275556
rect 519538 275544 519544 275556
rect 519596 275544 519602 275596
rect 519722 275544 519728 275596
rect 519780 275584 519786 275596
rect 522942 275584 522948 275596
rect 519780 275556 522948 275584
rect 519780 275544 519786 275556
rect 522942 275544 522948 275556
rect 523000 275544 523006 275596
rect 524248 275584 524276 275692
rect 527358 275680 527364 275732
rect 527416 275720 527422 275732
rect 619082 275720 619088 275732
rect 527416 275692 619088 275720
rect 527416 275680 527422 275692
rect 619082 275680 619088 275692
rect 619140 275680 619146 275732
rect 530486 275584 530492 275596
rect 524248 275556 530492 275584
rect 530486 275544 530492 275556
rect 530544 275544 530550 275596
rect 530762 275544 530768 275596
rect 530820 275584 530826 275596
rect 534902 275584 534908 275596
rect 530820 275556 534908 275584
rect 530820 275544 530826 275556
rect 534902 275544 534908 275556
rect 534960 275544 534966 275596
rect 538030 275544 538036 275596
rect 538088 275584 538094 275596
rect 626166 275584 626172 275596
rect 538088 275556 626172 275584
rect 538088 275544 538094 275556
rect 626166 275544 626172 275556
rect 626224 275544 626230 275596
rect 467708 275420 502012 275448
rect 467708 275408 467714 275420
rect 504358 275408 504364 275460
rect 504416 275448 504422 275460
rect 538214 275448 538220 275460
rect 504416 275420 538220 275448
rect 504416 275408 504422 275420
rect 538214 275408 538220 275420
rect 538272 275408 538278 275460
rect 540974 275448 540980 275460
rect 538416 275420 540980 275448
rect 353996 275284 354674 275312
rect 353996 275272 354002 275284
rect 356330 275272 356336 275324
rect 356388 275312 356394 275324
rect 368474 275312 368480 275324
rect 356388 275284 368480 275312
rect 356388 275272 356394 275284
rect 368474 275272 368480 275284
rect 368532 275272 368538 275324
rect 375098 275272 375104 275324
rect 375156 275312 375162 275324
rect 403986 275312 403992 275324
rect 375156 275284 403992 275312
rect 375156 275272 375162 275284
rect 403986 275272 403992 275284
rect 404044 275272 404050 275324
rect 411254 275272 411260 275324
rect 411312 275312 411318 275324
rect 455966 275312 455972 275324
rect 411312 275284 455972 275312
rect 411312 275272 411318 275284
rect 455966 275272 455972 275284
rect 456024 275272 456030 275324
rect 456150 275272 456156 275324
rect 456208 275312 456214 275324
rect 512178 275312 512184 275324
rect 456208 275284 512184 275312
rect 456208 275272 456214 275284
rect 512178 275272 512184 275284
rect 512236 275272 512242 275324
rect 519354 275312 519360 275324
rect 512380 275284 519360 275312
rect 339000 275148 345014 275176
rect 339000 275136 339006 275148
rect 420914 275136 420920 275188
rect 420972 275176 420978 275188
rect 434714 275176 434720 275188
rect 420972 275148 434720 275176
rect 420972 275136 420978 275148
rect 434714 275136 434720 275148
rect 434772 275136 434778 275188
rect 437474 275136 437480 275188
rect 437532 275176 437538 275188
rect 450078 275176 450084 275188
rect 437532 275148 450084 275176
rect 437532 275136 437538 275148
rect 450078 275136 450084 275148
rect 450136 275136 450142 275188
rect 456794 275136 456800 275188
rect 456852 275176 456858 275188
rect 467834 275176 467840 275188
rect 456852 275148 467840 275176
rect 456852 275136 456858 275148
rect 467834 275136 467840 275148
rect 467892 275136 467898 275188
rect 468202 275136 468208 275188
rect 468260 275176 468266 275188
rect 494514 275176 494520 275188
rect 468260 275148 494520 275176
rect 468260 275136 468266 275148
rect 494514 275136 494520 275148
rect 494572 275136 494578 275188
rect 494698 275136 494704 275188
rect 494756 275176 494762 275188
rect 512380 275176 512408 275284
rect 519354 275272 519360 275284
rect 519412 275272 519418 275324
rect 519538 275272 519544 275324
rect 519596 275312 519602 275324
rect 537570 275312 537576 275324
rect 519596 275284 537576 275312
rect 519596 275272 519602 275284
rect 537570 275272 537576 275284
rect 537628 275272 537634 275324
rect 537754 275272 537760 275324
rect 537812 275312 537818 275324
rect 538416 275312 538444 275420
rect 540974 275408 540980 275420
rect 541032 275408 541038 275460
rect 541158 275408 541164 275460
rect 541216 275448 541222 275460
rect 544286 275448 544292 275460
rect 541216 275420 544292 275448
rect 541216 275408 541222 275420
rect 544286 275408 544292 275420
rect 544344 275408 544350 275460
rect 544470 275408 544476 275460
rect 544528 275448 544534 275460
rect 546034 275448 546040 275460
rect 544528 275420 546040 275448
rect 544528 275408 544534 275420
rect 546034 275408 546040 275420
rect 546092 275408 546098 275460
rect 546218 275408 546224 275460
rect 546276 275448 546282 275460
rect 641622 275448 641628 275460
rect 546276 275420 641628 275448
rect 546276 275408 546282 275420
rect 641622 275408 641628 275420
rect 641680 275408 641686 275460
rect 537812 275284 538444 275312
rect 537812 275272 537818 275284
rect 538582 275272 538588 275324
rect 538640 275312 538646 275324
rect 633342 275312 633348 275324
rect 538640 275284 633348 275312
rect 538640 275272 538646 275284
rect 633342 275272 633348 275284
rect 633400 275272 633406 275324
rect 590746 275176 590752 275188
rect 494756 275148 512408 275176
rect 512472 275148 590752 275176
rect 494756 275136 494762 275148
rect 224218 275068 224224 275120
rect 224276 275108 224282 275120
rect 226150 275108 226156 275120
rect 224276 275080 226156 275108
rect 224276 275068 224282 275080
rect 226150 275068 226156 275080
rect 226208 275068 226214 275120
rect 294046 275068 294052 275120
rect 294104 275108 294110 275120
rect 295150 275108 295156 275120
rect 294104 275080 295156 275108
rect 294104 275068 294110 275080
rect 295150 275068 295156 275080
rect 295208 275068 295214 275120
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 182082 275040 182088 275052
rect 135680 275012 182088 275040
rect 135680 275000 135686 275012
rect 182082 275000 182088 275012
rect 182140 275000 182146 275052
rect 449894 275000 449900 275052
rect 449952 275040 449958 275052
rect 460658 275040 460664 275052
rect 449952 275012 460664 275040
rect 449952 275000 449958 275012
rect 460658 275000 460664 275012
rect 460716 275000 460722 275052
rect 488534 275000 488540 275052
rect 488592 275040 488598 275052
rect 492582 275040 492588 275052
rect 488592 275012 492588 275040
rect 488592 275000 488598 275012
rect 492582 275000 492588 275012
rect 492640 275000 492646 275052
rect 494698 275000 494704 275052
rect 494756 275040 494762 275052
rect 498562 275040 498568 275052
rect 494756 275012 498568 275040
rect 494756 275000 494762 275012
rect 498562 275000 498568 275012
rect 498620 275000 498626 275052
rect 505094 275000 505100 275052
rect 505152 275040 505158 275052
rect 506842 275040 506848 275052
rect 505152 275012 506848 275040
rect 505152 275000 505158 275012
rect 506842 275000 506848 275012
rect 506900 275000 506906 275052
rect 507026 275000 507032 275052
rect 507084 275040 507090 275052
rect 512472 275040 512500 275148
rect 590746 275136 590752 275148
rect 590804 275136 590810 275188
rect 611354 275136 611360 275188
rect 611412 275176 611418 275188
rect 616782 275176 616788 275188
rect 611412 275148 616788 275176
rect 611412 275136 611418 275148
rect 616782 275136 616788 275148
rect 616840 275136 616846 275188
rect 619174 275136 619180 275188
rect 619232 275176 619238 275188
rect 623866 275176 623872 275188
rect 619232 275148 623872 275176
rect 619232 275136 619238 275148
rect 623866 275136 623872 275148
rect 623924 275136 623930 275188
rect 507084 275012 512500 275040
rect 507084 275000 507090 275012
rect 514018 275000 514024 275052
rect 514076 275040 514082 275052
rect 583662 275040 583668 275052
rect 514076 275012 583668 275040
rect 514076 275000 514082 275012
rect 583662 275000 583668 275012
rect 583720 275000 583726 275052
rect 71774 274932 71780 274984
rect 71832 274972 71838 274984
rect 73798 274972 73804 274984
rect 71832 274944 73804 274972
rect 71832 274932 71838 274944
rect 73798 274932 73804 274944
rect 73856 274932 73862 274984
rect 277486 274932 277492 274984
rect 277544 274972 277550 274984
rect 284294 274972 284300 274984
rect 277544 274944 284300 274972
rect 277544 274932 277550 274944
rect 284294 274932 284300 274944
rect 284352 274932 284358 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136542 274904 136548 274916
rect 129700 274876 136548 274904
rect 129700 274864 129706 274876
rect 136542 274864 136548 274876
rect 136600 274864 136606 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 185578 274904 185584 274916
rect 149848 274876 185584 274904
rect 149848 274864 149854 274876
rect 185578 274864 185584 274876
rect 185636 274864 185642 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 293402 274904 293408 274916
rect 289320 274876 293408 274904
rect 289320 274864 289326 274876
rect 293402 274864 293408 274876
rect 293460 274864 293466 274916
rect 471790 274864 471796 274916
rect 471848 274904 471854 274916
rect 523126 274904 523132 274916
rect 471848 274876 523132 274904
rect 471848 274864 471854 274876
rect 523126 274864 523132 274876
rect 523184 274864 523190 274916
rect 523310 274864 523316 274916
rect 523368 274904 523374 274916
rect 597830 274904 597836 274916
rect 523368 274876 597836 274904
rect 523368 274864 523374 274876
rect 597830 274864 597836 274876
rect 597888 274864 597894 274916
rect 283374 274796 283380 274848
rect 283432 274836 283438 274848
rect 289078 274836 289084 274848
rect 283432 274808 289084 274836
rect 283432 274796 283438 274808
rect 289078 274796 289084 274808
rect 289136 274796 289142 274848
rect 404262 274796 404268 274848
rect 404320 274836 404326 274848
rect 407482 274836 407488 274848
rect 404320 274808 407488 274836
rect 404320 274796 404326 274808
rect 407482 274796 407488 274808
rect 407540 274796 407546 274848
rect 426250 274796 426256 274848
rect 426308 274836 426314 274848
rect 432322 274836 432328 274848
rect 426308 274808 432328 274836
rect 426308 274796 426314 274808
rect 432322 274796 432328 274808
rect 432380 274796 432386 274848
rect 105998 274728 106004 274780
rect 106056 274768 106062 274780
rect 110414 274768 110420 274780
rect 106056 274740 110420 274768
rect 106056 274728 106062 274740
rect 110414 274728 110420 274740
rect 110472 274728 110478 274780
rect 140314 274728 140320 274780
rect 140372 274768 140378 274780
rect 144638 274768 144644 274780
rect 140372 274740 144644 274768
rect 140372 274728 140378 274740
rect 144638 274728 144644 274740
rect 144696 274728 144702 274780
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149882 274768 149888 274780
rect 146260 274740 149888 274768
rect 146260 274728 146266 274740
rect 149882 274728 149888 274740
rect 149940 274728 149946 274780
rect 435634 274728 435640 274780
rect 435692 274768 435698 274780
rect 439406 274768 439412 274780
rect 435692 274740 439412 274768
rect 435692 274728 435698 274740
rect 439406 274728 439412 274740
rect 439464 274728 439470 274780
rect 453942 274728 453948 274780
rect 454000 274768 454006 274780
rect 457162 274768 457168 274780
rect 454000 274740 457168 274768
rect 454000 274728 454006 274740
rect 457162 274728 457168 274740
rect 457220 274728 457226 274780
rect 464338 274728 464344 274780
rect 464396 274768 464402 274780
rect 471330 274768 471336 274780
rect 464396 274740 471336 274768
rect 464396 274728 464402 274740
rect 471330 274728 471336 274740
rect 471388 274728 471394 274780
rect 482922 274728 482928 274780
rect 482980 274768 482986 274780
rect 538674 274768 538680 274780
rect 482980 274740 538680 274768
rect 482980 274728 482986 274740
rect 538674 274728 538680 274740
rect 538732 274728 538738 274780
rect 539042 274728 539048 274780
rect 539100 274768 539106 274780
rect 545850 274768 545856 274780
rect 539100 274740 545856 274768
rect 539100 274728 539106 274740
rect 545850 274728 545856 274740
rect 545908 274728 545914 274780
rect 546034 274728 546040 274780
rect 546092 274768 546098 274780
rect 558822 274768 558828 274780
rect 546092 274740 558828 274768
rect 546092 274728 546098 274740
rect 558822 274728 558828 274740
rect 558880 274728 558886 274780
rect 570782 274728 570788 274780
rect 570840 274768 570846 274780
rect 570840 274740 571196 274768
rect 570840 274728 570846 274740
rect 66990 274660 66996 274712
rect 67048 274700 67054 274712
rect 71038 274700 71044 274712
rect 67048 274672 71044 274700
rect 67048 274660 67054 274672
rect 71038 274660 71044 274672
rect 71096 274660 71102 274712
rect 90634 274660 90640 274712
rect 90692 274700 90698 274712
rect 95878 274700 95884 274712
rect 90692 274672 95884 274700
rect 90692 274660 90698 274672
rect 95878 274660 95884 274672
rect 95936 274660 95942 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163130 274700 163136 274712
rect 161624 274672 163136 274700
rect 161624 274660 161630 274672
rect 163130 274660 163136 274672
rect 163188 274660 163194 274712
rect 170122 274660 170128 274712
rect 170180 274700 170186 274712
rect 173158 274700 173164 274712
rect 170180 274672 173164 274700
rect 170180 274660 170186 274672
rect 173158 274660 173164 274672
rect 173216 274660 173222 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 187142 274700 187148 274712
rect 185268 274672 187148 274700
rect 185268 274660 185274 274672
rect 187142 274660 187148 274672
rect 187200 274660 187206 274712
rect 238478 274660 238484 274712
rect 238536 274700 238542 274712
rect 239766 274700 239772 274712
rect 238536 274672 239772 274700
rect 238536 274660 238542 274672
rect 239766 274660 239772 274672
rect 239824 274660 239830 274712
rect 285766 274660 285772 274712
rect 285824 274700 285830 274712
rect 286962 274700 286968 274712
rect 285824 274672 286968 274700
rect 285824 274660 285830 274672
rect 286962 274660 286968 274672
rect 287020 274660 287026 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 360286 274660 360292 274712
rect 360344 274700 360350 274712
rect 363782 274700 363788 274712
rect 360344 274672 363788 274700
rect 360344 274660 360350 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 367094 274660 367100 274712
rect 367152 274700 367158 274712
rect 369670 274700 369676 274712
rect 367152 274672 369676 274700
rect 367152 274660 367158 274672
rect 369670 274660 369676 274672
rect 369728 274660 369734 274712
rect 386046 274660 386052 274712
rect 386104 274700 386110 274712
rect 389726 274700 389732 274712
rect 386104 274672 389732 274700
rect 386104 274660 386110 274672
rect 389726 274660 389732 274672
rect 389784 274660 389790 274712
rect 407114 274660 407120 274712
rect 407172 274700 407178 274712
rect 411070 274700 411076 274712
rect 407172 274672 411076 274700
rect 407172 274660 407178 274672
rect 411070 274660 411076 274672
rect 411128 274660 411134 274712
rect 104802 274592 104808 274644
rect 104860 274632 104866 274644
rect 157610 274632 157616 274644
rect 104860 274604 157616 274632
rect 104860 274592 104866 274604
rect 157610 274592 157616 274604
rect 157668 274592 157674 274644
rect 195882 274592 195888 274644
rect 195940 274632 195946 274644
rect 206278 274632 206284 274644
rect 195940 274604 206284 274632
rect 195940 274592 195946 274604
rect 206278 274592 206284 274604
rect 206336 274592 206342 274644
rect 424962 274592 424968 274644
rect 425020 274632 425026 274644
rect 474918 274632 474924 274644
rect 425020 274604 474924 274632
rect 425020 274592 425026 274604
rect 474918 274592 474924 274604
rect 474976 274592 474982 274644
rect 475378 274592 475384 274644
rect 475436 274632 475442 274644
rect 538122 274632 538128 274644
rect 475436 274604 538128 274632
rect 475436 274592 475442 274604
rect 538122 274592 538128 274604
rect 538180 274592 538186 274644
rect 539042 274592 539048 274644
rect 539100 274632 539106 274644
rect 570966 274632 570972 274644
rect 539100 274604 570972 274632
rect 539100 274592 539106 274604
rect 570966 274592 570972 274604
rect 571024 274592 571030 274644
rect 571168 274632 571196 274740
rect 571794 274632 571800 274644
rect 571168 274604 571800 274632
rect 571794 274592 571800 274604
rect 571852 274592 571858 274644
rect 577774 274632 577780 274644
rect 576826 274604 577780 274632
rect 121362 274456 121368 274508
rect 121420 274496 121426 274508
rect 176746 274496 176752 274508
rect 121420 274468 176752 274496
rect 121420 274456 121426 274468
rect 176746 274456 176752 274468
rect 176804 274456 176810 274508
rect 182910 274456 182916 274508
rect 182968 274496 182974 274508
rect 199654 274496 199660 274508
rect 182968 274468 199660 274496
rect 182968 274456 182974 274468
rect 199654 274456 199660 274468
rect 199712 274456 199718 274508
rect 210050 274456 210056 274508
rect 210108 274496 210114 274508
rect 237834 274496 237840 274508
rect 210108 274468 237840 274496
rect 210108 274456 210114 274468
rect 237834 274456 237840 274468
rect 237892 274456 237898 274508
rect 392578 274456 392584 274508
rect 392636 274496 392642 274508
rect 402790 274496 402796 274508
rect 392636 274468 402796 274496
rect 392636 274456 392642 274468
rect 402790 274456 402796 274468
rect 402848 274456 402854 274508
rect 406838 274456 406844 274508
rect 406896 274496 406902 274508
rect 437474 274496 437480 274508
rect 406896 274468 437480 274496
rect 406896 274456 406902 274468
rect 437474 274456 437480 274468
rect 437532 274456 437538 274508
rect 440878 274456 440884 274508
rect 440936 274496 440942 274508
rect 493778 274496 493784 274508
rect 440936 274468 493784 274496
rect 440936 274456 440942 274468
rect 493778 274456 493784 274468
rect 493836 274456 493842 274508
rect 496354 274456 496360 274508
rect 496412 274496 496418 274508
rect 576826 274496 576854 274604
rect 577774 274592 577780 274604
rect 577832 274592 577838 274644
rect 496412 274468 576854 274496
rect 496412 274456 496418 274468
rect 585778 274456 585784 274508
rect 585836 274496 585842 274508
rect 585836 274468 586514 274496
rect 585836 274456 585842 274468
rect 101306 274320 101312 274372
rect 101364 274360 101370 274372
rect 160922 274360 160928 274372
rect 101364 274332 160928 274360
rect 101364 274320 101370 274332
rect 160922 274320 160928 274332
rect 160980 274320 160986 274372
rect 187786 274320 187792 274372
rect 187844 274360 187850 274372
rect 220906 274360 220912 274372
rect 187844 274332 220912 274360
rect 187844 274320 187850 274332
rect 220906 274320 220912 274332
rect 220964 274320 220970 274372
rect 362862 274320 362868 274372
rect 362920 274360 362926 274372
rect 386230 274360 386236 274372
rect 362920 274332 386236 274360
rect 362920 274320 362926 274332
rect 386230 274320 386236 274332
rect 386288 274320 386294 274372
rect 395890 274320 395896 274372
rect 395948 274360 395954 274372
rect 420914 274360 420920 274372
rect 395948 274332 420920 274360
rect 395948 274320 395954 274332
rect 420914 274320 420920 274332
rect 420972 274320 420978 274372
rect 471238 274320 471244 274372
rect 471296 274360 471302 274372
rect 491478 274360 491484 274372
rect 471296 274332 491484 274360
rect 471296 274320 471302 274332
rect 491478 274320 491484 274332
rect 491536 274320 491542 274372
rect 492490 274320 492496 274372
rect 492548 274360 492554 274372
rect 570782 274360 570788 274372
rect 492548 274332 570788 274360
rect 492548 274320 492554 274332
rect 570782 274320 570788 274332
rect 570840 274320 570846 274372
rect 570966 274320 570972 274372
rect 571024 274360 571030 274372
rect 586054 274360 586060 274372
rect 571024 274332 586060 274360
rect 571024 274320 571030 274332
rect 586054 274320 586060 274332
rect 586112 274320 586118 274372
rect 586486 274360 586514 274468
rect 601418 274360 601424 274372
rect 586486 274332 601424 274360
rect 601418 274320 601424 274332
rect 601476 274320 601482 274372
rect 84746 274184 84752 274236
rect 84804 274224 84810 274236
rect 148318 274224 148324 274236
rect 84804 274196 148324 274224
rect 84804 274184 84810 274196
rect 148318 274184 148324 274196
rect 148376 274184 148382 274236
rect 160094 274184 160100 274236
rect 160152 274224 160158 274236
rect 164234 274224 164240 274236
rect 160152 274196 164240 274224
rect 160152 274184 160158 274196
rect 164234 274184 164240 274196
rect 164292 274184 164298 274236
rect 176930 274184 176936 274236
rect 176988 274224 176994 274236
rect 214650 274224 214656 274236
rect 176988 274196 214656 274224
rect 176988 274184 176994 274196
rect 214650 274184 214656 274196
rect 214708 274184 214714 274236
rect 220538 274184 220544 274236
rect 220596 274224 220602 274236
rect 240594 274224 240600 274236
rect 220596 274196 240600 274224
rect 220596 274184 220602 274196
rect 240594 274184 240600 274196
rect 240652 274184 240658 274236
rect 342898 274184 342904 274236
rect 342956 274224 342962 274236
rect 347222 274224 347228 274236
rect 342956 274196 347228 274224
rect 342956 274184 342962 274196
rect 347222 274184 347228 274196
rect 347280 274184 347286 274236
rect 366910 274184 366916 274236
rect 366968 274224 366974 274236
rect 389174 274224 389180 274236
rect 366968 274196 389180 274224
rect 366968 274184 366974 274196
rect 389174 274184 389180 274196
rect 389232 274184 389238 274236
rect 390278 274184 390284 274236
rect 390336 274224 390342 274236
rect 426434 274224 426440 274236
rect 390336 274196 426440 274224
rect 390336 274184 390342 274196
rect 426434 274184 426440 274196
rect 426492 274184 426498 274236
rect 438762 274184 438768 274236
rect 438820 274224 438826 274236
rect 496170 274224 496176 274236
rect 438820 274196 496176 274224
rect 438820 274184 438826 274196
rect 496170 274184 496176 274196
rect 496228 274184 496234 274236
rect 501966 274184 501972 274236
rect 502024 274224 502030 274236
rect 502024 274196 518296 274224
rect 502024 274184 502030 274196
rect 82354 274048 82360 274100
rect 82412 274088 82418 274100
rect 145558 274088 145564 274100
rect 82412 274060 145564 274088
rect 82412 274048 82418 274060
rect 145558 274048 145564 274060
rect 145616 274048 145622 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 200666 274088 200672 274100
rect 158128 274060 200672 274088
rect 158128 274048 158134 274060
rect 200666 274048 200672 274060
rect 200724 274048 200730 274100
rect 206554 274048 206560 274100
rect 206612 274088 206618 274100
rect 235442 274088 235448 274100
rect 206612 274060 235448 274088
rect 206612 274048 206618 274060
rect 235442 274048 235448 274060
rect 235500 274048 235506 274100
rect 239582 274048 239588 274100
rect 239640 274088 239646 274100
rect 258626 274088 258632 274100
rect 239640 274060 258632 274088
rect 239640 274048 239646 274060
rect 258626 274048 258632 274060
rect 258684 274048 258690 274100
rect 360102 274048 360108 274100
rect 360160 274088 360166 274100
rect 383838 274088 383844 274100
rect 360160 274060 383844 274088
rect 360160 274048 360166 274060
rect 383838 274048 383844 274060
rect 383896 274048 383902 274100
rect 384942 274048 384948 274100
rect 385000 274088 385006 274100
rect 419350 274088 419356 274100
rect 385000 274060 419356 274088
rect 385000 274048 385006 274060
rect 419350 274048 419356 274060
rect 419408 274048 419414 274100
rect 421558 274048 421564 274100
rect 421616 274088 421622 274100
rect 458358 274088 458364 274100
rect 421616 274060 458364 274088
rect 421616 274048 421622 274060
rect 458358 274048 458364 274060
rect 458416 274048 458422 274100
rect 459370 274048 459376 274100
rect 459428 274088 459434 274100
rect 516594 274088 516600 274100
rect 459428 274060 516600 274088
rect 459428 274048 459434 274060
rect 516594 274048 516600 274060
rect 516652 274048 516658 274100
rect 518268 274088 518296 274196
rect 518434 274184 518440 274236
rect 518492 274224 518498 274236
rect 602522 274224 602528 274236
rect 518492 274196 602528 274224
rect 518492 274184 518498 274196
rect 602522 274184 602528 274196
rect 602580 274184 602586 274236
rect 613378 274184 613384 274236
rect 613436 274224 613442 274236
rect 615586 274224 615592 274236
rect 613436 274196 615592 274224
rect 613436 274184 613442 274196
rect 615586 274184 615592 274196
rect 615644 274184 615650 274236
rect 533890 274088 533896 274100
rect 518268 274060 533896 274088
rect 533890 274048 533896 274060
rect 533948 274048 533954 274100
rect 534028 274048 534034 274100
rect 534086 274088 534092 274100
rect 619174 274088 619180 274100
rect 534086 274060 619180 274088
rect 534086 274048 534092 274060
rect 619174 274048 619180 274060
rect 619232 274048 619238 274100
rect 77202 273912 77208 273964
rect 77260 273952 77266 273964
rect 143534 273952 143540 273964
rect 77260 273924 143540 273952
rect 77260 273912 77266 273924
rect 143534 273912 143540 273924
rect 143592 273912 143598 273964
rect 145006 273912 145012 273964
rect 145064 273952 145070 273964
rect 192478 273952 192484 273964
rect 145064 273924 192484 273952
rect 145064 273912 145070 273924
rect 192478 273912 192484 273924
rect 192536 273912 192542 273964
rect 193490 273912 193496 273964
rect 193548 273952 193554 273964
rect 226334 273952 226340 273964
rect 193548 273924 226340 273952
rect 193548 273912 193554 273924
rect 226334 273912 226340 273924
rect 226392 273912 226398 273964
rect 234890 273912 234896 273964
rect 234948 273952 234954 273964
rect 255498 273952 255504 273964
rect 234948 273924 255504 273952
rect 234948 273912 234954 273924
rect 255498 273912 255504 273924
rect 255556 273912 255562 273964
rect 256142 273912 256148 273964
rect 256200 273952 256206 273964
rect 270586 273952 270592 273964
rect 256200 273924 270592 273952
rect 256200 273912 256206 273924
rect 270586 273912 270592 273924
rect 270644 273912 270650 273964
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280798 273952 280804 273964
rect 271564 273924 280804 273952
rect 271564 273912 271570 273924
rect 280798 273912 280804 273924
rect 280856 273912 280862 273964
rect 346302 273912 346308 273964
rect 346360 273952 346366 273964
rect 362586 273952 362592 273964
rect 346360 273924 362592 273952
rect 346360 273912 346366 273924
rect 362586 273912 362592 273924
rect 362644 273912 362650 273964
rect 377766 273912 377772 273964
rect 377824 273952 377830 273964
rect 408678 273952 408684 273964
rect 377824 273924 408684 273952
rect 377824 273912 377830 273924
rect 408678 273912 408684 273924
rect 408736 273912 408742 273964
rect 413922 273912 413928 273964
rect 413980 273952 413986 273964
rect 449894 273952 449900 273964
rect 413980 273924 449900 273952
rect 413980 273912 413986 273924
rect 449894 273912 449900 273924
rect 449952 273912 449958 273964
rect 451090 273912 451096 273964
rect 451148 273952 451154 273964
rect 513834 273952 513840 273964
rect 451148 273924 513840 273952
rect 451148 273912 451154 273924
rect 513834 273912 513840 273924
rect 513892 273912 513898 273964
rect 517054 273912 517060 273964
rect 517112 273952 517118 273964
rect 524230 273952 524236 273964
rect 517112 273924 524236 273952
rect 517112 273912 517118 273924
rect 524230 273912 524236 273924
rect 524288 273912 524294 273964
rect 524414 273912 524420 273964
rect 524472 273952 524478 273964
rect 613194 273952 613200 273964
rect 524472 273924 613200 273952
rect 524472 273912 524478 273924
rect 613194 273912 613200 273924
rect 613252 273912 613258 273964
rect 123754 273776 123760 273828
rect 123812 273816 123818 273828
rect 177482 273816 177488 273828
rect 123812 273788 177488 273816
rect 123812 273776 123818 273788
rect 177482 273776 177488 273788
rect 177540 273776 177546 273828
rect 426894 273776 426900 273828
rect 426952 273816 426958 273828
rect 477218 273816 477224 273828
rect 426952 273788 477224 273816
rect 426952 273776 426958 273788
rect 477218 273776 477224 273788
rect 477276 273776 477282 273828
rect 491202 273776 491208 273828
rect 491260 273816 491266 273828
rect 570598 273816 570604 273828
rect 491260 273788 570604 273816
rect 491260 273776 491266 273788
rect 570598 273776 570604 273788
rect 570656 273776 570662 273828
rect 587158 273816 587164 273828
rect 576826 273788 587164 273816
rect 280982 273708 280988 273760
rect 281040 273748 281046 273760
rect 287514 273748 287520 273760
rect 281040 273720 287520 273748
rect 281040 273708 281046 273720
rect 287514 273708 287520 273720
rect 287572 273708 287578 273760
rect 134426 273640 134432 273692
rect 134484 273680 134490 273692
rect 185026 273680 185032 273692
rect 134484 273652 185032 273680
rect 134484 273640 134490 273652
rect 185026 273640 185032 273652
rect 185084 273640 185090 273692
rect 460014 273640 460020 273692
rect 460072 273680 460078 273692
rect 484302 273680 484308 273692
rect 460072 273652 484308 273680
rect 460072 273640 460078 273652
rect 484302 273640 484308 273652
rect 484360 273640 484366 273692
rect 487982 273640 487988 273692
rect 488040 273680 488046 273692
rect 565906 273680 565912 273692
rect 488040 273652 565912 273680
rect 488040 273640 488046 273652
rect 565906 273640 565912 273652
rect 565964 273640 565970 273692
rect 570598 273640 570604 273692
rect 570656 273680 570662 273692
rect 576826 273680 576854 273788
rect 587158 273776 587164 273788
rect 587216 273776 587222 273828
rect 570656 273652 576854 273680
rect 570656 273640 570662 273652
rect 144638 273504 144644 273556
rect 144696 273544 144702 273556
rect 187786 273544 187792 273556
rect 144696 273516 187792 273544
rect 144696 273504 144702 273516
rect 187786 273504 187792 273516
rect 187844 273504 187850 273556
rect 429010 273504 429016 273556
rect 429068 273544 429074 273556
rect 482002 273544 482008 273556
rect 429068 273516 482008 273544
rect 429068 273504 429074 273516
rect 482002 273504 482008 273516
rect 482060 273504 482066 273556
rect 487062 273504 487068 273556
rect 487120 273544 487126 273556
rect 563514 273544 563520 273556
rect 487120 273516 563520 273544
rect 487120 273504 487126 273516
rect 563514 273504 563520 273516
rect 563572 273504 563578 273556
rect 481358 273368 481364 273420
rect 481416 273408 481422 273420
rect 556430 273408 556436 273420
rect 481416 273380 556436 273408
rect 481416 273368 481422 273380
rect 556430 273368 556436 273380
rect 556488 273368 556494 273420
rect 347038 273232 347044 273284
rect 347096 273272 347102 273284
rect 349614 273272 349620 273284
rect 347096 273244 349620 273272
rect 347096 273232 347102 273244
rect 349614 273232 349620 273244
rect 349672 273232 349678 273284
rect 350258 273232 350264 273284
rect 350316 273272 350322 273284
rect 356330 273272 356336 273284
rect 350316 273244 356336 273272
rect 350316 273232 350322 273244
rect 356330 273232 356336 273244
rect 356388 273232 356394 273284
rect 409138 273232 409144 273284
rect 409196 273272 409202 273284
rect 409874 273272 409880 273284
rect 409196 273244 409880 273272
rect 409196 273232 409202 273244
rect 409874 273232 409880 273244
rect 409932 273232 409938 273284
rect 114278 273164 114284 273216
rect 114336 273204 114342 273216
rect 169018 273204 169024 273216
rect 114336 273176 169024 273204
rect 114336 273164 114342 273176
rect 169018 273164 169024 273176
rect 169076 273164 169082 273216
rect 211982 273204 211988 273216
rect 200086 273176 211988 273204
rect 104986 273028 104992 273080
rect 105044 273068 105050 273080
rect 163314 273068 163320 273080
rect 105044 273040 163320 273068
rect 105044 273028 105050 273040
rect 163314 273028 163320 273040
rect 163372 273028 163378 273080
rect 167546 273028 167552 273080
rect 167604 273068 167610 273080
rect 184198 273068 184204 273080
rect 167604 273040 184204 273068
rect 167604 273028 167610 273040
rect 184198 273028 184204 273040
rect 184256 273028 184262 273080
rect 187602 273028 187608 273080
rect 187660 273068 187666 273080
rect 200086 273068 200114 273176
rect 211982 273164 211988 273176
rect 212040 273164 212046 273216
rect 419166 273164 419172 273216
rect 419224 273204 419230 273216
rect 456794 273204 456800 273216
rect 419224 273176 456800 273204
rect 419224 273164 419230 273176
rect 456794 273164 456800 273176
rect 456852 273164 456858 273216
rect 463510 273164 463516 273216
rect 463568 273204 463574 273216
rect 486878 273204 486884 273216
rect 463568 273176 486884 273204
rect 463568 273164 463574 273176
rect 486878 273164 486884 273176
rect 486936 273164 486942 273216
rect 493318 273164 493324 273216
rect 493376 273204 493382 273216
rect 574186 273204 574192 273216
rect 493376 273176 574192 273204
rect 493376 273164 493382 273176
rect 574186 273164 574192 273176
rect 574244 273164 574250 273216
rect 578878 273164 578884 273216
rect 578936 273204 578942 273216
rect 594334 273204 594340 273216
rect 578936 273176 594340 273204
rect 578936 273164 578942 273176
rect 594334 273164 594340 273176
rect 594392 273164 594398 273216
rect 187660 273040 200114 273068
rect 187660 273028 187666 273040
rect 211246 273028 211252 273080
rect 211304 273068 211310 273080
rect 220078 273068 220084 273080
rect 211304 273040 220084 273068
rect 211304 273028 211310 273040
rect 220078 273028 220084 273040
rect 220136 273028 220142 273080
rect 382918 273028 382924 273080
rect 382976 273068 382982 273080
rect 392118 273068 392124 273080
rect 382976 273040 392124 273068
rect 382976 273028 382982 273040
rect 392118 273028 392124 273040
rect 392176 273028 392182 273080
rect 403986 273028 403992 273080
rect 404044 273068 404050 273080
rect 429194 273068 429200 273080
rect 404044 273040 429200 273068
rect 404044 273028 404050 273040
rect 429194 273028 429200 273040
rect 429252 273028 429258 273080
rect 434622 273028 434628 273080
rect 434680 273068 434686 273080
rect 488718 273068 488724 273080
rect 434680 273040 488724 273068
rect 434680 273028 434686 273040
rect 488718 273028 488724 273040
rect 488776 273028 488782 273080
rect 496630 273028 496636 273080
rect 496688 273068 496694 273080
rect 578510 273068 578516 273080
rect 496688 273040 578516 273068
rect 496688 273028 496694 273040
rect 578510 273028 578516 273040
rect 578568 273028 578574 273080
rect 580258 273028 580264 273080
rect 580316 273068 580322 273080
rect 640426 273068 640432 273080
rect 580316 273040 640432 273068
rect 580316 273028 580322 273040
rect 640426 273028 640432 273040
rect 640484 273028 640490 273080
rect 78858 272892 78864 272944
rect 78916 272932 78922 272944
rect 138658 272932 138664 272944
rect 78916 272904 138664 272932
rect 78916 272892 78922 272904
rect 138658 272892 138664 272904
rect 138716 272892 138722 272944
rect 141786 272892 141792 272944
rect 141844 272932 141850 272944
rect 189810 272932 189816 272944
rect 141844 272904 189816 272932
rect 141844 272892 141850 272904
rect 189810 272892 189816 272904
rect 189868 272892 189874 272944
rect 191190 272892 191196 272944
rect 191248 272932 191254 272944
rect 224862 272932 224868 272944
rect 191248 272904 224868 272932
rect 191248 272892 191254 272904
rect 224862 272892 224868 272904
rect 224920 272892 224926 272944
rect 288066 272892 288072 272944
rect 288124 272932 288130 272944
rect 290458 272932 290464 272944
rect 288124 272904 290464 272932
rect 288124 272892 288130 272904
rect 290458 272892 290464 272904
rect 290516 272892 290522 272944
rect 373166 272892 373172 272944
rect 373224 272932 373230 272944
rect 382642 272932 382648 272944
rect 373224 272904 382648 272932
rect 373224 272892 373230 272904
rect 382642 272892 382648 272904
rect 382700 272892 382706 272944
rect 388622 272932 388628 272944
rect 383626 272904 388628 272932
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 156046 272796 156052 272808
rect 94280 272768 156052 272796
rect 94280 272756 94286 272768
rect 156046 272756 156052 272768
rect 156104 272756 156110 272808
rect 180518 272756 180524 272808
rect 180576 272796 180582 272808
rect 217226 272796 217232 272808
rect 180576 272768 217232 272796
rect 180576 272756 180582 272768
rect 217226 272756 217232 272768
rect 217284 272756 217290 272808
rect 228818 272756 228824 272808
rect 228876 272796 228882 272808
rect 249058 272796 249064 272808
rect 228876 272768 249064 272796
rect 228876 272756 228882 272768
rect 249058 272756 249064 272768
rect 249116 272756 249122 272808
rect 352926 272756 352932 272808
rect 352984 272796 352990 272808
rect 372982 272796 372988 272808
rect 352984 272768 372988 272796
rect 352984 272756 352990 272768
rect 372982 272756 372988 272768
rect 373040 272756 373046 272808
rect 380526 272756 380532 272808
rect 380584 272796 380590 272808
rect 383626 272796 383654 272904
rect 388622 272892 388628 272904
rect 388680 272892 388686 272944
rect 391842 272892 391848 272944
rect 391900 272932 391906 272944
rect 410058 272932 410064 272944
rect 391900 272904 410064 272932
rect 391900 272892 391906 272904
rect 410058 272892 410064 272904
rect 410116 272892 410122 272944
rect 412450 272892 412456 272944
rect 412508 272932 412514 272944
rect 453942 272932 453948 272944
rect 412508 272904 453948 272932
rect 412508 272892 412514 272904
rect 453942 272892 453948 272904
rect 454000 272892 454006 272944
rect 458082 272892 458088 272944
rect 458140 272932 458146 272944
rect 521838 272932 521844 272944
rect 458140 272904 521844 272932
rect 458140 272892 458146 272904
rect 521838 272892 521844 272904
rect 521896 272892 521902 272944
rect 524368 272932 524374 272944
rect 523604 272904 524374 272932
rect 394510 272796 394516 272808
rect 380584 272768 383654 272796
rect 388456 272768 394516 272796
rect 380584 272756 380590 272768
rect 87138 272620 87144 272672
rect 87196 272660 87202 272672
rect 151998 272660 152004 272672
rect 87196 272632 152004 272660
rect 87196 272620 87202 272632
rect 151998 272620 152004 272632
rect 152056 272620 152062 272672
rect 168650 272620 168656 272672
rect 168708 272660 168714 272672
rect 208486 272660 208492 272672
rect 168708 272632 208492 272660
rect 168708 272620 168714 272632
rect 208486 272620 208492 272632
rect 208544 272620 208550 272672
rect 217410 272620 217416 272672
rect 217468 272660 217474 272672
rect 242158 272660 242164 272672
rect 217468 272632 242164 272660
rect 217468 272620 217474 272632
rect 242158 272620 242164 272632
rect 242216 272620 242222 272672
rect 242342 272620 242348 272672
rect 242400 272660 242406 272672
rect 259546 272660 259552 272672
rect 242400 272632 259552 272660
rect 242400 272620 242406 272632
rect 259546 272620 259552 272632
rect 259604 272620 259610 272672
rect 331030 272620 331036 272672
rect 331088 272660 331094 272672
rect 342438 272660 342444 272672
rect 331088 272632 342444 272660
rect 331088 272620 331094 272632
rect 342438 272620 342444 272632
rect 342496 272620 342502 272672
rect 368382 272620 368388 272672
rect 368440 272660 368446 272672
rect 388456 272660 388484 272768
rect 394510 272756 394516 272768
rect 394568 272756 394574 272808
rect 397270 272756 397276 272808
rect 397328 272796 397334 272808
rect 418338 272796 418344 272808
rect 397328 272768 418344 272796
rect 397328 272756 397334 272768
rect 418338 272756 418344 272768
rect 418396 272756 418402 272808
rect 426066 272756 426072 272808
rect 426124 272796 426130 272808
rect 478414 272796 478420 272808
rect 426124 272768 478420 272796
rect 426124 272756 426130 272768
rect 478414 272756 478420 272768
rect 478472 272756 478478 272808
rect 482554 272756 482560 272808
rect 482612 272796 482618 272808
rect 523604 272796 523632 272904
rect 524368 272892 524374 272904
rect 524426 272892 524432 272944
rect 524506 272892 524512 272944
rect 524564 272932 524570 272944
rect 611354 272932 611360 272944
rect 524564 272904 611360 272932
rect 524564 272892 524570 272904
rect 611354 272892 611360 272904
rect 611412 272892 611418 272944
rect 606110 272796 606116 272808
rect 482612 272768 523632 272796
rect 523696 272768 606116 272796
rect 482612 272756 482618 272768
rect 368440 272632 388484 272660
rect 368440 272620 368446 272632
rect 388622 272620 388628 272672
rect 388680 272660 388686 272672
rect 393590 272660 393596 272672
rect 388680 272632 393596 272660
rect 388680 272620 388686 272632
rect 393590 272620 393596 272632
rect 393648 272620 393654 272672
rect 393958 272620 393964 272672
rect 394016 272660 394022 272672
rect 406286 272660 406292 272672
rect 394016 272632 406292 272660
rect 394016 272620 394022 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 408402 272620 408408 272672
rect 408460 272660 408466 272672
rect 452470 272660 452476 272672
rect 408460 272632 452476 272660
rect 408460 272620 408466 272632
rect 452470 272620 452476 272632
rect 452528 272620 452534 272672
rect 453850 272620 453856 272672
rect 453908 272660 453914 272672
rect 516410 272660 516416 272672
rect 453908 272632 516416 272660
rect 453908 272620 453914 272632
rect 516410 272620 516416 272632
rect 516468 272620 516474 272672
rect 516594 272620 516600 272672
rect 516652 272660 516658 272672
rect 523696 272660 523724 272768
rect 606110 272756 606116 272768
rect 606168 272756 606174 272808
rect 516652 272632 523724 272660
rect 516652 272620 516658 272632
rect 524322 272620 524328 272672
rect 524380 272660 524386 272672
rect 524506 272660 524512 272672
rect 524380 272632 524512 272660
rect 524380 272620 524386 272632
rect 524506 272620 524512 272632
rect 524564 272620 524570 272672
rect 524874 272620 524880 272672
rect 524932 272660 524938 272672
rect 614390 272660 614396 272672
rect 524932 272632 614396 272660
rect 524932 272620 524938 272632
rect 614390 272620 614396 272632
rect 614448 272620 614454 272672
rect 77662 272484 77668 272536
rect 77720 272524 77726 272536
rect 145098 272524 145104 272536
rect 77720 272496 145104 272524
rect 77720 272484 77726 272496
rect 145098 272484 145104 272496
rect 145156 272484 145162 272536
rect 152182 272484 152188 272536
rect 152240 272524 152246 272536
rect 197538 272524 197544 272536
rect 152240 272496 197544 272524
rect 152240 272484 152246 272496
rect 197538 272484 197544 272496
rect 197596 272484 197602 272536
rect 199470 272484 199476 272536
rect 199528 272524 199534 272536
rect 230566 272524 230572 272536
rect 199528 272496 230572 272524
rect 199528 272484 199534 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 252738 272524 252744 272536
rect 231452 272496 252744 272524
rect 231452 272484 231458 272496
rect 252738 272484 252744 272496
rect 252796 272484 252802 272536
rect 252922 272484 252928 272536
rect 252980 272524 252986 272536
rect 267734 272524 267740 272536
rect 252980 272496 267740 272524
rect 252980 272484 252986 272496
rect 267734 272484 267740 272496
rect 267792 272484 267798 272536
rect 268010 272484 268016 272536
rect 268068 272524 268074 272536
rect 278774 272524 278780 272536
rect 268068 272496 278780 272524
rect 268068 272484 268074 272496
rect 278774 272484 278780 272496
rect 278832 272484 278838 272536
rect 279786 272484 279792 272536
rect 279844 272524 279850 272536
rect 287146 272524 287152 272536
rect 279844 272496 287152 272524
rect 279844 272484 279850 272496
rect 287146 272484 287152 272496
rect 287204 272484 287210 272536
rect 338022 272484 338028 272536
rect 338080 272524 338086 272536
rect 351914 272524 351920 272536
rect 338080 272496 351920 272524
rect 338080 272484 338086 272496
rect 351914 272484 351920 272496
rect 351972 272484 351978 272536
rect 358630 272484 358636 272536
rect 358688 272524 358694 272536
rect 380342 272524 380348 272536
rect 358688 272496 380348 272524
rect 358688 272484 358694 272496
rect 380342 272484 380348 272496
rect 380400 272484 380406 272536
rect 380710 272484 380716 272536
rect 380768 272524 380774 272536
rect 413370 272524 413376 272536
rect 380768 272496 413376 272524
rect 380768 272484 380774 272496
rect 413370 272484 413376 272496
rect 413428 272484 413434 272536
rect 415118 272484 415124 272536
rect 415176 272524 415182 272536
rect 461854 272524 461860 272536
rect 415176 272496 461860 272524
rect 415176 272484 415182 272496
rect 461854 272484 461860 272496
rect 461912 272484 461918 272536
rect 463326 272484 463332 272536
rect 463384 272524 463390 272536
rect 524506 272524 524512 272536
rect 463384 272496 524512 272524
rect 463384 272484 463390 272496
rect 524506 272484 524512 272496
rect 524564 272484 524570 272536
rect 524690 272484 524696 272536
rect 524748 272524 524754 272536
rect 533982 272524 533988 272536
rect 524748 272496 533988 272524
rect 524748 272484 524754 272496
rect 533982 272484 533988 272496
rect 534040 272484 534046 272536
rect 534166 272484 534172 272536
rect 534224 272524 534230 272536
rect 632146 272524 632152 272536
rect 534224 272496 632152 272524
rect 534224 272484 534230 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 127342 272348 127348 272400
rect 127400 272388 127406 272400
rect 179874 272388 179880 272400
rect 127400 272360 179880 272388
rect 127400 272348 127406 272360
rect 179874 272348 179880 272360
rect 179932 272348 179938 272400
rect 439314 272348 439320 272400
rect 439372 272388 439378 272400
rect 473722 272388 473728 272400
rect 439372 272360 473728 272388
rect 439372 272348 439378 272360
rect 473722 272348 473728 272360
rect 473780 272348 473786 272400
rect 474642 272348 474648 272400
rect 474700 272388 474706 272400
rect 495434 272388 495440 272400
rect 474700 272360 495440 272388
rect 474700 272348 474706 272360
rect 495434 272348 495440 272360
rect 495492 272348 495498 272400
rect 501598 272348 501604 272400
rect 501656 272388 501662 272400
rect 581270 272388 581276 272400
rect 501656 272360 581276 272388
rect 501656 272348 501662 272360
rect 581270 272348 581276 272360
rect 581328 272348 581334 272400
rect 139118 272212 139124 272264
rect 139176 272252 139182 272264
rect 141418 272252 141424 272264
rect 139176 272224 141424 272252
rect 139176 272212 139182 272224
rect 141418 272212 141424 272224
rect 141476 272212 141482 272264
rect 143902 272212 143908 272264
rect 143960 272252 143966 272264
rect 190730 272252 190736 272264
rect 143960 272224 190736 272252
rect 143960 272212 143966 272224
rect 190730 272212 190736 272224
rect 190788 272212 190794 272264
rect 451918 272212 451924 272264
rect 451976 272252 451982 272264
rect 480806 272252 480812 272264
rect 451976 272224 480812 272252
rect 451976 272212 451982 272224
rect 480806 272212 480812 272224
rect 480864 272212 480870 272264
rect 488350 272212 488356 272264
rect 488408 272252 488414 272264
rect 567102 272252 567108 272264
rect 488408 272224 567108 272252
rect 488408 272212 488414 272224
rect 567102 272212 567108 272224
rect 567160 272212 567166 272264
rect 153286 272076 153292 272128
rect 153344 272116 153350 272128
rect 171778 272116 171784 272128
rect 153344 272088 171784 272116
rect 153344 272076 153350 272088
rect 171778 272076 171784 272088
rect 171836 272076 171842 272128
rect 473078 272076 473084 272128
rect 473136 272116 473142 272128
rect 482922 272116 482928 272128
rect 473136 272088 482928 272116
rect 473136 272076 473142 272088
rect 482922 272076 482928 272088
rect 482980 272076 482986 272128
rect 483382 272076 483388 272128
rect 483440 272116 483446 272128
rect 560018 272116 560024 272128
rect 483440 272088 560024 272116
rect 483440 272076 483446 272088
rect 560018 272076 560024 272088
rect 560076 272076 560082 272128
rect 478414 271940 478420 271992
rect 478472 271980 478478 271992
rect 552474 271980 552480 271992
rect 478472 271952 552480 271980
rect 478472 271940 478478 271952
rect 552474 271940 552480 271952
rect 552532 271940 552538 271992
rect 552842 271940 552848 271992
rect 552900 271980 552906 271992
rect 580074 271980 580080 271992
rect 552900 271952 580080 271980
rect 552900 271940 552906 271952
rect 580074 271940 580080 271952
rect 580132 271940 580138 271992
rect 110414 271804 110420 271856
rect 110472 271844 110478 271856
rect 164970 271844 164976 271856
rect 110472 271816 164976 271844
rect 110472 271804 110478 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 175826 271804 175832 271856
rect 175884 271844 175890 271856
rect 207658 271844 207664 271856
rect 175884 271816 207664 271844
rect 175884 271804 175890 271816
rect 207658 271804 207664 271816
rect 207716 271804 207722 271856
rect 214834 271804 214840 271856
rect 214892 271844 214898 271856
rect 221458 271844 221464 271856
rect 214892 271816 221464 271844
rect 214892 271804 214898 271816
rect 221458 271804 221464 271816
rect 221516 271804 221522 271856
rect 222102 271804 222108 271856
rect 222160 271844 222166 271856
rect 232130 271844 232136 271856
rect 222160 271816 232136 271844
rect 222160 271804 222166 271816
rect 232130 271804 232136 271816
rect 232188 271804 232194 271856
rect 356514 271804 356520 271856
rect 356572 271844 356578 271856
rect 358998 271844 359004 271856
rect 356572 271816 359004 271844
rect 356572 271804 356578 271816
rect 358998 271804 359004 271816
rect 359056 271804 359062 271856
rect 394326 271804 394332 271856
rect 394384 271844 394390 271856
rect 426250 271844 426256 271856
rect 394384 271816 426256 271844
rect 394384 271804 394390 271816
rect 426250 271804 426256 271816
rect 426308 271804 426314 271856
rect 427078 271804 427084 271856
rect 427136 271844 427142 271856
rect 433518 271844 433524 271856
rect 427136 271816 433524 271844
rect 427136 271804 427142 271816
rect 433518 271804 433524 271816
rect 433576 271804 433582 271856
rect 447778 271804 447784 271856
rect 447836 271844 447842 271856
rect 504542 271844 504548 271856
rect 447836 271816 504548 271844
rect 447836 271804 447842 271816
rect 504542 271804 504548 271816
rect 504600 271804 504606 271856
rect 504726 271804 504732 271856
rect 504784 271844 504790 271856
rect 589550 271844 589556 271856
rect 504784 271816 589556 271844
rect 504784 271804 504790 271816
rect 589550 271804 589556 271816
rect 589608 271804 589614 271856
rect 596634 271844 596640 271856
rect 591316 271816 596640 271844
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 93026 271668 93032 271720
rect 93084 271708 93090 271720
rect 120718 271708 120724 271720
rect 93084 271680 120724 271708
rect 93084 271668 93090 271680
rect 120718 271668 120724 271680
rect 120776 271668 120782 271720
rect 120902 271668 120908 271720
rect 120960 271708 120966 271720
rect 175274 271708 175280 271720
rect 120960 271680 175280 271708
rect 120960 271668 120966 271680
rect 175274 271668 175280 271680
rect 175332 271668 175338 271720
rect 192294 271668 192300 271720
rect 192352 271708 192358 271720
rect 225506 271708 225512 271720
rect 192352 271680 225512 271708
rect 192352 271668 192358 271680
rect 225506 271668 225512 271680
rect 225564 271668 225570 271720
rect 237466 271668 237472 271720
rect 237524 271708 237530 271720
rect 243722 271708 243728 271720
rect 237524 271680 243728 271708
rect 237524 271668 237530 271680
rect 243722 271668 243728 271680
rect 243780 271668 243786 271720
rect 355318 271668 355324 271720
rect 355376 271708 355382 271720
rect 374362 271708 374368 271720
rect 355376 271680 374368 271708
rect 355376 271668 355382 271680
rect 374362 271668 374368 271680
rect 374420 271668 374426 271720
rect 387702 271668 387708 271720
rect 387760 271708 387766 271720
rect 421374 271708 421380 271720
rect 387760 271680 421380 271708
rect 387760 271668 387766 271680
rect 421374 271668 421380 271680
rect 421432 271668 421438 271720
rect 421742 271668 421748 271720
rect 421800 271708 421806 271720
rect 438210 271708 438216 271720
rect 421800 271680 438216 271708
rect 421800 271668 421806 271680
rect 438210 271668 438216 271680
rect 438268 271668 438274 271720
rect 442902 271668 442908 271720
rect 442960 271708 442966 271720
rect 500494 271708 500500 271720
rect 442960 271680 500500 271708
rect 442960 271668 442966 271680
rect 500494 271668 500500 271680
rect 500552 271668 500558 271720
rect 500862 271668 500868 271720
rect 500920 271708 500926 271720
rect 508038 271708 508044 271720
rect 500920 271680 508044 271708
rect 500920 271668 500926 271680
rect 508038 271668 508044 271680
rect 508096 271668 508102 271720
rect 508958 271668 508964 271720
rect 509016 271708 509022 271720
rect 591316 271708 591344 271816
rect 596634 271804 596640 271816
rect 596692 271804 596698 271856
rect 509016 271680 591344 271708
rect 509016 271668 509022 271680
rect 591482 271668 591488 271720
rect 591540 271708 591546 271720
rect 603718 271708 603724 271720
rect 591540 271680 603724 271708
rect 591540 271668 591546 271680
rect 603718 271668 603724 271680
rect 603776 271668 603782 271720
rect 111978 271532 111984 271584
rect 112036 271572 112042 271584
rect 168374 271572 168380 271584
rect 112036 271544 168380 271572
rect 112036 271532 112042 271544
rect 168374 271532 168380 271544
rect 168432 271532 168438 271584
rect 173434 271532 173440 271584
rect 173492 271572 173498 271584
rect 212626 271572 212632 271584
rect 173492 271544 212632 271572
rect 173492 271532 173498 271544
rect 212626 271532 212632 271544
rect 212684 271532 212690 271584
rect 226150 271532 226156 271584
rect 226208 271572 226214 271584
rect 247218 271572 247224 271584
rect 226208 271544 247224 271572
rect 226208 271532 226214 271544
rect 247218 271532 247224 271544
rect 247276 271532 247282 271584
rect 259730 271532 259736 271584
rect 259788 271572 259794 271584
rect 272610 271572 272616 271584
rect 259788 271544 272616 271572
rect 259788 271532 259794 271544
rect 272610 271532 272616 271544
rect 272668 271532 272674 271584
rect 372522 271532 372528 271584
rect 372580 271572 372586 271584
rect 400398 271572 400404 271584
rect 372580 271544 400404 271572
rect 372580 271532 372586 271544
rect 400398 271532 400404 271544
rect 400456 271532 400462 271584
rect 409782 271532 409788 271584
rect 409840 271572 409846 271584
rect 443730 271572 443736 271584
rect 409840 271544 443736 271572
rect 409840 271532 409846 271544
rect 443730 271532 443736 271544
rect 443788 271532 443794 271584
rect 453298 271532 453304 271584
rect 453356 271572 453362 271584
rect 511534 271572 511540 271584
rect 453356 271544 511540 271572
rect 453356 271532 453362 271544
rect 511534 271532 511540 271544
rect 511592 271532 511598 271584
rect 511902 271532 511908 271584
rect 511960 271572 511966 271584
rect 600222 271572 600228 271584
rect 511960 271544 600228 271572
rect 511960 271532 511966 271544
rect 600222 271532 600228 271544
rect 600280 271532 600286 271584
rect 607858 271532 607864 271584
rect 607916 271572 607922 271584
rect 643922 271572 643928 271584
rect 607916 271544 643928 271572
rect 607916 271532 607922 271544
rect 643922 271532 643928 271544
rect 643980 271532 643986 271584
rect 89714 271396 89720 271448
rect 89772 271436 89778 271448
rect 152642 271436 152648 271448
rect 89772 271408 152648 271436
rect 89772 271396 89778 271408
rect 152642 271396 152648 271408
rect 152700 271396 152706 271448
rect 165154 271396 165160 271448
rect 165212 271436 165218 271448
rect 205726 271436 205732 271448
rect 165212 271408 205732 271436
rect 165212 271396 165218 271408
rect 205726 271396 205732 271408
rect 205784 271396 205790 271448
rect 223574 271396 223580 271448
rect 223632 271436 223638 271448
rect 247402 271436 247408 271448
rect 223632 271408 247408 271436
rect 223632 271396 223638 271408
rect 247402 271396 247408 271408
rect 247460 271396 247466 271448
rect 247862 271396 247868 271448
rect 247920 271436 247926 271448
rect 264330 271436 264336 271448
rect 247920 271408 264336 271436
rect 247920 271396 247926 271408
rect 264330 271396 264336 271408
rect 264388 271396 264394 271448
rect 334618 271396 334624 271448
rect 334676 271436 334682 271448
rect 341334 271436 341340 271448
rect 334676 271408 341340 271436
rect 334676 271396 334682 271408
rect 341334 271396 341340 271408
rect 341392 271396 341398 271448
rect 342162 271396 342168 271448
rect 342220 271436 342226 271448
rect 356698 271436 356704 271448
rect 342220 271408 356704 271436
rect 342220 271396 342226 271408
rect 356698 271396 356704 271408
rect 356756 271396 356762 271448
rect 360838 271396 360844 271448
rect 360896 271436 360902 271448
rect 381538 271436 381544 271448
rect 360896 271408 381544 271436
rect 360896 271396 360902 271408
rect 381538 271396 381544 271408
rect 381596 271396 381602 271448
rect 397914 271396 397920 271448
rect 397972 271436 397978 271448
rect 427078 271436 427084 271448
rect 397972 271408 427084 271436
rect 397972 271396 397978 271408
rect 427078 271396 427084 271408
rect 427136 271396 427142 271448
rect 427262 271396 427268 271448
rect 427320 271436 427326 271448
rect 427320 271408 436784 271436
rect 427320 271396 427326 271408
rect 72970 271260 72976 271312
rect 73028 271300 73034 271312
rect 142154 271300 142160 271312
rect 73028 271272 142160 271300
rect 73028 271260 73034 271272
rect 142154 271260 142160 271272
rect 142212 271260 142218 271312
rect 150986 271260 150992 271312
rect 151044 271300 151050 271312
rect 195974 271300 195980 271312
rect 151044 271272 195980 271300
rect 151044 271260 151050 271272
rect 195974 271260 195980 271272
rect 196032 271260 196038 271312
rect 215938 271260 215944 271312
rect 215996 271300 216002 271312
rect 242066 271300 242072 271312
rect 215996 271272 242072 271300
rect 215996 271260 216002 271272
rect 242066 271260 242072 271272
rect 242124 271260 242130 271312
rect 243170 271260 243176 271312
rect 243228 271300 243234 271312
rect 261018 271300 261024 271312
rect 243228 271272 261024 271300
rect 243228 271260 243234 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 275094 271260 275100 271312
rect 275152 271300 275158 271312
rect 283466 271300 283472 271312
rect 275152 271272 283472 271300
rect 275152 271260 275158 271272
rect 283466 271260 283472 271272
rect 283524 271260 283530 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 325510 271260 325516 271312
rect 325568 271300 325574 271312
rect 334158 271300 334164 271312
rect 325568 271272 334164 271300
rect 325568 271260 325574 271272
rect 334158 271260 334164 271272
rect 334216 271260 334222 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355502 271300 355508 271312
rect 340656 271272 355508 271300
rect 340656 271260 340662 271272
rect 355502 271260 355508 271272
rect 355560 271260 355566 271312
rect 364150 271260 364156 271312
rect 364208 271300 364214 271312
rect 386046 271300 386052 271312
rect 364208 271272 386052 271300
rect 364208 271260 364214 271272
rect 386046 271260 386052 271272
rect 386104 271260 386110 271312
rect 400122 271260 400128 271312
rect 400180 271300 400186 271312
rect 435634 271300 435640 271312
rect 400180 271272 435640 271300
rect 400180 271260 400186 271272
rect 435634 271260 435640 271272
rect 435692 271260 435698 271312
rect 436756 271300 436784 271408
rect 436922 271396 436928 271448
rect 436980 271436 436986 271448
rect 454770 271436 454776 271448
rect 436980 271408 454776 271436
rect 436980 271396 436986 271408
rect 454770 271396 454776 271408
rect 454828 271396 454834 271448
rect 457438 271396 457444 271448
rect 457496 271436 457502 271448
rect 511718 271436 511724 271448
rect 457496 271408 511724 271436
rect 457496 271396 457502 271408
rect 511718 271396 511724 271408
rect 511776 271396 511782 271448
rect 515122 271436 515128 271448
rect 512196 271408 515128 271436
rect 448882 271300 448888 271312
rect 436756 271272 448888 271300
rect 448882 271260 448888 271272
rect 448940 271260 448946 271312
rect 454678 271260 454684 271312
rect 454736 271300 454742 271312
rect 512196 271300 512224 271408
rect 515122 271396 515128 271408
rect 515180 271396 515186 271448
rect 515306 271396 515312 271448
rect 515364 271436 515370 271448
rect 518618 271436 518624 271448
rect 515364 271408 518624 271436
rect 515364 271396 515370 271408
rect 518618 271396 518624 271408
rect 518676 271396 518682 271448
rect 520090 271396 520096 271448
rect 520148 271436 520154 271448
rect 523954 271436 523960 271448
rect 520148 271408 523960 271436
rect 520148 271396 520154 271408
rect 523954 271396 523960 271408
rect 524012 271396 524018 271448
rect 524138 271396 524144 271448
rect 524196 271436 524202 271448
rect 524196 271408 529244 271436
rect 524196 271396 524202 271408
rect 454736 271272 512224 271300
rect 454736 271260 454742 271272
rect 514478 271260 514484 271312
rect 514536 271300 514542 271312
rect 529014 271300 529020 271312
rect 514536 271272 529020 271300
rect 514536 271260 514542 271272
rect 529014 271260 529020 271272
rect 529072 271260 529078 271312
rect 529216 271300 529244 271408
rect 529382 271396 529388 271448
rect 529440 271436 529446 271448
rect 610802 271436 610808 271448
rect 529440 271408 610808 271436
rect 529440 271396 529446 271408
rect 610802 271396 610808 271408
rect 610860 271396 610866 271448
rect 617978 271300 617984 271312
rect 529216 271272 617984 271300
rect 617978 271260 617984 271272
rect 618036 271260 618042 271312
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 208854 271124 208860 271176
rect 208912 271164 208918 271176
rect 237466 271164 237472 271176
rect 208912 271136 237472 271164
rect 208912 271124 208918 271136
rect 237466 271124 237472 271136
rect 237524 271124 237530 271176
rect 240778 271124 240784 271176
rect 240836 271164 240842 271176
rect 259822 271164 259828 271176
rect 240836 271136 259828 271164
rect 240836 271124 240842 271136
rect 259822 271124 259828 271136
rect 259880 271124 259886 271176
rect 262122 271124 262128 271176
rect 262180 271164 262186 271176
rect 274634 271164 274640 271176
rect 262180 271136 274640 271164
rect 262180 271124 262186 271136
rect 274634 271124 274640 271136
rect 274692 271124 274698 271176
rect 276290 271124 276296 271176
rect 276348 271164 276354 271176
rect 284478 271164 284484 271176
rect 276348 271136 284484 271164
rect 276348 271124 276354 271136
rect 284478 271124 284484 271136
rect 284536 271124 284542 271176
rect 333882 271124 333888 271176
rect 333940 271164 333946 271176
rect 344462 271164 344468 271176
rect 333940 271136 344468 271164
rect 333940 271124 333946 271136
rect 344462 271124 344468 271136
rect 344520 271124 344526 271176
rect 344646 271124 344652 271176
rect 344704 271164 344710 271176
rect 350718 271164 350724 271176
rect 344704 271136 350724 271164
rect 344704 271124 344710 271136
rect 350718 271124 350724 271136
rect 350776 271124 350782 271176
rect 351822 271124 351828 271176
rect 351880 271164 351886 271176
rect 372062 271164 372068 271176
rect 351880 271136 372068 271164
rect 351880 271124 351886 271136
rect 372062 271124 372068 271136
rect 372120 271124 372126 271176
rect 379422 271124 379428 271176
rect 379480 271164 379486 271176
rect 407114 271164 407120 271176
rect 379480 271136 407120 271164
rect 379480 271124 379486 271136
rect 407114 271124 407120 271136
rect 407172 271124 407178 271176
rect 416590 271124 416596 271176
rect 416648 271164 416654 271176
rect 463970 271164 463976 271176
rect 416648 271136 463976 271164
rect 416648 271124 416654 271136
rect 463970 271124 463976 271136
rect 464028 271124 464034 271176
rect 464522 271124 464528 271176
rect 464580 271164 464586 271176
rect 524506 271164 524512 271176
rect 464580 271136 524512 271164
rect 464580 271124 464586 271136
rect 524506 271124 524512 271136
rect 524564 271124 524570 271176
rect 524690 271124 524696 271176
rect 524748 271164 524754 271176
rect 529382 271164 529388 271176
rect 524748 271136 529388 271164
rect 524748 271124 524754 271136
rect 529382 271124 529388 271136
rect 529440 271124 529446 271176
rect 529566 271124 529572 271176
rect 529624 271164 529630 271176
rect 532786 271164 532792 271176
rect 529624 271136 532792 271164
rect 529624 271124 529630 271136
rect 532786 271124 532792 271136
rect 532844 271124 532850 271176
rect 533154 271124 533160 271176
rect 533212 271164 533218 271176
rect 621474 271164 621480 271176
rect 533212 271136 621480 271164
rect 533212 271124 533218 271136
rect 621474 271124 621480 271136
rect 621532 271124 621538 271176
rect 621658 271124 621664 271176
rect 621716 271164 621722 271176
rect 636838 271164 636844 271176
rect 621716 271136 636844 271164
rect 621716 271124 621722 271136
rect 636838 271124 636844 271136
rect 636896 271124 636902 271176
rect 128538 270988 128544 271040
rect 128596 271028 128602 271040
rect 181346 271028 181352 271040
rect 128596 271000 181352 271028
rect 128596 270988 128602 271000
rect 181346 270988 181352 271000
rect 181404 270988 181410 271040
rect 189994 270988 190000 271040
rect 190052 271028 190058 271040
rect 216122 271028 216128 271040
rect 190052 271000 216128 271028
rect 190052 270988 190058 271000
rect 216122 270988 216128 271000
rect 216180 270988 216186 271040
rect 381538 270988 381544 271040
rect 381596 271028 381602 271040
rect 399202 271028 399208 271040
rect 381596 271000 399208 271028
rect 381596 270988 381602 271000
rect 399202 270988 399208 271000
rect 399260 270988 399266 271040
rect 401318 270988 401324 271040
rect 401376 271028 401382 271040
rect 401376 271000 422294 271028
rect 401376 270988 401382 271000
rect 130838 270852 130844 270904
rect 130896 270892 130902 270904
rect 182450 270892 182456 270904
rect 130896 270864 182456 270892
rect 130896 270852 130902 270864
rect 182450 270852 182456 270864
rect 182508 270852 182514 270904
rect 200482 270852 200488 270904
rect 200540 270892 200546 270904
rect 224218 270892 224224 270904
rect 200540 270864 224224 270892
rect 200540 270852 200546 270864
rect 224218 270852 224224 270864
rect 224276 270852 224282 270904
rect 389082 270852 389088 270904
rect 389140 270892 389146 270904
rect 415302 270892 415308 270904
rect 389140 270864 415308 270892
rect 389140 270852 389146 270864
rect 415302 270852 415308 270864
rect 415360 270852 415366 270904
rect 422266 270892 422294 271000
rect 425698 270988 425704 271040
rect 425756 271028 425762 271040
rect 427262 271028 427268 271040
rect 425756 271000 427268 271028
rect 425756 270988 425762 271000
rect 427262 270988 427268 271000
rect 427320 270988 427326 271040
rect 431678 270988 431684 271040
rect 431736 271028 431742 271040
rect 485498 271028 485504 271040
rect 431736 271000 485504 271028
rect 431736 270988 431742 271000
rect 485498 270988 485504 271000
rect 485556 270988 485562 271040
rect 488718 270988 488724 271040
rect 488776 271028 488782 271040
rect 551738 271028 551744 271040
rect 488776 271000 551744 271028
rect 488776 270988 488782 271000
rect 551738 270988 551744 271000
rect 551796 270988 551802 271040
rect 552658 270988 552664 271040
rect 552716 271028 552722 271040
rect 591482 271028 591488 271040
rect 552716 271000 591488 271028
rect 552716 270988 552722 271000
rect 591482 270988 591488 271000
rect 591540 270988 591546 271040
rect 427814 270892 427820 270904
rect 422266 270864 427820 270892
rect 427814 270852 427820 270864
rect 427872 270852 427878 270904
rect 435358 270852 435364 270904
rect 435416 270892 435422 270904
rect 436922 270892 436928 270904
rect 435416 270864 436928 270892
rect 435416 270852 435422 270864
rect 436922 270852 436928 270864
rect 436980 270852 436986 270904
rect 445018 270852 445024 270904
rect 445076 270892 445082 270904
rect 497366 270892 497372 270904
rect 445076 270864 497372 270892
rect 445076 270852 445082 270864
rect 497366 270852 497372 270864
rect 497424 270852 497430 270904
rect 507670 270852 507676 270904
rect 507728 270892 507734 270904
rect 522022 270892 522028 270904
rect 507728 270864 522028 270892
rect 507728 270852 507734 270864
rect 522022 270852 522028 270864
rect 522080 270852 522086 270904
rect 524782 270852 524788 270904
rect 524840 270892 524846 270904
rect 593138 270892 593144 270904
rect 524840 270864 593144 270892
rect 524840 270852 524846 270864
rect 593138 270852 593144 270864
rect 593196 270852 593202 270904
rect 137922 270716 137928 270768
rect 137980 270756 137986 270768
rect 187878 270756 187884 270768
rect 137980 270728 187884 270756
rect 137980 270716 137986 270728
rect 187878 270716 187884 270728
rect 187936 270716 187942 270768
rect 433150 270716 433156 270768
rect 433208 270756 433214 270768
rect 456978 270756 456984 270768
rect 433208 270728 456984 270756
rect 433208 270716 433214 270728
rect 456978 270716 456984 270728
rect 457036 270716 457042 270768
rect 465718 270716 465724 270768
rect 465776 270756 465782 270768
rect 526254 270756 526260 270768
rect 465776 270728 526260 270756
rect 465776 270716 465782 270728
rect 526254 270716 526260 270728
rect 526312 270716 526318 270768
rect 526438 270716 526444 270768
rect 526496 270756 526502 270768
rect 528646 270756 528652 270768
rect 526496 270728 528652 270756
rect 526496 270716 526502 270728
rect 528646 270716 528652 270728
rect 528704 270716 528710 270768
rect 529014 270716 529020 270768
rect 529072 270756 529078 270768
rect 529072 270728 539088 270756
rect 529072 270716 529078 270728
rect 116670 270580 116676 270632
rect 116728 270620 116734 270632
rect 151078 270620 151084 270632
rect 116728 270592 151084 270620
rect 116728 270580 116734 270592
rect 151078 270580 151084 270592
rect 151136 270580 151142 270632
rect 237282 270580 237288 270632
rect 237340 270620 237346 270632
rect 237340 270592 237512 270620
rect 237340 270580 237346 270592
rect 115842 270444 115848 270496
rect 115900 270484 115906 270496
rect 171226 270484 171232 270496
rect 115900 270456 171232 270484
rect 115900 270444 115906 270456
rect 171226 270444 171232 270456
rect 171284 270444 171290 270496
rect 173158 270444 173164 270496
rect 173216 270484 173222 270496
rect 210142 270484 210148 270496
rect 173216 270456 210148 270484
rect 173216 270444 173222 270456
rect 210142 270444 210148 270456
rect 210200 270444 210206 270496
rect 210786 270444 210792 270496
rect 210844 270484 210850 270496
rect 211798 270484 211804 270496
rect 210844 270456 211804 270484
rect 210844 270444 210850 270456
rect 211798 270444 211804 270456
rect 211856 270444 211862 270496
rect 233142 270444 233148 270496
rect 233200 270484 233206 270496
rect 237282 270484 237288 270496
rect 233200 270456 237288 270484
rect 233200 270444 233206 270456
rect 237282 270444 237288 270456
rect 237340 270444 237346 270496
rect 237484 270484 237512 270592
rect 428458 270580 428464 270632
rect 428516 270620 428522 270632
rect 466638 270620 466644 270632
rect 428516 270592 466644 270620
rect 428516 270580 428522 270592
rect 466638 270580 466644 270592
rect 466696 270580 466702 270632
rect 477494 270580 477500 270632
rect 477552 270620 477558 270632
rect 538858 270620 538864 270632
rect 477552 270592 538864 270620
rect 477552 270580 477558 270592
rect 538858 270580 538864 270592
rect 538916 270580 538922 270632
rect 539060 270620 539088 270728
rect 540514 270716 540520 270768
rect 540572 270756 540578 270768
rect 543550 270756 543556 270768
rect 540572 270728 543556 270756
rect 540572 270716 540578 270728
rect 543550 270716 543556 270728
rect 543608 270716 543614 270768
rect 543688 270716 543694 270768
rect 543746 270756 543752 270768
rect 607306 270756 607312 270768
rect 543746 270728 607312 270756
rect 543746 270716 543752 270728
rect 607306 270716 607312 270728
rect 607364 270716 607370 270768
rect 552658 270620 552664 270632
rect 539060 270592 552664 270620
rect 552658 270580 552664 270592
rect 552716 270580 552722 270632
rect 252002 270484 252008 270496
rect 237484 270456 252008 270484
rect 252002 270444 252008 270456
rect 252060 270444 252066 270496
rect 292850 270444 292856 270496
rect 292908 270484 292914 270496
rect 296254 270484 296260 270496
rect 292908 270456 296260 270484
rect 292908 270444 292914 270456
rect 296254 270444 296260 270456
rect 296312 270444 296318 270496
rect 359734 270444 359740 270496
rect 359792 270484 359798 270496
rect 376754 270484 376760 270496
rect 359792 270456 376760 270484
rect 359792 270444 359798 270456
rect 376754 270444 376760 270456
rect 376812 270444 376818 270496
rect 377582 270444 377588 270496
rect 377640 270484 377646 270496
rect 394694 270484 394700 270496
rect 377640 270456 394700 270484
rect 377640 270444 377646 270456
rect 394694 270444 394700 270456
rect 394752 270444 394758 270496
rect 397086 270444 397092 270496
rect 397144 270484 397150 270496
rect 423674 270484 423680 270496
rect 397144 270456 423680 270484
rect 397144 270444 397150 270456
rect 423674 270444 423680 270456
rect 423732 270444 423738 270496
rect 424594 270444 424600 270496
rect 424652 270484 424658 270496
rect 476298 270484 476304 270496
rect 424652 270456 476304 270484
rect 424652 270444 424658 270456
rect 476298 270444 476304 270456
rect 476356 270444 476362 270496
rect 479242 270444 479248 270496
rect 479300 270484 479306 270496
rect 552198 270484 552204 270496
rect 479300 270456 552204 270484
rect 479300 270444 479306 270456
rect 552198 270444 552204 270456
rect 552256 270444 552262 270496
rect 552382 270444 552388 270496
rect 552440 270484 552446 270496
rect 564434 270484 564440 270496
rect 552440 270456 564440 270484
rect 552440 270444 552446 270456
rect 564434 270444 564440 270456
rect 564492 270444 564498 270496
rect 110230 270308 110236 270360
rect 110288 270348 110294 270360
rect 167914 270348 167920 270360
rect 110288 270320 167920 270348
rect 110288 270308 110294 270320
rect 167914 270308 167920 270320
rect 167972 270308 167978 270360
rect 172422 270308 172428 270360
rect 172480 270348 172486 270360
rect 208670 270348 208676 270360
rect 172480 270320 208676 270348
rect 172480 270308 172486 270320
rect 208670 270308 208676 270320
rect 208728 270308 208734 270360
rect 212442 270308 212448 270360
rect 212500 270348 212506 270360
rect 239950 270348 239956 270360
rect 212500 270320 239956 270348
rect 212500 270308 212506 270320
rect 239950 270308 239956 270320
rect 240008 270308 240014 270360
rect 253842 270308 253848 270360
rect 253900 270348 253906 270360
rect 265066 270348 265072 270360
rect 253900 270320 265072 270348
rect 253900 270308 253906 270320
rect 265066 270308 265072 270320
rect 265124 270308 265130 270360
rect 291654 270308 291660 270360
rect 291712 270348 291718 270360
rect 295518 270348 295524 270360
rect 291712 270320 295524 270348
rect 291712 270308 291718 270320
rect 295518 270308 295524 270320
rect 295576 270308 295582 270360
rect 348418 270308 348424 270360
rect 348476 270348 348482 270360
rect 363046 270348 363052 270360
rect 348476 270320 363052 270348
rect 348476 270308 348482 270320
rect 363046 270308 363052 270320
rect 363104 270308 363110 270360
rect 364978 270308 364984 270360
rect 365036 270348 365042 270360
rect 390554 270348 390560 270360
rect 365036 270320 390560 270348
rect 365036 270308 365042 270320
rect 390554 270308 390560 270320
rect 390612 270308 390618 270360
rect 392302 270308 392308 270360
rect 392360 270348 392366 270360
rect 429378 270348 429384 270360
rect 392360 270320 429384 270348
rect 392360 270308 392366 270320
rect 429378 270308 429384 270320
rect 429436 270308 429442 270360
rect 429562 270308 429568 270360
rect 429620 270348 429626 270360
rect 483106 270348 483112 270360
rect 429620 270320 483112 270348
rect 429620 270308 429626 270320
rect 483106 270308 483112 270320
rect 483164 270308 483170 270360
rect 486694 270308 486700 270360
rect 486752 270348 486758 270360
rect 490374 270348 490380 270360
rect 486752 270320 490380 270348
rect 486752 270308 486758 270320
rect 490374 270308 490380 270320
rect 490432 270308 490438 270360
rect 490558 270308 490564 270360
rect 490616 270348 490622 270360
rect 560294 270348 560300 270360
rect 490616 270320 560300 270348
rect 490616 270308 490622 270320
rect 560294 270308 560300 270320
rect 560352 270308 560358 270360
rect 316954 270240 316960 270292
rect 317012 270280 317018 270292
rect 321554 270280 321560 270292
rect 317012 270252 321560 270280
rect 317012 270240 317018 270252
rect 321554 270240 321560 270252
rect 321612 270240 321618 270292
rect 339310 270240 339316 270292
rect 339368 270280 339374 270292
rect 341518 270280 341524 270292
rect 339368 270252 341524 270280
rect 339368 270240 339374 270252
rect 341518 270240 341524 270252
rect 341576 270240 341582 270292
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 166902 270172 166908 270224
rect 166960 270212 166966 270224
rect 207382 270212 207388 270224
rect 166960 270184 207388 270212
rect 166960 270172 166966 270184
rect 207382 270172 207388 270184
rect 207440 270172 207446 270224
rect 213822 270172 213828 270224
rect 213880 270212 213886 270224
rect 240502 270212 240508 270224
rect 213880 270184 240508 270212
rect 213880 270172 213886 270184
rect 240502 270172 240508 270184
rect 240560 270172 240566 270224
rect 249610 270172 249616 270224
rect 249668 270212 249674 270224
rect 263318 270212 263324 270224
rect 249668 270184 263324 270212
rect 249668 270172 249674 270184
rect 263318 270172 263324 270184
rect 263376 270172 263382 270224
rect 269206 270172 269212 270224
rect 269264 270212 269270 270224
rect 279694 270212 279700 270224
rect 269264 270184 279700 270212
rect 269264 270172 269270 270184
rect 279694 270172 279700 270184
rect 279752 270172 279758 270224
rect 321922 270172 321928 270224
rect 321980 270212 321986 270224
rect 328454 270212 328460 270224
rect 321980 270184 328460 270212
rect 321980 270172 321986 270184
rect 328454 270172 328460 270184
rect 328512 270172 328518 270224
rect 341794 270172 341800 270224
rect 341852 270212 341858 270224
rect 357434 270212 357440 270224
rect 341852 270184 357440 270212
rect 341852 270172 341858 270184
rect 357434 270172 357440 270184
rect 357492 270172 357498 270224
rect 369394 270172 369400 270224
rect 369452 270212 369458 270224
rect 396074 270212 396080 270224
rect 369452 270184 396080 270212
rect 369452 270172 369458 270184
rect 396074 270172 396080 270184
rect 396132 270172 396138 270224
rect 403066 270172 403072 270224
rect 403124 270212 403130 270224
rect 444374 270212 444380 270224
rect 403124 270184 444380 270212
rect 403124 270172 403130 270184
rect 444374 270172 444380 270184
rect 444432 270172 444438 270224
rect 446950 270172 446956 270224
rect 447008 270212 447014 270224
rect 504174 270212 504180 270224
rect 447008 270184 504180 270212
rect 447008 270172 447014 270184
rect 504174 270172 504180 270184
rect 504232 270172 504238 270224
rect 504358 270172 504364 270224
rect 504416 270212 504422 270224
rect 504416 270184 528692 270212
rect 504416 270172 504422 270184
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 528664 270144 528692 270184
rect 528922 270172 528928 270224
rect 528980 270212 528986 270224
rect 533522 270212 533528 270224
rect 528980 270184 533528 270212
rect 528980 270172 528986 270184
rect 533522 270172 533528 270184
rect 533580 270172 533586 270224
rect 533982 270172 533988 270224
rect 534040 270212 534046 270224
rect 626534 270212 626540 270224
rect 534040 270184 626540 270212
rect 534040 270172 534046 270184
rect 626534 270172 626540 270184
rect 626592 270172 626598 270224
rect 528664 270116 528784 270144
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 146662 270036 146668 270088
rect 146720 270076 146726 270088
rect 151354 270076 151360 270088
rect 146720 270048 151360 270076
rect 146720 270036 146726 270048
rect 151354 270036 151360 270048
rect 151412 270036 151418 270088
rect 153838 270076 153844 270088
rect 151786 270048 153844 270076
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 142614 269940 142620 269952
rect 75880 269912 142620 269940
rect 75880 269900 75886 269912
rect 142614 269900 142620 269912
rect 142672 269900 142678 269952
rect 143350 269900 143356 269952
rect 143408 269940 143414 269952
rect 151786 269940 151814 270048
rect 153838 270036 153844 270048
rect 153896 270036 153902 270088
rect 159910 270036 159916 270088
rect 159968 270076 159974 270088
rect 202690 270076 202696 270088
rect 159968 270048 202696 270076
rect 159968 270036 159974 270048
rect 202690 270036 202696 270048
rect 202748 270036 202754 270088
rect 205542 270036 205548 270088
rect 205600 270076 205606 270088
rect 234982 270076 234988 270088
rect 205600 270048 234988 270076
rect 205600 270036 205606 270048
rect 234982 270036 234988 270048
rect 235040 270036 235046 270088
rect 239766 270036 239772 270088
rect 239824 270076 239830 270088
rect 253198 270076 253204 270088
rect 239824 270048 253204 270076
rect 239824 270036 239830 270048
rect 253198 270036 253204 270048
rect 253256 270036 253262 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 323578 270036 323584 270088
rect 323636 270076 323642 270088
rect 331214 270076 331220 270088
rect 323636 270048 331220 270076
rect 323636 270036 323642 270048
rect 331214 270036 331220 270048
rect 331272 270036 331278 270088
rect 354214 270036 354220 270088
rect 354272 270076 354278 270088
rect 375374 270076 375380 270088
rect 354272 270048 375380 270076
rect 354272 270036 354278 270048
rect 375374 270036 375380 270048
rect 375432 270036 375438 270088
rect 376570 270036 376576 270088
rect 376628 270076 376634 270088
rect 404262 270076 404268 270088
rect 376628 270048 404268 270076
rect 376628 270036 376634 270048
rect 404262 270036 404268 270048
rect 404320 270036 404326 270088
rect 417142 270036 417148 270088
rect 417200 270076 417206 270088
rect 465074 270076 465080 270088
rect 417200 270048 465080 270076
rect 417200 270036 417206 270048
rect 465074 270036 465080 270048
rect 465132 270036 465138 270088
rect 465994 270036 466000 270088
rect 466052 270076 466058 270088
rect 528462 270076 528468 270088
rect 466052 270048 528468 270076
rect 466052 270036 466058 270048
rect 528462 270036 528468 270048
rect 528520 270036 528526 270088
rect 528756 270076 528784 270116
rect 538858 270076 538864 270088
rect 528756 270048 538864 270076
rect 538858 270036 538864 270048
rect 538916 270036 538922 270088
rect 540974 270036 540980 270088
rect 541032 270076 541038 270088
rect 541802 270076 541808 270088
rect 541032 270048 541808 270076
rect 541032 270036 541038 270048
rect 541802 270036 541808 270048
rect 541860 270036 541866 270088
rect 541986 270036 541992 270088
rect 542044 270076 542050 270088
rect 633618 270076 633624 270088
rect 542044 270048 633624 270076
rect 542044 270036 542050 270048
rect 633618 270036 633624 270048
rect 633676 270036 633682 270088
rect 143408 269912 151814 269940
rect 143408 269900 143414 269912
rect 154482 269900 154488 269952
rect 154540 269940 154546 269952
rect 198182 269940 198188 269952
rect 154540 269912 198188 269940
rect 154540 269900 154546 269912
rect 198182 269900 198188 269912
rect 198240 269900 198246 269952
rect 198642 269900 198648 269952
rect 198700 269940 198706 269952
rect 230014 269940 230020 269952
rect 198700 269912 230020 269940
rect 198700 269900 198706 269912
rect 230014 269900 230020 269912
rect 230072 269900 230078 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 252370 269940 252376 269952
rect 230440 269912 252376 269940
rect 230440 269900 230446 269912
rect 252370 269900 252376 269912
rect 252428 269900 252434 269952
rect 258442 269900 258448 269952
rect 258500 269940 258506 269952
rect 272242 269940 272248 269952
rect 258500 269912 272248 269940
rect 258500 269900 258506 269912
rect 272242 269900 272248 269912
rect 272300 269900 272306 269952
rect 273070 269900 273076 269952
rect 273128 269940 273134 269952
rect 282178 269940 282184 269952
rect 273128 269912 282184 269940
rect 273128 269900 273134 269912
rect 282178 269900 282184 269912
rect 282236 269900 282242 269952
rect 286778 269900 286784 269952
rect 286836 269940 286842 269952
rect 292114 269940 292120 269952
rect 286836 269912 292120 269940
rect 286836 269900 286842 269912
rect 292114 269900 292120 269912
rect 292172 269900 292178 269952
rect 331674 269900 331680 269952
rect 331732 269940 331738 269952
rect 336734 269940 336740 269952
rect 331732 269912 336740 269940
rect 331732 269900 331738 269912
rect 336734 269900 336740 269912
rect 336792 269900 336798 269952
rect 347590 269900 347596 269952
rect 347648 269940 347654 269952
rect 365714 269940 365720 269952
rect 347648 269912 365720 269940
rect 347648 269900 347654 269912
rect 365714 269900 365720 269912
rect 365772 269900 365778 269952
rect 372338 269900 372344 269952
rect 372396 269940 372402 269952
rect 401778 269940 401784 269952
rect 372396 269912 401784 269940
rect 372396 269900 372402 269912
rect 401778 269900 401784 269912
rect 401836 269900 401842 269952
rect 413002 269900 413008 269952
rect 413060 269940 413066 269952
rect 459554 269940 459560 269952
rect 413060 269912 459560 269940
rect 413060 269900 413066 269912
rect 459554 269900 459560 269912
rect 459612 269900 459618 269952
rect 461854 269900 461860 269952
rect 461912 269940 461918 269952
rect 528646 269940 528652 269952
rect 461912 269912 528652 269940
rect 461912 269900 461918 269912
rect 528646 269900 528652 269912
rect 528704 269900 528710 269952
rect 529750 269900 529756 269952
rect 529808 269940 529814 269952
rect 530762 269940 530768 269952
rect 529808 269912 530768 269940
rect 529808 269900 529814 269912
rect 530762 269900 530768 269912
rect 530820 269900 530826 269952
rect 530946 269900 530952 269952
rect 531004 269940 531010 269952
rect 532970 269940 532976 269952
rect 531004 269912 532976 269940
rect 531004 269900 531010 269912
rect 532970 269900 532976 269912
rect 533028 269900 533034 269952
rect 536558 269900 536564 269952
rect 536616 269940 536622 269952
rect 630674 269940 630680 269952
rect 536616 269912 630680 269940
rect 536616 269900 536622 269912
rect 630674 269900 630680 269912
rect 630732 269900 630738 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 139946 269764 139952 269816
rect 140004 269804 140010 269816
rect 181162 269804 181168 269816
rect 140004 269776 181168 269804
rect 140004 269764 140010 269776
rect 181162 269764 181168 269776
rect 181220 269764 181226 269816
rect 182082 269764 182088 269816
rect 182140 269804 182146 269816
rect 186958 269804 186964 269816
rect 182140 269776 186964 269804
rect 182140 269764 182146 269776
rect 186958 269764 186964 269776
rect 187016 269764 187022 269816
rect 187326 269764 187332 269816
rect 187384 269804 187390 269816
rect 191926 269804 191932 269816
rect 187384 269776 191932 269804
rect 187384 269764 187390 269776
rect 191926 269764 191932 269776
rect 191984 269764 191990 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 84102 269628 84108 269680
rect 84160 269668 84166 269680
rect 119798 269668 119804 269680
rect 84160 269640 119804 269668
rect 84160 269628 84166 269640
rect 119798 269628 119804 269640
rect 119856 269628 119862 269680
rect 173710 269668 173716 269680
rect 122806 269640 173716 269668
rect 119062 269492 119068 269544
rect 119120 269532 119126 269544
rect 122806 269532 122834 269640
rect 173710 269628 173716 269640
rect 173768 269628 173774 269680
rect 184750 269628 184756 269680
rect 184808 269668 184814 269680
rect 213822 269668 213828 269680
rect 184808 269640 213828 269668
rect 184808 269628 184814 269640
rect 213822 269628 213828 269640
rect 213880 269628 213886 269680
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 251450 269764 251456 269816
rect 251508 269804 251514 269816
rect 267274 269804 267280 269816
rect 251508 269776 267280 269804
rect 251508 269764 251514 269776
rect 267274 269764 267280 269776
rect 267332 269764 267338 269816
rect 270310 269764 270316 269816
rect 270368 269804 270374 269816
rect 280522 269804 280528 269816
rect 270368 269776 280528 269804
rect 270368 269764 270374 269776
rect 280522 269764 280528 269776
rect 280580 269764 280586 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318794 269804 318800 269816
rect 314528 269776 318800 269804
rect 314528 269764 314534 269776
rect 318794 269764 318800 269776
rect 318852 269764 318858 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335906 269804 335912 269816
rect 326948 269776 335912 269804
rect 326948 269764 326954 269776
rect 335906 269764 335912 269776
rect 335964 269764 335970 269816
rect 336826 269764 336832 269816
rect 336884 269804 336890 269816
rect 350534 269804 350540 269816
rect 336884 269776 350540 269804
rect 336884 269764 336890 269776
rect 350534 269764 350540 269776
rect 350592 269764 350598 269816
rect 356698 269764 356704 269816
rect 356756 269804 356762 269816
rect 378134 269804 378140 269816
rect 356756 269776 378140 269804
rect 356756 269764 356762 269776
rect 378134 269764 378140 269776
rect 378192 269764 378198 269816
rect 385678 269764 385684 269816
rect 385736 269804 385742 269816
rect 419534 269804 419540 269816
rect 385736 269776 419540 269804
rect 385736 269764 385742 269776
rect 419534 269764 419540 269776
rect 419592 269764 419598 269816
rect 419994 269764 420000 269816
rect 420052 269804 420058 269816
rect 468018 269804 468024 269816
rect 420052 269776 468024 269804
rect 420052 269764 420058 269776
rect 468018 269764 468024 269776
rect 468076 269764 468082 269816
rect 470962 269764 470968 269816
rect 471020 269804 471026 269816
rect 537478 269804 537484 269816
rect 471020 269776 537484 269804
rect 471020 269764 471026 269776
rect 537478 269764 537484 269776
rect 537536 269764 537542 269816
rect 538858 269764 538864 269816
rect 538916 269804 538922 269816
rect 552290 269804 552296 269816
rect 538916 269776 552296 269804
rect 538916 269764 538922 269776
rect 552290 269764 552296 269776
rect 552348 269764 552354 269816
rect 552474 269764 552480 269816
rect 552532 269804 552538 269816
rect 641898 269804 641904 269816
rect 552532 269776 641904 269804
rect 552532 269764 552538 269776
rect 641898 269764 641904 269776
rect 641956 269764 641962 269816
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 253198 269628 253204 269680
rect 253256 269668 253262 269680
rect 258166 269668 258172 269680
rect 253256 269640 258172 269668
rect 253256 269628 253262 269640
rect 258166 269628 258172 269640
rect 258224 269628 258230 269680
rect 329650 269628 329656 269680
rect 329708 269668 329714 269680
rect 339494 269668 339500 269680
rect 329708 269640 339500 269668
rect 329708 269628 329714 269640
rect 339494 269628 339500 269640
rect 339552 269628 339558 269680
rect 351638 269628 351644 269680
rect 351696 269668 351702 269680
rect 364334 269668 364340 269680
rect 351696 269640 364340 269668
rect 351696 269628 351702 269640
rect 364334 269628 364340 269640
rect 364392 269628 364398 269680
rect 384022 269628 384028 269680
rect 384080 269668 384086 269680
rect 388162 269668 388168 269680
rect 384080 269640 388168 269668
rect 384080 269628 384086 269640
rect 388162 269628 388168 269640
rect 388220 269628 388226 269680
rect 394694 269628 394700 269680
rect 394752 269668 394758 269680
rect 416774 269668 416780 269680
rect 394752 269640 416780 269668
rect 394752 269628 394758 269640
rect 416774 269628 416780 269640
rect 416832 269628 416838 269680
rect 427354 269628 427360 269680
rect 427412 269668 427418 269680
rect 478874 269668 478880 269680
rect 427412 269640 478880 269668
rect 427412 269628 427418 269640
rect 478874 269628 478880 269640
rect 478932 269628 478938 269680
rect 484210 269628 484216 269680
rect 484268 269668 484274 269680
rect 490558 269668 490564 269680
rect 484268 269640 490564 269668
rect 484268 269628 484274 269640
rect 490558 269628 490564 269640
rect 490616 269628 490622 269680
rect 490742 269628 490748 269680
rect 490800 269668 490806 269680
rect 504358 269668 504364 269680
rect 490800 269640 504364 269668
rect 490800 269628 490806 269640
rect 504358 269628 504364 269640
rect 504416 269628 504422 269680
rect 504542 269628 504548 269680
rect 504600 269668 504606 269680
rect 553026 269668 553032 269680
rect 504600 269640 553032 269668
rect 504600 269628 504606 269640
rect 553026 269628 553032 269640
rect 553084 269628 553090 269680
rect 558914 269628 558920 269680
rect 558972 269668 558978 269680
rect 572714 269668 572720 269680
rect 558972 269640 572720 269668
rect 558972 269628 558978 269640
rect 572714 269628 572720 269640
rect 572772 269628 572778 269680
rect 119120 269504 122834 269532
rect 119120 269492 119126 269504
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 187326 269532 187332 269544
rect 183520 269504 187332 269532
rect 183520 269492 183526 269504
rect 187326 269492 187332 269504
rect 187384 269492 187390 269544
rect 208302 269492 208308 269544
rect 208360 269532 208366 269544
rect 230750 269532 230756 269544
rect 208360 269504 230756 269532
rect 208360 269492 208366 269504
rect 230750 269492 230756 269504
rect 230808 269492 230814 269544
rect 401594 269492 401600 269544
rect 401652 269532 401658 269544
rect 430574 269532 430580 269544
rect 401652 269504 430580 269532
rect 401652 269492 401658 269504
rect 430574 269492 430580 269504
rect 430632 269492 430638 269544
rect 449894 269492 449900 269544
rect 449952 269532 449958 269544
rect 471974 269532 471980 269544
rect 449952 269504 471980 269532
rect 449952 269492 449958 269504
rect 471974 269492 471980 269504
rect 472032 269492 472038 269544
rect 474274 269492 474280 269544
rect 474332 269532 474338 269544
rect 474332 269504 537340 269532
rect 474332 269492 474338 269504
rect 118602 269356 118608 269408
rect 118660 269396 118666 269408
rect 166902 269396 166908 269408
rect 118660 269368 166908 269396
rect 118660 269356 118666 269368
rect 166902 269356 166908 269368
rect 166960 269356 166966 269408
rect 335630 269356 335636 269408
rect 335688 269396 335694 269408
rect 343818 269396 343824 269408
rect 335688 269368 343824 269396
rect 335688 269356 335694 269368
rect 343818 269356 343824 269368
rect 343876 269356 343882 269408
rect 404354 269356 404360 269408
rect 404412 269396 404418 269408
rect 426618 269396 426624 269408
rect 404412 269368 426624 269396
rect 404412 269356 404418 269368
rect 426618 269356 426624 269368
rect 426676 269356 426682 269408
rect 457714 269356 457720 269408
rect 457772 269396 457778 269408
rect 471790 269396 471796 269408
rect 457772 269368 471796 269396
rect 457772 269356 457778 269368
rect 471790 269356 471796 269368
rect 471848 269356 471854 269408
rect 476758 269356 476764 269408
rect 476816 269396 476822 269408
rect 537312 269396 537340 269504
rect 537478 269492 537484 269544
rect 537536 269532 537542 269544
rect 540974 269532 540980 269544
rect 537536 269504 540980 269532
rect 537536 269492 537542 269504
rect 540974 269492 540980 269504
rect 541032 269492 541038 269544
rect 541342 269492 541348 269544
rect 541400 269532 541406 269544
rect 552382 269532 552388 269544
rect 541400 269504 552388 269532
rect 541400 269492 541406 269504
rect 552382 269492 552388 269504
rect 552440 269492 552446 269544
rect 568574 269532 568580 269544
rect 552768 269504 568580 269532
rect 552768 269464 552796 269504
rect 568574 269492 568580 269504
rect 568632 269492 568638 269544
rect 552584 269436 552796 269464
rect 546218 269396 546224 269408
rect 476816 269368 537248 269396
rect 537312 269368 546224 269396
rect 476816 269356 476822 269368
rect 136818 269220 136824 269272
rect 136876 269260 136882 269272
rect 182174 269260 182180 269272
rect 136876 269232 182180 269260
rect 136876 269220 136882 269232
rect 182174 269220 182180 269232
rect 182232 269220 182238 269272
rect 264882 269220 264888 269272
rect 264940 269260 264946 269272
rect 269114 269260 269120 269272
rect 264940 269232 269120 269260
rect 264940 269220 264946 269232
rect 269114 269220 269120 269232
rect 269172 269220 269178 269272
rect 321094 269220 321100 269272
rect 321152 269260 321158 269272
rect 327902 269260 327908 269272
rect 321152 269232 327908 269260
rect 321152 269220 321158 269232
rect 327902 269220 327908 269232
rect 327960 269220 327966 269272
rect 468754 269220 468760 269272
rect 468812 269260 468818 269272
rect 537018 269260 537024 269272
rect 468812 269232 537024 269260
rect 468812 269220 468818 269232
rect 537018 269220 537024 269232
rect 537076 269220 537082 269272
rect 537220 269260 537248 269368
rect 546218 269356 546224 269368
rect 546276 269356 546282 269408
rect 546402 269356 546408 269408
rect 546460 269396 546466 269408
rect 551922 269396 551928 269408
rect 546460 269368 551928 269396
rect 546460 269356 546466 269368
rect 551922 269356 551928 269368
rect 551980 269356 551986 269408
rect 552584 269396 552612 269436
rect 552124 269368 552612 269396
rect 549438 269260 549444 269272
rect 537220 269232 549444 269260
rect 549438 269220 549444 269232
rect 549496 269220 549502 269272
rect 549622 269220 549628 269272
rect 549680 269260 549686 269272
rect 552124 269260 552152 269368
rect 553026 269356 553032 269408
rect 553084 269396 553090 269408
rect 557534 269396 557540 269408
rect 553084 269368 557540 269396
rect 553084 269356 553090 269368
rect 557534 269356 557540 269368
rect 557592 269356 557598 269408
rect 549680 269232 552152 269260
rect 549680 269220 549686 269232
rect 552290 269220 552296 269272
rect 552348 269260 552354 269272
rect 607582 269260 607588 269272
rect 552348 269232 607588 269260
rect 552348 269220 552354 269232
rect 607582 269220 607588 269232
rect 607640 269220 607646 269272
rect 282730 269084 282736 269136
rect 282788 269124 282794 269136
rect 288802 269124 288808 269136
rect 282788 269096 288808 269124
rect 282788 269084 282794 269096
rect 288802 269084 288808 269096
rect 288860 269084 288866 269136
rect 295334 269084 295340 269136
rect 295392 269124 295398 269136
rect 297542 269124 297548 269136
rect 295392 269096 297548 269124
rect 295392 269084 295398 269096
rect 297542 269084 297548 269096
rect 297600 269084 297606 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 434438 269084 434444 269136
rect 434496 269124 434502 269136
rect 489914 269124 489920 269136
rect 434496 269096 489920 269124
rect 434496 269084 434502 269096
rect 489914 269084 489920 269096
rect 489972 269084 489978 269136
rect 108942 269016 108948 269068
rect 109000 269056 109006 269068
rect 166258 269056 166264 269068
rect 109000 269028 166264 269056
rect 109000 269016 109006 269028
rect 166258 269016 166264 269028
rect 166316 269016 166322 269068
rect 185578 269016 185584 269068
rect 185636 269056 185642 269068
rect 196894 269056 196900 269068
rect 185636 269028 196900 269056
rect 185636 269016 185642 269028
rect 196894 269016 196900 269028
rect 196952 269016 196958 269068
rect 251082 269016 251088 269068
rect 251140 269056 251146 269068
rect 256510 269056 256516 269068
rect 251140 269028 256516 269056
rect 251140 269016 251146 269028
rect 256510 269016 256516 269028
rect 256568 269016 256574 269068
rect 422294 269056 422300 269068
rect 412606 269028 422300 269056
rect 86862 268880 86868 268932
rect 86920 268920 86926 268932
rect 144730 268920 144736 268932
rect 86920 268892 144736 268920
rect 86920 268880 86926 268892
rect 144730 268880 144736 268892
rect 144788 268880 144794 268932
rect 179322 268880 179328 268932
rect 179380 268920 179386 268932
rect 215938 268920 215944 268932
rect 179380 268892 215944 268920
rect 179380 268880 179386 268892
rect 215938 268880 215944 268892
rect 215996 268880 216002 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 400582 268920 400588 268932
rect 382424 268892 400588 268920
rect 382424 268880 382430 268892
rect 400582 268880 400588 268892
rect 400640 268880 400646 268932
rect 102502 268744 102508 268796
rect 102560 268784 102566 268796
rect 162946 268784 162952 268796
rect 102560 268756 162952 268784
rect 102560 268744 102566 268756
rect 162946 268744 162952 268756
rect 163004 268744 163010 268796
rect 163130 268744 163136 268796
rect 163188 268784 163194 268796
rect 203518 268784 203524 268796
rect 163188 268756 203524 268784
rect 163188 268744 163194 268756
rect 203518 268744 203524 268756
rect 203576 268744 203582 268796
rect 203978 268744 203984 268796
rect 204036 268784 204042 268796
rect 227714 268784 227720 268796
rect 204036 268756 227720 268784
rect 204036 268744 204042 268756
rect 227714 268744 227720 268756
rect 227772 268744 227778 268796
rect 227898 268744 227904 268796
rect 227956 268784 227962 268796
rect 250714 268784 250720 268796
rect 227956 268756 250720 268784
rect 227956 268744 227962 268756
rect 250714 268744 250720 268756
rect 250772 268744 250778 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 412606 268784 412634 269028
rect 422294 269016 422300 269028
rect 422352 269016 422358 269068
rect 503254 269016 503260 269068
rect 503312 269056 503318 269068
rect 581454 269056 581460 269068
rect 503312 269028 581460 269056
rect 503312 269016 503318 269028
rect 581454 269016 581460 269028
rect 581512 269016 581518 269068
rect 581638 269016 581644 269068
rect 581696 269056 581702 269068
rect 584122 269056 584128 269068
rect 581696 269028 584128 269056
rect 581696 269016 581702 269028
rect 584122 269016 584128 269028
rect 584180 269016 584186 269068
rect 590654 269016 590660 269068
rect 590712 269056 590718 269068
rect 590712 269028 596174 269056
rect 590712 269016 590718 269028
rect 418982 268880 418988 268932
rect 419040 268920 419046 268932
rect 440234 268920 440240 268932
rect 419040 268892 440240 268920
rect 419040 268880 419046 268892
rect 440234 268880 440240 268892
rect 440292 268880 440298 268932
rect 443638 268880 443644 268932
rect 443696 268920 443702 268932
rect 502426 268920 502432 268932
rect 443696 268892 502432 268920
rect 443696 268880 443702 268892
rect 502426 268880 502432 268892
rect 502484 268880 502490 268932
rect 503438 268880 503444 268932
rect 503496 268920 503502 268932
rect 505094 268920 505100 268932
rect 503496 268892 505100 268920
rect 503496 268880 503502 268892
rect 505094 268880 505100 268892
rect 505152 268880 505158 268932
rect 508498 268880 508504 268932
rect 508556 268920 508562 268932
rect 594794 268920 594800 268932
rect 508556 268892 594800 268920
rect 508556 268880 508562 268892
rect 594794 268880 594800 268892
rect 594852 268880 594858 268932
rect 387392 268756 412634 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268796
rect 422352 268784 422358 268796
rect 436094 268784 436100 268796
rect 422352 268756 436100 268784
rect 422352 268744 422358 268756
rect 436094 268744 436100 268756
rect 436152 268744 436158 268796
rect 441154 268744 441160 268796
rect 441212 268784 441218 268796
rect 499574 268784 499580 268796
rect 441212 268756 499580 268784
rect 441212 268744 441218 268756
rect 499574 268744 499580 268756
rect 499632 268744 499638 268796
rect 500678 268744 500684 268796
rect 500736 268784 500742 268796
rect 581270 268784 581276 268796
rect 500736 268756 581276 268784
rect 500736 268744 500742 268756
rect 581270 268744 581276 268756
rect 581328 268744 581334 268796
rect 581638 268744 581644 268796
rect 581696 268784 581702 268796
rect 596146 268784 596174 269028
rect 598842 268784 598848 268796
rect 581696 268756 590884 268784
rect 596146 268756 598848 268784
rect 581696 268744 581702 268756
rect 590856 268716 590884 268756
rect 598842 268744 598848 268756
rect 598900 268744 598906 268796
rect 590856 268688 590976 268716
rect 99282 268608 99288 268660
rect 99340 268648 99346 268660
rect 160462 268648 160468 268660
rect 99340 268620 160468 268648
rect 99340 268608 99346 268620
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 162762 268608 162768 268660
rect 162820 268648 162826 268660
rect 205174 268648 205180 268660
rect 162820 268620 205180 268648
rect 162820 268608 162826 268620
rect 205174 268608 205180 268620
rect 205232 268608 205238 268660
rect 219526 268608 219532 268660
rect 219584 268648 219590 268660
rect 244918 268648 244924 268660
rect 219584 268620 244924 268648
rect 219584 268608 219590 268620
rect 244918 268608 244924 268620
rect 244976 268608 244982 268660
rect 363046 268608 363052 268660
rect 363104 268648 363110 268660
rect 386414 268648 386420 268660
rect 363104 268620 386420 268648
rect 363104 268608 363110 268620
rect 386414 268608 386420 268620
rect 386472 268608 386478 268660
rect 400582 268608 400588 268660
rect 400640 268648 400646 268660
rect 441614 268648 441620 268660
rect 400640 268620 441620 268648
rect 400640 268608 400646 268620
rect 441614 268608 441620 268620
rect 441672 268608 441678 268660
rect 442718 268608 442724 268660
rect 442776 268648 442782 268660
rect 445754 268648 445760 268660
rect 442776 268620 445760 268648
rect 442776 268608 442782 268620
rect 445754 268608 445760 268620
rect 445812 268608 445818 268660
rect 446582 268608 446588 268660
rect 446640 268648 446646 268660
rect 503438 268648 503444 268660
rect 446640 268620 503444 268648
rect 446640 268608 446646 268620
rect 503438 268608 503444 268620
rect 503496 268608 503502 268660
rect 504174 268608 504180 268660
rect 504232 268648 504238 268660
rect 504232 268620 504588 268648
rect 504232 268608 504238 268620
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 155862 268472 155868 268524
rect 155920 268512 155926 268524
rect 200206 268512 200212 268524
rect 155920 268484 200212 268512
rect 155920 268472 155926 268484
rect 200206 268472 200212 268484
rect 200264 268472 200270 268524
rect 202966 268472 202972 268524
rect 203024 268512 203030 268524
rect 233326 268512 233332 268524
rect 203024 268484 233332 268512
rect 203024 268472 203030 268484
rect 233326 268472 233332 268484
rect 233384 268472 233390 268524
rect 245562 268472 245568 268524
rect 245620 268512 245626 268524
rect 263134 268512 263140 268524
rect 245620 268484 263140 268512
rect 245620 268472 245626 268484
rect 263134 268472 263140 268484
rect 263192 268472 263198 268524
rect 263502 268472 263508 268524
rect 263560 268512 263566 268524
rect 275554 268512 275560 268524
rect 263560 268484 275560 268512
rect 263560 268472 263566 268484
rect 275554 268472 275560 268484
rect 275612 268472 275618 268524
rect 333514 268472 333520 268524
rect 333572 268512 333578 268524
rect 345106 268512 345112 268524
rect 333572 268484 345112 268512
rect 333572 268472 333578 268484
rect 345106 268472 345112 268484
rect 345164 268472 345170 268524
rect 345934 268472 345940 268524
rect 345992 268512 345998 268524
rect 360286 268512 360292 268524
rect 345992 268484 360292 268512
rect 345992 268472 345998 268484
rect 360286 268472 360292 268484
rect 360344 268472 360350 268524
rect 361022 268472 361028 268524
rect 361080 268512 361086 268524
rect 369854 268512 369860 268524
rect 361080 268484 369860 268512
rect 361080 268472 361086 268484
rect 369854 268472 369860 268484
rect 369912 268472 369918 268524
rect 370314 268472 370320 268524
rect 370372 268512 370378 268524
rect 397454 268512 397460 268524
rect 370372 268484 397460 268512
rect 370372 268472 370378 268484
rect 397454 268472 397460 268484
rect 397512 268472 397518 268524
rect 402238 268472 402244 268524
rect 402296 268512 402302 268524
rect 443270 268512 443276 268524
rect 402296 268484 443276 268512
rect 402296 268472 402302 268484
rect 443270 268472 443276 268484
rect 443328 268472 443334 268524
rect 448606 268472 448612 268524
rect 448664 268512 448670 268524
rect 504358 268512 504364 268524
rect 448664 268484 504364 268512
rect 448664 268472 448670 268484
rect 504358 268472 504364 268484
rect 504416 268472 504422 268524
rect 504560 268512 504588 268620
rect 506106 268608 506112 268660
rect 506164 268648 506170 268660
rect 514018 268648 514024 268660
rect 506164 268620 514024 268648
rect 506164 268608 506170 268620
rect 514018 268608 514024 268620
rect 514076 268608 514082 268660
rect 514202 268608 514208 268660
rect 514260 268648 514266 268660
rect 590654 268648 590660 268660
rect 514260 268620 590660 268648
rect 514260 268608 514266 268620
rect 590654 268608 590660 268620
rect 590712 268608 590718 268660
rect 590948 268648 590976 268688
rect 608686 268648 608692 268660
rect 590948 268620 608692 268648
rect 608686 268608 608692 268620
rect 608744 268608 608750 268660
rect 504560 268484 519124 268512
rect 66254 268336 66260 268388
rect 66312 268376 66318 268388
rect 137278 268376 137284 268388
rect 66312 268348 137284 268376
rect 66312 268336 66318 268348
rect 137278 268336 137284 268348
rect 137336 268336 137342 268388
rect 147582 268336 147588 268388
rect 147640 268376 147646 268388
rect 193582 268376 193588 268388
rect 147640 268348 193588 268376
rect 147640 268336 147646 268348
rect 193582 268336 193588 268348
rect 193640 268336 193646 268388
rect 197262 268336 197268 268388
rect 197320 268376 197326 268388
rect 229186 268376 229192 268388
rect 197320 268348 229192 268376
rect 197320 268336 197326 268348
rect 229186 268336 229192 268348
rect 229244 268336 229250 268388
rect 233694 268336 233700 268388
rect 233752 268376 233758 268388
rect 254854 268376 254860 268388
rect 233752 268348 254860 268376
rect 233752 268336 233758 268348
rect 254854 268336 254860 268348
rect 254912 268336 254918 268388
rect 255314 268336 255320 268388
rect 255372 268376 255378 268388
rect 269758 268376 269764 268388
rect 255372 268348 269764 268376
rect 255372 268336 255378 268348
rect 269758 268336 269764 268348
rect 269816 268336 269822 268388
rect 322750 268336 322756 268388
rect 322808 268376 322814 268388
rect 329834 268376 329840 268388
rect 322808 268348 329840 268376
rect 322808 268336 322814 268348
rect 329834 268336 329840 268348
rect 329892 268336 329898 268388
rect 335170 268336 335176 268388
rect 335228 268376 335234 268388
rect 347774 268376 347780 268388
rect 335228 268348 347780 268376
rect 335228 268336 335234 268348
rect 347774 268336 347780 268348
rect 347832 268336 347838 268388
rect 350074 268336 350080 268388
rect 350132 268376 350138 268388
rect 367094 268376 367100 268388
rect 350132 268348 367100 268376
rect 350132 268336 350138 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 374914 268336 374920 268388
rect 374972 268376 374978 268388
rect 404538 268376 404544 268388
rect 374972 268348 404544 268376
rect 374972 268336 374978 268348
rect 404538 268336 404544 268348
rect 404596 268336 404602 268388
rect 407206 268336 407212 268388
rect 407264 268376 407270 268388
rect 451458 268376 451464 268388
rect 407264 268348 451464 268376
rect 407264 268336 407270 268348
rect 451458 268336 451464 268348
rect 451516 268336 451522 268388
rect 461026 268336 461032 268388
rect 461084 268376 461090 268388
rect 518894 268376 518900 268388
rect 461084 268348 518900 268376
rect 461084 268336 461090 268348
rect 518894 268336 518900 268348
rect 518952 268336 518958 268388
rect 519096 268376 519124 268484
rect 519354 268472 519360 268524
rect 519412 268512 519418 268524
rect 533890 268512 533896 268524
rect 519412 268484 533896 268512
rect 519412 268472 519418 268484
rect 533890 268472 533896 268484
rect 533948 268472 533954 268524
rect 534028 268472 534034 268524
rect 534086 268512 534092 268524
rect 619634 268512 619640 268524
rect 534086 268484 619640 268512
rect 534086 268472 534092 268484
rect 619634 268472 619640 268484
rect 619692 268472 619698 268524
rect 520274 268376 520280 268388
rect 519096 268348 520280 268376
rect 520274 268336 520280 268348
rect 520332 268336 520338 268388
rect 520458 268336 520464 268388
rect 520516 268376 520522 268388
rect 526990 268376 526996 268388
rect 520516 268348 526996 268376
rect 520516 268336 520522 268348
rect 526990 268336 526996 268348
rect 527048 268336 527054 268388
rect 527174 268336 527180 268388
rect 527232 268376 527238 268388
rect 547506 268376 547512 268388
rect 527232 268348 547512 268376
rect 527232 268336 527238 268348
rect 547506 268336 547512 268348
rect 547564 268336 547570 268388
rect 547690 268336 547696 268388
rect 547748 268376 547754 268388
rect 638954 268376 638960 268388
rect 547748 268348 638960 268376
rect 547748 268336 547754 268348
rect 638954 268336 638960 268348
rect 639012 268336 639018 268388
rect 122742 268200 122748 268252
rect 122800 268240 122806 268252
rect 176194 268240 176200 268252
rect 122800 268212 176200 268240
rect 122800 268200 122806 268212
rect 176194 268200 176200 268212
rect 176252 268200 176258 268252
rect 436186 268200 436192 268252
rect 436244 268240 436250 268252
rect 436244 268212 480668 268240
rect 436244 268200 436250 268212
rect 480640 268172 480668 268212
rect 480990 268200 480996 268252
rect 481048 268240 481054 268252
rect 504174 268240 504180 268252
rect 481048 268212 504180 268240
rect 481048 268200 481054 268212
rect 504174 268200 504180 268212
rect 504232 268200 504238 268252
rect 504358 268200 504364 268252
rect 504416 268240 504422 268252
rect 509602 268240 509608 268252
rect 504416 268212 509608 268240
rect 504416 268200 504422 268212
rect 509602 268200 509608 268212
rect 509660 268200 509666 268252
rect 510706 268200 510712 268252
rect 510764 268240 510770 268252
rect 513834 268240 513840 268252
rect 510764 268212 513840 268240
rect 510764 268200 510770 268212
rect 513834 268200 513840 268212
rect 513892 268200 513898 268252
rect 514018 268200 514024 268252
rect 514076 268240 514082 268252
rect 591022 268240 591028 268252
rect 514076 268212 591028 268240
rect 514076 268200 514082 268212
rect 591022 268200 591028 268212
rect 591080 268200 591086 268252
rect 480640 268144 480760 268172
rect 133782 268064 133788 268116
rect 133840 268104 133846 268116
rect 183646 268104 183652 268116
rect 133840 268076 183652 268104
rect 133840 268064 133846 268076
rect 183646 268064 183652 268076
rect 183704 268064 183710 268116
rect 420454 268064 420460 268116
rect 420512 268104 420518 268116
rect 469030 268104 469036 268116
rect 420512 268076 469036 268104
rect 420512 268064 420518 268076
rect 469030 268064 469036 268076
rect 469088 268064 469094 268116
rect 469214 268064 469220 268116
rect 469272 268104 469278 268116
rect 480438 268104 480444 268116
rect 469272 268076 480444 268104
rect 469272 268064 469278 268076
rect 480438 268064 480444 268076
rect 480496 268064 480502 268116
rect 480732 268104 480760 268144
rect 488534 268104 488540 268116
rect 480732 268076 488540 268104
rect 488534 268064 488540 268076
rect 488592 268064 488598 268116
rect 491478 268064 491484 268116
rect 491536 268104 491542 268116
rect 494698 268104 494704 268116
rect 491536 268076 494704 268104
rect 491536 268064 491542 268076
rect 494698 268064 494704 268076
rect 494756 268064 494762 268116
rect 499114 268064 499120 268116
rect 499172 268104 499178 268116
rect 579614 268104 579620 268116
rect 499172 268076 579620 268104
rect 499172 268064 499178 268076
rect 579614 268064 579620 268076
rect 579672 268064 579678 268116
rect 581454 268064 581460 268116
rect 581512 268104 581518 268116
rect 587894 268104 587900 268116
rect 581512 268076 587900 268104
rect 581512 268064 581518 268076
rect 587894 268064 587900 268076
rect 587952 268064 587958 268116
rect 125502 267928 125508 267980
rect 125560 267968 125566 267980
rect 147582 267968 147588 267980
rect 125560 267940 147588 267968
rect 125560 267928 125566 267940
rect 147582 267928 147588 267940
rect 147640 267928 147646 267980
rect 437842 267928 437848 267980
rect 437900 267968 437906 267980
rect 468202 267968 468208 267980
rect 437900 267940 468208 267968
rect 437900 267928 437906 267940
rect 468202 267928 468208 267940
rect 468260 267928 468266 267980
rect 533890 267968 533896 267980
rect 470566 267940 533896 267968
rect 431954 267792 431960 267844
rect 432012 267832 432018 267844
rect 447134 267832 447140 267844
rect 432012 267804 447140 267832
rect 432012 267792 432018 267804
rect 447134 267792 447140 267804
rect 447192 267792 447198 267844
rect 470566 267832 470594 267940
rect 533890 267928 533896 267940
rect 533948 267928 533954 267980
rect 534028 267928 534034 267980
rect 534086 267968 534092 267980
rect 581638 267968 581644 267980
rect 534086 267940 581644 267968
rect 534086 267928 534092 267940
rect 581638 267928 581644 267940
rect 581696 267928 581702 267980
rect 467944 267804 470594 267832
rect 95878 267656 95884 267708
rect 95936 267696 95942 267708
rect 154666 267696 154672 267708
rect 95936 267668 154672 267696
rect 95936 267656 95942 267668
rect 154666 267656 154672 267668
rect 154724 267656 154730 267708
rect 162118 267656 162124 267708
rect 162176 267696 162182 267708
rect 169570 267696 169576 267708
rect 162176 267668 169576 267696
rect 162176 267656 162182 267668
rect 169570 267656 169576 267668
rect 169628 267656 169634 267708
rect 171778 267656 171784 267708
rect 171836 267696 171842 267708
rect 199378 267696 199384 267708
rect 171836 267668 199384 267696
rect 171836 267656 171842 267668
rect 199378 267656 199384 267668
rect 199436 267656 199442 267708
rect 207658 267656 207664 267708
rect 207716 267696 207722 267708
rect 213454 267696 213460 267708
rect 207716 267668 213460 267696
rect 207716 267656 207722 267668
rect 213454 267656 213460 267668
rect 213512 267656 213518 267708
rect 216122 267656 216128 267708
rect 216180 267696 216186 267708
rect 223390 267696 223396 267708
rect 216180 267668 223396 267696
rect 216180 267656 216186 267668
rect 223390 267656 223396 267668
rect 223448 267656 223454 267708
rect 368198 267656 368204 267708
rect 368256 267696 368262 267708
rect 377582 267696 377588 267708
rect 368256 267668 377588 267696
rect 368256 267656 368262 267668
rect 377582 267656 377588 267668
rect 377640 267656 377646 267708
rect 388162 267656 388168 267708
rect 388220 267696 388226 267708
rect 397086 267696 397092 267708
rect 388220 267668 397092 267696
rect 388220 267656 388226 267668
rect 397086 267656 397092 267668
rect 397144 267656 397150 267708
rect 398098 267656 398104 267708
rect 398156 267696 398162 267708
rect 421742 267696 421748 267708
rect 398156 267668 421748 267696
rect 398156 267656 398162 267668
rect 421742 267656 421748 267668
rect 421800 267656 421806 267708
rect 430390 267656 430396 267708
rect 430448 267696 430454 267708
rect 460014 267696 460020 267708
rect 430448 267668 460020 267696
rect 430448 267656 430454 267668
rect 460014 267656 460020 267668
rect 460072 267656 460078 267708
rect 460198 267656 460204 267708
rect 460256 267696 460262 267708
rect 465534 267696 465540 267708
rect 460256 267668 465540 267696
rect 460256 267656 460262 267668
rect 465534 267656 465540 267668
rect 465592 267656 465598 267708
rect 466822 267656 466828 267708
rect 466880 267696 466886 267708
rect 467944 267696 467972 267804
rect 489178 267792 489184 267844
rect 489236 267832 489242 267844
rect 567654 267832 567660 267844
rect 489236 267804 567660 267832
rect 489236 267792 489242 267804
rect 567654 267792 567660 267804
rect 567712 267792 567718 267844
rect 579614 267792 579620 267844
rect 579672 267832 579678 267844
rect 582374 267832 582380 267844
rect 579672 267804 582380 267832
rect 579672 267792 579678 267804
rect 582374 267792 582380 267804
rect 582432 267792 582438 267844
rect 466880 267668 467972 267696
rect 466880 267656 466886 267668
rect 470134 267656 470140 267708
rect 470192 267696 470198 267708
rect 518802 267696 518808 267708
rect 470192 267668 518808 267696
rect 470192 267656 470198 267668
rect 518802 267656 518808 267668
rect 518860 267656 518866 267708
rect 518986 267656 518992 267708
rect 519044 267696 519050 267708
rect 533982 267696 533988 267708
rect 519044 267668 533988 267696
rect 519044 267656 519050 267668
rect 533982 267656 533988 267668
rect 534040 267656 534046 267708
rect 534166 267656 534172 267708
rect 534224 267696 534230 267708
rect 537018 267696 537024 267708
rect 534224 267668 537024 267696
rect 534224 267656 534230 267668
rect 537018 267656 537024 267668
rect 537076 267656 537082 267708
rect 537202 267656 537208 267708
rect 537260 267696 537266 267708
rect 539042 267696 539048 267708
rect 537260 267668 539048 267696
rect 537260 267656 537266 267668
rect 539042 267656 539048 267668
rect 539100 267656 539106 267708
rect 539686 267656 539692 267708
rect 539744 267696 539750 267708
rect 543550 267696 543556 267708
rect 539744 267668 543556 267696
rect 539744 267656 539750 267668
rect 543550 267656 543556 267668
rect 543608 267656 543614 267708
rect 543688 267656 543694 267708
rect 543746 267696 543752 267708
rect 546402 267696 546408 267708
rect 543746 267668 546408 267696
rect 543746 267656 543752 267668
rect 546402 267656 546408 267668
rect 546460 267656 546466 267708
rect 546586 267656 546592 267708
rect 546644 267696 546650 267708
rect 580258 267696 580264 267708
rect 546644 267668 580264 267696
rect 546644 267656 546650 267668
rect 580258 267656 580264 267668
rect 580316 267656 580322 267708
rect 88978 267520 88984 267572
rect 89036 267560 89042 267572
rect 144546 267560 144552 267572
rect 89036 267532 144552 267560
rect 89036 267520 89042 267532
rect 144546 267520 144552 267532
rect 144604 267520 144610 267572
rect 144914 267520 144920 267572
rect 144972 267560 144978 267572
rect 150526 267560 150532 267572
rect 144972 267532 150532 267560
rect 144972 267520 144978 267532
rect 150526 267520 150532 267532
rect 150584 267520 150590 267572
rect 151078 267520 151084 267572
rect 151136 267560 151142 267572
rect 172882 267560 172888 267572
rect 151136 267532 172888 267560
rect 151136 267520 151142 267532
rect 172882 267520 172888 267532
rect 172940 267520 172946 267572
rect 187142 267520 187148 267572
rect 187200 267560 187206 267572
rect 221734 267560 221740 267572
rect 187200 267532 221740 267560
rect 187200 267520 187206 267532
rect 221734 267520 221740 267532
rect 221792 267520 221798 267572
rect 227714 267520 227720 267572
rect 227772 267560 227778 267572
rect 234154 267560 234160 267572
rect 227772 267532 234160 267560
rect 227772 267520 227778 267532
rect 234154 267520 234160 267532
rect 234212 267520 234218 267572
rect 313642 267520 313648 267572
rect 313700 267560 313706 267572
rect 317782 267560 317788 267572
rect 313700 267532 317788 267560
rect 313700 267520 313706 267532
rect 317782 267520 317788 267532
rect 317840 267520 317846 267572
rect 370774 267520 370780 267572
rect 370832 267560 370838 267572
rect 381538 267560 381544 267572
rect 370832 267532 381544 267560
rect 370832 267520 370838 267532
rect 381538 267520 381544 267532
rect 381596 267520 381602 267572
rect 383194 267520 383200 267572
rect 383252 267560 383258 267572
rect 394694 267560 394700 267572
rect 383252 267532 394700 267560
rect 383252 267520 383258 267532
rect 394694 267520 394700 267532
rect 394752 267520 394758 267572
rect 397086 267520 397092 267572
rect 397144 267560 397150 267572
rect 422294 267560 422300 267572
rect 397144 267532 422300 267560
rect 397144 267520 397150 267532
rect 422294 267520 422300 267532
rect 422352 267520 422358 267572
rect 443454 267520 443460 267572
rect 443512 267560 443518 267572
rect 449894 267560 449900 267572
rect 443512 267532 449900 267560
rect 443512 267520 443518 267532
rect 449894 267520 449900 267532
rect 449952 267520 449958 267572
rect 450078 267520 450084 267572
rect 450136 267560 450142 267572
rect 481542 267560 481548 267572
rect 450136 267532 481548 267560
rect 450136 267520 450142 267532
rect 481542 267520 481548 267532
rect 481600 267520 481606 267572
rect 481726 267520 481732 267572
rect 481784 267560 481790 267572
rect 503070 267560 503076 267572
rect 481784 267532 503076 267560
rect 481784 267520 481790 267532
rect 503070 267520 503076 267532
rect 503128 267520 503134 267572
rect 504174 267520 504180 267572
rect 504232 267560 504238 267572
rect 504232 267532 504588 267560
rect 504232 267520 504238 267532
rect 107562 267384 107568 267436
rect 107620 267424 107626 267436
rect 167086 267424 167092 267436
rect 107620 267396 167092 267424
rect 107620 267384 107626 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 167730 267384 167736 267436
rect 167788 267424 167794 267436
rect 204346 267424 204352 267436
rect 167788 267396 204352 267424
rect 167788 267384 167794 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 211982 267384 211988 267436
rect 212040 267424 212046 267436
rect 222562 267424 222568 267436
rect 212040 267396 222568 267424
rect 212040 267384 212046 267396
rect 222562 267384 222568 267396
rect 222620 267384 222626 267436
rect 224218 267384 224224 267436
rect 224276 267424 224282 267436
rect 231670 267424 231676 267436
rect 224276 267396 231676 267424
rect 224276 267384 224282 267396
rect 231670 267384 231676 267396
rect 231728 267384 231734 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 246574 267424 246580 267436
rect 233936 267396 246580 267424
rect 233936 267384 233942 267396
rect 246574 267384 246580 267396
rect 246632 267384 246638 267436
rect 334342 267384 334348 267436
rect 334400 267424 334406 267436
rect 342898 267424 342904 267436
rect 334400 267396 342904 267424
rect 334400 267384 334406 267396
rect 342898 267384 342904 267396
rect 342956 267384 342962 267436
rect 350902 267384 350908 267436
rect 350960 267424 350966 267436
rect 361022 267424 361028 267436
rect 350960 267396 361028 267424
rect 350960 267384 350966 267396
rect 361022 267384 361028 267396
rect 361080 267384 361086 267436
rect 365806 267384 365812 267436
rect 365864 267424 365870 267436
rect 382918 267424 382924 267436
rect 365864 267396 382924 267424
rect 365864 267384 365870 267396
rect 382918 267384 382924 267396
rect 382976 267384 382982 267436
rect 390646 267384 390652 267436
rect 390704 267424 390710 267436
rect 404354 267424 404360 267436
rect 390704 267396 404360 267424
rect 390704 267384 390710 267396
rect 404354 267384 404360 267396
rect 404412 267384 404418 267436
rect 409598 267384 409604 267436
rect 409656 267424 409662 267436
rect 435358 267424 435364 267436
rect 409656 267396 435364 267424
rect 409656 267384 409662 267396
rect 435358 267384 435364 267396
rect 435416 267384 435422 267436
rect 440326 267384 440332 267436
rect 440384 267424 440390 267436
rect 485728 267424 485734 267436
rect 440384 267396 485734 267424
rect 440384 267384 440390 267396
rect 485728 267384 485734 267396
rect 485786 267384 485792 267436
rect 485866 267384 485872 267436
rect 485924 267424 485930 267436
rect 487062 267424 487068 267436
rect 485924 267396 487068 267424
rect 485924 267384 485930 267396
rect 487062 267384 487068 267396
rect 487120 267384 487126 267436
rect 487246 267384 487252 267436
rect 487304 267424 487310 267436
rect 491478 267424 491484 267436
rect 487304 267396 491484 267424
rect 487304 267384 487310 267396
rect 491478 267384 491484 267396
rect 491536 267384 491542 267436
rect 491662 267384 491668 267436
rect 491720 267424 491726 267436
rect 492490 267424 492496 267436
rect 491720 267396 492496 267424
rect 491720 267384 491726 267396
rect 492490 267384 492496 267396
rect 492548 267384 492554 267436
rect 492674 267384 492680 267436
rect 492732 267424 492738 267436
rect 504358 267424 504364 267436
rect 492732 267396 504364 267424
rect 492732 267384 492738 267396
rect 504358 267384 504364 267396
rect 504416 267384 504422 267436
rect 504560 267424 504588 267532
rect 506474 267520 506480 267572
rect 506532 267560 506538 267572
rect 507210 267560 507216 267572
rect 506532 267532 507216 267560
rect 506532 267520 506538 267532
rect 507210 267520 507216 267532
rect 507268 267520 507274 267572
rect 507394 267520 507400 267572
rect 507452 267560 507458 267572
rect 578878 267560 578884 267572
rect 507452 267532 578884 267560
rect 507452 267520 507458 267532
rect 578878 267520 578884 267532
rect 578936 267520 578942 267572
rect 552842 267424 552848 267436
rect 504560 267396 552848 267424
rect 552842 267384 552848 267396
rect 552900 267384 552906 267436
rect 100662 267248 100668 267300
rect 100720 267288 100726 267300
rect 159818 267288 159824 267300
rect 100720 267260 159824 267288
rect 100720 267248 100726 267260
rect 159818 267248 159824 267260
rect 159876 267248 159882 267300
rect 166902 267248 166908 267300
rect 166960 267288 166966 267300
rect 174538 267288 174544 267300
rect 166960 267260 174544 267288
rect 166960 267248 166966 267260
rect 174538 267248 174544 267260
rect 174596 267248 174602 267300
rect 175090 267248 175096 267300
rect 175148 267288 175154 267300
rect 214282 267288 214288 267300
rect 175148 267260 214288 267288
rect 175148 267248 175154 267260
rect 214282 267248 214288 267260
rect 214340 267248 214346 267300
rect 220078 267248 220084 267300
rect 220136 267288 220142 267300
rect 239122 267288 239128 267300
rect 220136 267260 239128 267288
rect 220136 267248 220142 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 254578 267248 254584 267300
rect 254636 267288 254642 267300
rect 262306 267288 262312 267300
rect 254636 267260 262312 267288
rect 254636 267248 254642 267260
rect 262306 267248 262312 267260
rect 262364 267248 262370 267300
rect 312814 267248 312820 267300
rect 312872 267288 312878 267300
rect 316034 267288 316040 267300
rect 312872 267260 316040 267288
rect 312872 267248 312878 267260
rect 316034 267248 316040 267260
rect 316092 267248 316098 267300
rect 343450 267248 343456 267300
rect 343508 267288 343514 267300
rect 353938 267288 353944 267300
rect 343508 267260 353944 267288
rect 343508 267248 343514 267260
rect 353938 267248 353944 267260
rect 353996 267248 354002 267300
rect 363322 267248 363328 267300
rect 363380 267288 363386 267300
rect 370498 267288 370504 267300
rect 363380 267260 370504 267288
rect 363380 267248 363386 267260
rect 370498 267248 370504 267260
rect 370556 267248 370562 267300
rect 375742 267248 375748 267300
rect 375800 267288 375806 267300
rect 393958 267288 393964 267300
rect 375800 267260 393964 267288
rect 375800 267248 375806 267260
rect 393958 267248 393964 267260
rect 394016 267248 394022 267300
rect 399754 267248 399760 267300
rect 399812 267288 399818 267300
rect 418982 267288 418988 267300
rect 399812 267260 418988 267288
rect 399812 267248 399818 267260
rect 418982 267248 418988 267260
rect 419040 267248 419046 267300
rect 421282 267248 421288 267300
rect 421340 267288 421346 267300
rect 464338 267288 464344 267300
rect 421340 267260 464344 267288
rect 421340 267248 421346 267260
rect 464338 267248 464344 267260
rect 464396 267248 464402 267300
rect 465166 267248 465172 267300
rect 465224 267288 465230 267300
rect 480898 267288 480904 267300
rect 465224 267260 480904 267288
rect 465224 267248 465230 267260
rect 480898 267248 480904 267260
rect 480956 267248 480962 267300
rect 481082 267248 481088 267300
rect 481140 267288 481146 267300
rect 518802 267288 518808 267300
rect 481140 267260 518808 267288
rect 481140 267248 481146 267260
rect 518802 267248 518808 267260
rect 518860 267248 518866 267300
rect 518986 267248 518992 267300
rect 519044 267288 519050 267300
rect 533890 267288 533896 267300
rect 519044 267260 533896 267288
rect 519044 267248 519050 267260
rect 533890 267248 533896 267260
rect 533948 267248 533954 267300
rect 534028 267248 534034 267300
rect 534086 267288 534092 267300
rect 538858 267288 538864 267300
rect 534086 267260 538864 267288
rect 534086 267248 534092 267260
rect 538858 267248 538864 267260
rect 538916 267248 538922 267300
rect 539042 267248 539048 267300
rect 539100 267288 539106 267300
rect 621658 267288 621664 267300
rect 539100 267260 621664 267288
rect 539100 267248 539106 267260
rect 621658 267248 621664 267260
rect 621716 267248 621722 267300
rect 71038 267112 71044 267164
rect 71096 267152 71102 267164
rect 138106 267152 138112 267164
rect 71096 267124 138112 267152
rect 71096 267112 71102 267124
rect 138106 267112 138112 267124
rect 138164 267112 138170 267164
rect 141418 267112 141424 267164
rect 141476 267152 141482 267164
rect 141476 267124 142154 267152
rect 141476 267112 141482 267124
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 141418 267016 141424 267028
rect 73856 266988 141424 267016
rect 73856 266976 73862 266988
rect 141418 266976 141424 266988
rect 141476 266976 141482 267028
rect 142126 267016 142154 267124
rect 144546 267112 144552 267164
rect 144604 267152 144610 267164
rect 147398 267152 147404 267164
rect 144604 267124 147404 267152
rect 144604 267112 144610 267124
rect 147398 267112 147404 267124
rect 147456 267112 147462 267164
rect 147582 267112 147588 267164
rect 147640 267152 147646 267164
rect 149054 267152 149060 267164
rect 147640 267124 149060 267152
rect 147640 267112 147646 267124
rect 149054 267112 149060 267124
rect 149112 267112 149118 267164
rect 149882 267112 149888 267164
rect 149940 267152 149946 267164
rect 194410 267152 194416 267164
rect 149940 267124 194416 267152
rect 149940 267112 149946 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 199654 267112 199660 267164
rect 199712 267152 199718 267164
rect 218422 267152 218428 267164
rect 199712 267124 218428 267152
rect 199712 267112 199718 267124
rect 218422 267112 218428 267124
rect 218480 267112 218486 267164
rect 221458 267112 221464 267164
rect 221516 267152 221522 267164
rect 241606 267152 241612 267164
rect 221516 267124 241612 267152
rect 221516 267112 221522 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 335998 267112 336004 267164
rect 336056 267152 336062 267164
rect 347038 267152 347044 267164
rect 336056 267124 347044 267152
rect 336056 267112 336062 267124
rect 347038 267112 347044 267124
rect 347096 267112 347102 267164
rect 355870 267112 355876 267164
rect 355928 267152 355934 267164
rect 369118 267152 369124 267164
rect 355928 267124 369124 267152
rect 355928 267112 355934 267124
rect 369118 267112 369124 267124
rect 369176 267112 369182 267164
rect 373258 267112 373264 267164
rect 373316 267152 373322 267164
rect 392578 267152 392584 267164
rect 373316 267124 392584 267152
rect 373316 267112 373322 267124
rect 392578 267112 392584 267124
rect 392636 267112 392642 267164
rect 404722 267112 404728 267164
rect 404780 267152 404786 267164
rect 431954 267152 431960 267164
rect 404780 267124 431960 267152
rect 404780 267112 404786 267124
rect 431954 267112 431960 267124
rect 432012 267112 432018 267164
rect 439498 267112 439504 267164
rect 439556 267152 439562 267164
rect 445018 267152 445024 267164
rect 439556 267124 445024 267152
rect 439556 267112 439562 267124
rect 445018 267112 445024 267124
rect 445076 267112 445082 267164
rect 445294 267112 445300 267164
rect 445352 267152 445358 267164
rect 450078 267152 450084 267164
rect 445352 267124 450084 267152
rect 445352 267112 445358 267124
rect 450078 267112 450084 267124
rect 450136 267112 450142 267164
rect 450262 267112 450268 267164
rect 450320 267152 450326 267164
rect 499574 267152 499580 267164
rect 450320 267124 499580 267152
rect 450320 267112 450326 267124
rect 499574 267112 499580 267124
rect 499632 267112 499638 267164
rect 499758 267112 499764 267164
rect 499816 267152 499822 267164
rect 504174 267152 504180 267164
rect 499816 267124 504180 267152
rect 499816 267112 499822 267124
rect 504174 267112 504180 267124
rect 504232 267112 504238 267164
rect 504358 267112 504364 267164
rect 504416 267152 504422 267164
rect 521746 267152 521752 267164
rect 504416 267124 521752 267152
rect 504416 267112 504422 267124
rect 521746 267112 521752 267124
rect 521804 267112 521810 267164
rect 585778 267152 585784 267164
rect 522960 267124 585784 267152
rect 184014 267016 184020 267028
rect 142126 266988 184020 267016
rect 184014 266976 184020 266988
rect 184072 266976 184078 267028
rect 184198 266976 184204 267028
rect 184256 267016 184262 267028
rect 184256 266988 190454 267016
rect 184256 266976 184262 266988
rect 132402 266840 132408 266892
rect 132460 266880 132466 266892
rect 184474 266880 184480 266892
rect 132460 266852 184480 266880
rect 132460 266840 132466 266852
rect 184474 266840 184480 266852
rect 184532 266840 184538 266892
rect 190426 266880 190454 266988
rect 193858 266976 193864 267028
rect 193916 267016 193922 267028
rect 201862 267016 201868 267028
rect 193916 266988 201868 267016
rect 193916 266976 193922 266988
rect 201862 266976 201868 266988
rect 201920 266976 201926 267028
rect 206278 266976 206284 267028
rect 206336 267016 206342 267028
rect 228358 267016 228364 267028
rect 206336 266988 228364 267016
rect 206336 266976 206342 266988
rect 228358 266976 228364 266988
rect 228416 266976 228422 267028
rect 237282 266976 237288 267028
rect 237340 267016 237346 267028
rect 254026 267016 254032 267028
rect 237340 266988 254032 267016
rect 237340 266976 237346 266988
rect 254026 266976 254032 266988
rect 254084 266976 254090 267028
rect 271414 267016 271420 267028
rect 258046 266988 271420 267016
rect 258046 266892 258074 266988
rect 271414 266976 271420 266988
rect 271472 266976 271478 267028
rect 276658 266976 276664 267028
rect 276716 267016 276722 267028
rect 278038 267016 278044 267028
rect 276716 266988 278044 267016
rect 276716 266976 276722 266988
rect 278038 266976 278044 266988
rect 278096 266976 278102 267028
rect 286962 266976 286968 267028
rect 287020 267016 287026 267028
rect 291286 267016 291292 267028
rect 287020 266988 291292 267016
rect 287020 266976 287026 266988
rect 291286 266976 291292 266988
rect 291344 266976 291350 267028
rect 295150 266976 295156 267028
rect 295208 267016 295214 267028
rect 297082 267016 297088 267028
rect 295208 266988 297088 267016
rect 295208 266976 295214 266988
rect 297082 266976 297088 266988
rect 297140 266976 297146 267028
rect 316126 266976 316132 267028
rect 316184 267016 316190 267028
rect 320174 267016 320180 267028
rect 316184 266988 320180 267016
rect 316184 266976 316190 266988
rect 320174 266976 320180 266988
rect 320232 266976 320238 267028
rect 324406 266976 324412 267028
rect 324464 267016 324470 267028
rect 332502 267016 332508 267028
rect 324464 266988 332508 267016
rect 324464 266976 324470 266988
rect 332502 266976 332508 266988
rect 332560 266976 332566 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 355318 267016 355324 267028
rect 353444 266988 355324 267016
rect 353444 266976 353450 266988
rect 355318 266976 355324 266988
rect 355376 266976 355382 267028
rect 378226 266976 378232 267028
rect 378284 267016 378290 267028
rect 409138 267016 409144 267028
rect 378284 266988 409144 267016
rect 378284 266976 378290 266988
rect 409138 266976 409144 266988
rect 409196 266976 409202 267028
rect 422110 266976 422116 267028
rect 422168 267016 422174 267028
rect 443454 267016 443460 267028
rect 422168 266988 443460 267016
rect 422168 266976 422174 266988
rect 443454 266976 443460 266988
rect 443512 266976 443518 267028
rect 451918 267016 451924 267028
rect 443748 266988 451924 267016
rect 209314 266880 209320 266892
rect 190426 266852 209320 266880
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 257982 266840 257988 266892
rect 258040 266852 258074 266892
rect 258040 266840 258046 266852
rect 320266 266840 320272 266892
rect 320324 266880 320330 266892
rect 327442 266880 327448 266892
rect 320324 266852 327448 266880
rect 320324 266840 320330 266852
rect 327442 266840 327448 266852
rect 327500 266840 327506 266892
rect 342622 266840 342628 266892
rect 342680 266880 342686 266892
rect 356514 266880 356520 266892
rect 342680 266852 356520 266880
rect 342680 266840 342686 266852
rect 356514 266840 356520 266852
rect 356572 266840 356578 266892
rect 359182 266840 359188 266892
rect 359240 266880 359246 266892
rect 359240 266852 364334 266880
rect 359240 266840 359246 266852
rect 265066 266772 265072 266824
rect 265124 266812 265130 266824
rect 268930 266812 268936 266824
rect 265124 266784 268936 266812
rect 265124 266772 265130 266784
rect 268930 266772 268936 266784
rect 268988 266772 268994 266824
rect 331858 266772 331864 266824
rect 331916 266812 331922 266824
rect 335630 266812 335636 266824
rect 331916 266784 335636 266812
rect 331916 266772 331922 266784
rect 335630 266772 335636 266784
rect 335688 266772 335694 266824
rect 120718 266704 120724 266756
rect 120776 266744 120782 266756
rect 157150 266744 157156 266756
rect 120776 266716 157156 266744
rect 120776 266704 120782 266716
rect 157150 266704 157156 266716
rect 157208 266704 157214 266756
rect 169018 266704 169024 266756
rect 169076 266744 169082 266756
rect 172054 266744 172060 266756
rect 169076 266716 172060 266744
rect 169076 266704 169082 266716
rect 172054 266704 172060 266716
rect 172112 266704 172118 266756
rect 184014 266704 184020 266756
rect 184072 266744 184078 266756
rect 189442 266744 189448 266756
rect 184072 266716 189448 266744
rect 184072 266704 184078 266716
rect 189442 266704 189448 266716
rect 189500 266704 189506 266756
rect 240686 266704 240692 266756
rect 240744 266744 240750 266756
rect 245746 266744 245752 266756
rect 240744 266716 245752 266744
rect 240744 266704 240750 266716
rect 245746 266704 245752 266716
rect 245804 266704 245810 266756
rect 249058 266704 249064 266756
rect 249116 266744 249122 266756
rect 251542 266744 251548 266756
rect 249116 266716 251548 266744
rect 249116 266704 249122 266716
rect 251542 266704 251548 266716
rect 251600 266704 251606 266756
rect 358354 266704 358360 266756
rect 358412 266744 358418 266756
rect 360838 266744 360844 266756
rect 358412 266716 360844 266744
rect 358412 266704 358418 266716
rect 360838 266704 360844 266716
rect 360896 266704 360902 266756
rect 330202 266636 330208 266688
rect 330260 266676 330266 266688
rect 334618 266676 334624 266688
rect 330260 266648 334624 266676
rect 330260 266636 330266 266648
rect 334618 266636 334624 266648
rect 334676 266636 334682 266688
rect 364306 266676 364334 266852
rect 393130 266840 393136 266892
rect 393188 266880 393194 266892
rect 401594 266880 401600 266892
rect 393188 266852 401600 266880
rect 393188 266840 393194 266852
rect 401594 266840 401600 266852
rect 401652 266840 401658 266892
rect 405550 266840 405556 266892
rect 405608 266880 405614 266892
rect 425698 266880 425704 266892
rect 405608 266852 425704 266880
rect 405608 266840 405614 266852
rect 425698 266840 425704 266852
rect 425756 266840 425762 266892
rect 428458 266880 428464 266892
rect 425900 266852 428464 266880
rect 412174 266704 412180 266756
rect 412232 266744 412238 266756
rect 412232 266716 412634 266744
rect 412232 266704 412238 266716
rect 373074 266676 373080 266688
rect 364306 266648 373080 266676
rect 373074 266636 373080 266648
rect 373132 266636 373138 266688
rect 138658 266568 138664 266620
rect 138716 266608 138722 266620
rect 138716 266580 145328 266608
rect 138716 266568 138722 266580
rect 119798 266432 119804 266484
rect 119856 266472 119862 266484
rect 144914 266472 144920 266484
rect 119856 266444 144920 266472
rect 119856 266432 119862 266444
rect 144914 266432 144920 266444
rect 144972 266432 144978 266484
rect 145300 266404 145328 266580
rect 149054 266568 149060 266620
rect 149112 266608 149118 266620
rect 179506 266608 179512 266620
rect 149112 266580 179512 266608
rect 149112 266568 149118 266580
rect 179506 266568 179512 266580
rect 179564 266568 179570 266620
rect 213822 266568 213828 266620
rect 213880 266608 213886 266620
rect 220078 266608 220084 266620
rect 213880 266580 220084 266608
rect 213880 266568 213886 266580
rect 220078 266568 220084 266580
rect 220136 266568 220142 266620
rect 245102 266568 245108 266620
rect 245160 266608 245166 266620
rect 249058 266608 249064 266620
rect 245160 266580 249064 266608
rect 245160 266568 245166 266580
rect 249058 266568 249064 266580
rect 249116 266568 249122 266620
rect 360838 266568 360844 266620
rect 360896 266608 360902 266620
rect 362218 266608 362224 266620
rect 360896 266580 362224 266608
rect 360896 266568 360902 266580
rect 362218 266568 362224 266580
rect 362276 266568 362282 266620
rect 412606 266608 412634 266716
rect 417970 266704 417976 266756
rect 418028 266744 418034 266756
rect 425900 266744 425928 266852
rect 428458 266840 428464 266852
rect 428516 266840 428522 266892
rect 435174 266840 435180 266892
rect 435232 266880 435238 266892
rect 439314 266880 439320 266892
rect 435232 266852 439320 266880
rect 435232 266840 435238 266852
rect 439314 266840 439320 266852
rect 439372 266840 439378 266892
rect 418028 266716 425928 266744
rect 418028 266704 418034 266716
rect 427906 266704 427912 266756
rect 427964 266744 427970 266756
rect 443748 266744 443776 266988
rect 451918 266976 451924 266988
rect 451976 266976 451982 267028
rect 455230 266976 455236 267028
rect 455288 267016 455294 267028
rect 460198 267016 460204 267028
rect 455288 266988 460204 267016
rect 455288 266976 455294 266988
rect 460198 266976 460204 266988
rect 460256 266976 460262 267028
rect 462314 266976 462320 267028
rect 462372 267016 462378 267028
rect 464982 267016 464988 267028
rect 462372 266988 464988 267016
rect 462372 266976 462378 266988
rect 464982 266976 464988 266988
rect 465040 266976 465046 267028
rect 465534 266976 465540 267028
rect 465592 267016 465598 267028
rect 512914 267016 512920 267028
rect 465592 266988 512920 267016
rect 465592 266976 465598 266988
rect 512914 266976 512920 266988
rect 512972 266976 512978 267028
rect 513374 266976 513380 267028
rect 513432 267016 513438 267028
rect 518802 267016 518808 267028
rect 513432 266988 518808 267016
rect 513432 266976 513438 266988
rect 518802 266976 518808 266988
rect 518860 266976 518866 267028
rect 518986 266976 518992 267028
rect 519044 267016 519050 267028
rect 520090 267016 520096 267028
rect 519044 266988 520096 267016
rect 519044 266976 519050 266988
rect 520090 266976 520096 266988
rect 520148 266976 520154 267028
rect 520274 266976 520280 267028
rect 520332 267016 520338 267028
rect 522960 267016 522988 267124
rect 585778 267112 585784 267124
rect 585836 267112 585842 267164
rect 520332 266988 522988 267016
rect 520332 266976 520338 266988
rect 523126 266976 523132 267028
rect 523184 267016 523190 267028
rect 524322 267016 524328 267028
rect 523184 266988 524328 267016
rect 523184 266976 523190 266988
rect 524322 266976 524328 266988
rect 524380 266976 524386 267028
rect 524782 266976 524788 267028
rect 524840 267016 524846 267028
rect 525702 267016 525708 267028
rect 524840 266988 525708 267016
rect 524840 266976 524846 266988
rect 525702 266976 525708 266988
rect 525760 266976 525766 267028
rect 525886 266976 525892 267028
rect 525944 267016 525950 267028
rect 613378 267016 613384 267028
rect 525944 266988 613384 267016
rect 525944 266976 525950 266988
rect 613378 266976 613384 266988
rect 613436 266976 613442 267028
rect 622394 267016 622400 267028
rect 615466 266988 622400 267016
rect 471238 266880 471244 266892
rect 427964 266716 443776 266744
rect 443840 266852 471244 266880
rect 427964 266704 427970 266716
rect 421558 266608 421564 266620
rect 412606 266580 421564 266608
rect 421558 266568 421564 266580
rect 421616 266568 421622 266620
rect 422938 266568 422944 266620
rect 422996 266608 423002 266620
rect 435174 266608 435180 266620
rect 422996 266580 435180 266608
rect 422996 266568 423002 266580
rect 435174 266568 435180 266580
rect 435232 266568 435238 266620
rect 435358 266568 435364 266620
rect 435416 266608 435422 266620
rect 443840 266608 443868 266852
rect 471238 266840 471244 266852
rect 471296 266840 471302 266892
rect 471624 266852 475608 266880
rect 449434 266704 449440 266756
rect 449492 266744 449498 266756
rect 449492 266716 451274 266744
rect 449492 266704 449498 266716
rect 435416 266580 443868 266608
rect 435416 266568 435422 266580
rect 145558 266500 145564 266552
rect 145616 266540 145622 266552
rect 148870 266540 148876 266552
rect 145616 266512 148876 266540
rect 145616 266500 145622 266512
rect 148870 266500 148876 266512
rect 148928 266500 148934 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 331674 266540 331680 266552
rect 327776 266512 331680 266540
rect 327776 266500 327782 266512
rect 331674 266500 331680 266512
rect 331732 266500 331738 266552
rect 346762 266500 346768 266552
rect 346820 266540 346826 266552
rect 351638 266540 351644 266552
rect 346820 266512 351644 266540
rect 346820 266500 346826 266512
rect 351638 266500 351644 266512
rect 351696 266500 351702 266552
rect 355042 266500 355048 266552
rect 355100 266540 355106 266552
rect 359734 266540 359740 266552
rect 355100 266512 359740 266540
rect 355100 266500 355106 266512
rect 359734 266500 359740 266512
rect 359792 266500 359798 266552
rect 394786 266500 394792 266552
rect 394844 266540 394850 266552
rect 397914 266540 397920 266552
rect 394844 266512 397920 266540
rect 394844 266500 394850 266512
rect 397914 266500 397920 266512
rect 397972 266500 397978 266552
rect 444466 266500 444472 266552
rect 444524 266540 444530 266552
rect 447778 266540 447784 266552
rect 444524 266512 447784 266540
rect 444524 266500 444530 266512
rect 447778 266500 447784 266512
rect 447836 266500 447842 266552
rect 451246 266540 451274 266716
rect 456426 266704 456432 266756
rect 456484 266744 456490 266756
rect 462314 266744 462320 266756
rect 456484 266716 462320 266744
rect 456484 266704 456490 266716
rect 462314 266704 462320 266716
rect 462372 266704 462378 266756
rect 464522 266744 464528 266756
rect 462516 266716 464528 266744
rect 452746 266636 452752 266688
rect 452804 266676 452810 266688
rect 456150 266676 456156 266688
rect 452804 266648 456156 266676
rect 452804 266636 452810 266648
rect 456150 266636 456156 266648
rect 456208 266636 456214 266688
rect 459186 266568 459192 266620
rect 459244 266608 459250 266620
rect 462516 266608 462544 266716
rect 464522 266704 464528 266716
rect 464580 266704 464586 266756
rect 464982 266704 464988 266756
rect 465040 266744 465046 266756
rect 469214 266744 469220 266756
rect 465040 266716 469220 266744
rect 465040 266704 465046 266716
rect 469214 266704 469220 266716
rect 469272 266704 469278 266756
rect 459244 266580 462544 266608
rect 459244 266568 459250 266580
rect 462682 266568 462688 266620
rect 462740 266608 462746 266620
rect 463510 266608 463516 266620
rect 462740 266580 463516 266608
rect 462740 266568 462746 266580
rect 463510 266568 463516 266580
rect 463568 266568 463574 266620
rect 464338 266568 464344 266620
rect 464396 266608 464402 266620
rect 465718 266608 465724 266620
rect 464396 266580 465724 266608
rect 464396 266568 464402 266580
rect 465718 266568 465724 266580
rect 465776 266568 465782 266620
rect 469306 266568 469312 266620
rect 469364 266608 469370 266620
rect 471624 266608 471652 266852
rect 471790 266704 471796 266756
rect 471848 266744 471854 266756
rect 475378 266744 475384 266756
rect 471848 266716 475384 266744
rect 471848 266704 471854 266716
rect 475378 266704 475384 266716
rect 475436 266704 475442 266756
rect 469364 266580 471652 266608
rect 469364 266568 469370 266580
rect 473446 266568 473452 266620
rect 473504 266608 473510 266620
rect 474642 266608 474648 266620
rect 473504 266580 474648 266608
rect 473504 266568 473510 266580
rect 474642 266568 474648 266580
rect 474700 266568 474706 266620
rect 475580 266608 475608 266852
rect 480898 266840 480904 266892
rect 480956 266880 480962 266892
rect 492674 266880 492680 266892
rect 480956 266852 492680 266880
rect 480956 266840 480962 266852
rect 492674 266840 492680 266852
rect 492732 266840 492738 266892
rect 497458 266840 497464 266892
rect 497516 266880 497522 266892
rect 499758 266880 499764 266892
rect 497516 266852 499764 266880
rect 497516 266840 497522 266852
rect 499758 266840 499764 266852
rect 499816 266840 499822 266892
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 500862 266880 500868 266892
rect 500000 266852 500868 266880
rect 500000 266840 500006 266852
rect 500862 266840 500868 266852
rect 500920 266840 500926 266892
rect 501046 266840 501052 266892
rect 501104 266880 501110 266892
rect 506382 266880 506388 266892
rect 501104 266852 506388 266880
rect 501104 266840 501110 266852
rect 506382 266840 506388 266852
rect 506440 266840 506446 266892
rect 506566 266840 506572 266892
rect 506624 266880 506630 266892
rect 507670 266880 507676 266892
rect 506624 266852 507676 266880
rect 506624 266840 506630 266852
rect 507670 266840 507676 266852
rect 507728 266840 507734 266892
rect 507854 266840 507860 266892
rect 507912 266880 507918 266892
rect 570598 266880 570604 266892
rect 507912 266852 570604 266880
rect 507912 266840 507918 266852
rect 570598 266840 570604 266852
rect 570656 266840 570662 266892
rect 615466 266880 615494 266988
rect 622394 266976 622400 266988
rect 622452 266976 622458 267028
rect 576826 266852 615494 266880
rect 475930 266704 475936 266756
rect 475988 266744 475994 266756
rect 481082 266744 481088 266756
rect 475988 266716 481088 266744
rect 475988 266704 475994 266716
rect 481082 266704 481088 266716
rect 481140 266704 481146 266756
rect 481542 266704 481548 266756
rect 481600 266744 481606 266756
rect 492306 266744 492312 266756
rect 481600 266716 492312 266744
rect 481600 266704 481606 266716
rect 492306 266704 492312 266716
rect 492364 266704 492370 266756
rect 492490 266704 492496 266756
rect 492548 266744 492554 266756
rect 492548 266716 552704 266744
rect 492548 266704 492554 266716
rect 477310 266608 477316 266620
rect 475580 266580 477316 266608
rect 477310 266568 477316 266580
rect 477368 266568 477374 266620
rect 477586 266568 477592 266620
rect 477644 266608 477650 266620
rect 485682 266608 485688 266620
rect 477644 266580 485688 266608
rect 477644 266568 477650 266580
rect 485682 266568 485688 266580
rect 485740 266568 485746 266620
rect 486050 266568 486056 266620
rect 486108 266608 486114 266620
rect 488718 266608 488724 266620
rect 486108 266580 488724 266608
rect 486108 266568 486114 266580
rect 488718 266568 488724 266580
rect 488776 266568 488782 266620
rect 490006 266568 490012 266620
rect 490064 266608 490070 266620
rect 534074 266608 534080 266620
rect 490064 266580 534080 266608
rect 490064 266568 490070 266580
rect 534074 266568 534080 266580
rect 534132 266568 534138 266620
rect 538674 266608 538680 266620
rect 534276 266580 538680 266608
rect 453298 266540 453304 266552
rect 451246 266512 453304 266540
rect 453298 266500 453304 266512
rect 453356 266500 453362 266552
rect 454402 266500 454408 266552
rect 454460 266540 454466 266552
rect 457438 266540 457444 266552
rect 454460 266512 457444 266540
rect 454460 266500 454466 266512
rect 457438 266500 457444 266512
rect 457496 266500 457502 266552
rect 159818 266432 159824 266484
rect 159876 266472 159882 266484
rect 162118 266472 162124 266484
rect 159876 266444 162124 266472
rect 159876 266432 159882 266444
rect 162118 266432 162124 266444
rect 162176 266432 162182 266484
rect 208670 266432 208676 266484
rect 208728 266472 208734 266484
rect 210970 266472 210976 266484
rect 208728 266444 210976 266472
rect 208728 266432 208734 266444
rect 210970 266432 210976 266444
rect 211028 266432 211034 266484
rect 361666 266432 361672 266484
rect 361724 266472 361730 266484
rect 362770 266472 362776 266484
rect 361724 266444 362776 266472
rect 361724 266432 361730 266444
rect 362770 266432 362776 266444
rect 362828 266432 362834 266484
rect 460198 266432 460204 266484
rect 460256 266472 460262 266484
rect 460256 266444 512224 266472
rect 460256 266432 460262 266444
rect 147214 266404 147220 266416
rect 145300 266376 147220 266404
rect 147214 266364 147220 266376
rect 147272 266364 147278 266416
rect 148318 266364 148324 266416
rect 148376 266404 148382 266416
rect 149698 266404 149704 266416
rect 148376 266376 149704 266404
rect 148376 266364 148382 266376
rect 149698 266364 149704 266376
rect 149756 266364 149762 266416
rect 156598 266364 156604 266416
rect 156656 266404 156662 266416
rect 159634 266404 159640 266416
rect 156656 266376 159640 266404
rect 156656 266364 156662 266376
rect 159634 266364 159640 266376
rect 159692 266364 159698 266416
rect 182174 266364 182180 266416
rect 182232 266404 182238 266416
rect 186130 266404 186136 266416
rect 182232 266376 186136 266404
rect 182232 266364 182238 266376
rect 186130 266364 186136 266376
rect 186188 266364 186194 266416
rect 202138 266364 202144 266416
rect 202196 266404 202202 266416
rect 206830 266404 206836 266416
rect 202196 266376 206836 266404
rect 202196 266364 202202 266376
rect 206830 266364 206836 266376
rect 206888 266364 206894 266416
rect 222838 266364 222844 266416
rect 222896 266404 222902 266416
rect 224218 266404 224224 266416
rect 222896 266376 224224 266404
rect 222896 266364 222902 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 230750 266364 230756 266416
rect 230808 266404 230814 266416
rect 236638 266404 236644 266416
rect 230808 266376 236644 266404
rect 230808 266364 230814 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 242250 266364 242256 266416
rect 242308 266404 242314 266416
rect 243262 266404 243268 266416
rect 242308 266376 243268 266404
rect 242308 266364 242314 266376
rect 243262 266364 243268 266376
rect 243320 266364 243326 266416
rect 252002 266364 252008 266416
rect 252060 266404 252066 266416
rect 257338 266404 257344 266416
rect 252060 266376 257344 266404
rect 252060 266364 252066 266376
rect 257338 266364 257344 266376
rect 257396 266364 257402 266416
rect 263318 266364 263324 266416
rect 263376 266404 263382 266416
rect 265618 266404 265624 266416
rect 263376 266376 265624 266404
rect 263376 266364 263382 266376
rect 265618 266364 265624 266376
rect 265676 266364 265682 266416
rect 269114 266364 269120 266416
rect 269172 266404 269178 266416
rect 276382 266404 276388 266416
rect 269172 266376 276388 266404
rect 269172 266364 269178 266376
rect 276382 266364 276388 266376
rect 276440 266364 276446 266416
rect 278590 266364 278596 266416
rect 278648 266404 278654 266416
rect 286318 266404 286324 266416
rect 278648 266376 286324 266404
rect 278648 266364 278654 266376
rect 286318 266364 286324 266376
rect 286376 266364 286382 266416
rect 290458 266364 290464 266416
rect 290516 266404 290522 266416
rect 292942 266404 292948 266416
rect 290516 266376 292948 266404
rect 290516 266364 290522 266376
rect 292942 266364 292948 266376
rect 293000 266364 293006 266416
rect 297910 266364 297916 266416
rect 297968 266404 297974 266416
rect 299566 266404 299572 266416
rect 297968 266376 299572 266404
rect 297968 266364 297974 266376
rect 299566 266364 299572 266376
rect 299624 266364 299630 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 312354 266364 312360 266416
rect 312412 266404 312418 266416
rect 314654 266404 314660 266416
rect 312412 266376 314660 266404
rect 312412 266364 312418 266376
rect 314654 266364 314660 266376
rect 314712 266364 314718 266416
rect 317782 266364 317788 266416
rect 317840 266404 317846 266416
rect 323118 266404 323124 266416
rect 317840 266376 323124 266404
rect 317840 266364 317846 266376
rect 323118 266364 323124 266376
rect 323176 266364 323182 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329466 266404 329472 266416
rect 328604 266376 329472 266404
rect 328604 266364 328610 266376
rect 329466 266364 329472 266376
rect 329524 266364 329530 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333882 266404 333888 266416
rect 332744 266376 333888 266404
rect 332744 266364 332750 266376
rect 333882 266364 333888 266376
rect 333940 266364 333946 266416
rect 340966 266364 340972 266416
rect 341024 266404 341030 266416
rect 342162 266404 342168 266416
rect 341024 266376 342168 266404
rect 341024 266364 341030 266376
rect 342162 266364 342168 266376
rect 342220 266364 342226 266416
rect 345106 266364 345112 266416
rect 345164 266404 345170 266416
rect 346302 266404 346308 266416
rect 345164 266376 346308 266404
rect 345164 266364 345170 266376
rect 346302 266364 346308 266376
rect 346360 266364 346366 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350258 266404 350264 266416
rect 349304 266376 350264 266404
rect 349304 266364 349310 266376
rect 350258 266364 350264 266376
rect 350316 266364 350322 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 358630 266404 358636 266416
rect 357584 266376 358636 266404
rect 357584 266364 357590 266376
rect 358630 266364 358636 266376
rect 358688 266364 358694 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368382 266404 368388 266416
rect 367520 266376 368388 266404
rect 367520 266364 367526 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375098 266404 375104 266416
rect 374144 266376 375104 266404
rect 374144 266364 374150 266376
rect 375098 266364 375104 266376
rect 375156 266364 375162 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412450 266404 412456 266416
rect 411404 266376 412456 266404
rect 411404 266364 411410 266376
rect 412450 266364 412456 266376
rect 412508 266364 412514 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 423766 266364 423772 266416
rect 423824 266404 423830 266416
rect 424962 266404 424968 266416
rect 423824 266376 424968 266404
rect 423824 266364 423830 266376
rect 424962 266364 424968 266376
rect 425020 266364 425026 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 426894 266404 426900 266416
rect 425480 266376 426900 266404
rect 425480 266364 425486 266376
rect 426894 266364 426900 266376
rect 426952 266364 426958 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 433702 266364 433708 266416
rect 433760 266404 433766 266416
rect 434622 266404 434628 266416
rect 433760 266376 434628 266404
rect 433760 266364 433766 266376
rect 434622 266364 434628 266376
rect 434680 266364 434686 266416
rect 437014 266364 437020 266416
rect 437072 266404 437078 266416
rect 440878 266404 440884 266416
rect 437072 266376 440884 266404
rect 437072 266364 437078 266376
rect 440878 266364 440884 266376
rect 440936 266364 440942 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 447778 266364 447784 266416
rect 447836 266404 447842 266416
rect 449158 266404 449164 266416
rect 447836 266376 449164 266404
rect 447836 266364 447842 266376
rect 449158 266364 449164 266376
rect 449216 266364 449222 266416
rect 451918 266364 451924 266416
rect 451976 266404 451982 266416
rect 454678 266404 454684 266416
rect 451976 266376 454684 266404
rect 451976 266364 451982 266376
rect 454678 266364 454684 266376
rect 454736 266364 454742 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 458082 266404 458088 266416
rect 456944 266376 458088 266404
rect 456944 266364 456950 266376
rect 458082 266364 458088 266376
rect 458140 266364 458146 266416
rect 458542 266364 458548 266416
rect 458600 266404 458606 266416
rect 459370 266404 459376 266416
rect 458600 266376 459376 266404
rect 458600 266364 458606 266376
rect 459370 266364 459376 266376
rect 459428 266364 459434 266416
rect 498562 266296 498568 266348
rect 498620 266336 498626 266348
rect 501598 266336 501604 266348
rect 498620 266308 501604 266336
rect 498620 266296 498626 266308
rect 501598 266296 501604 266308
rect 501656 266296 501662 266348
rect 502794 266296 502800 266348
rect 502852 266336 502858 266348
rect 507854 266336 507860 266348
rect 502852 266308 507860 266336
rect 502852 266296 502858 266308
rect 507854 266296 507860 266308
rect 507912 266296 507918 266348
rect 512196 266336 512224 266444
rect 512362 266432 512368 266484
rect 512420 266472 512426 266484
rect 513374 266472 513380 266484
rect 512420 266444 513380 266472
rect 512420 266432 512426 266444
rect 513374 266432 513380 266444
rect 513432 266432 513438 266484
rect 517330 266432 517336 266484
rect 517388 266472 517394 266484
rect 534276 266472 534304 266580
rect 538674 266568 538680 266580
rect 538732 266568 538738 266620
rect 538858 266568 538864 266620
rect 538916 266608 538922 266620
rect 552676 266608 552704 266716
rect 552842 266704 552848 266756
rect 552900 266744 552906 266756
rect 576826 266744 576854 266852
rect 552900 266716 576854 266744
rect 552900 266704 552906 266716
rect 558914 266608 558920 266620
rect 538916 266580 552612 266608
rect 552676 266580 558920 266608
rect 538916 266568 538922 266580
rect 517388 266444 534304 266472
rect 552584 266472 552612 266580
rect 558914 266568 558920 266580
rect 558972 266568 558978 266620
rect 552842 266472 552848 266484
rect 552584 266444 552848 266472
rect 517388 266432 517394 266444
rect 552842 266432 552848 266444
rect 552900 266432 552906 266484
rect 514662 266404 514668 266416
rect 513576 266376 514668 266404
rect 512196 266308 512316 266336
rect 512288 266268 512316 266308
rect 513576 266268 513604 266376
rect 514662 266364 514668 266376
rect 514720 266364 514726 266416
rect 514846 266364 514852 266416
rect 514904 266404 514910 266416
rect 516778 266404 516784 266416
rect 514904 266376 516784 266404
rect 514904 266364 514910 266376
rect 516778 266364 516784 266376
rect 516836 266364 516842 266416
rect 549622 266404 549628 266416
rect 534368 266376 549628 266404
rect 518802 266296 518808 266348
rect 518860 266336 518866 266348
rect 520274 266336 520280 266348
rect 518860 266308 520280 266336
rect 518860 266296 518866 266308
rect 520274 266296 520280 266308
rect 520332 266296 520338 266348
rect 522666 266296 522672 266348
rect 522724 266336 522730 266348
rect 525886 266336 525892 266348
rect 522724 266308 525892 266336
rect 522724 266296 522730 266308
rect 525886 266296 525892 266308
rect 525944 266296 525950 266348
rect 527634 266296 527640 266348
rect 527692 266336 527698 266348
rect 533890 266336 533896 266348
rect 527692 266308 533896 266336
rect 527692 266296 527698 266308
rect 533890 266296 533896 266308
rect 533948 266296 533954 266348
rect 534074 266296 534080 266348
rect 534132 266336 534138 266348
rect 534368 266336 534396 266376
rect 549622 266364 549628 266376
rect 549680 266364 549686 266416
rect 534132 266308 534396 266336
rect 534132 266296 534138 266308
rect 512288 266240 513604 266268
rect 475102 266024 475108 266076
rect 475160 266064 475166 266076
rect 547874 266064 547880 266076
rect 475160 266036 547880 266064
rect 475160 266024 475166 266036
rect 547874 266024 547880 266036
rect 547932 266024 547938 266076
rect 485038 265888 485044 265940
rect 485096 265928 485102 265940
rect 561674 265928 561680 265940
rect 485096 265900 561680 265928
rect 485096 265888 485102 265900
rect 561674 265888 561680 265900
rect 561732 265888 561738 265940
rect 494974 265752 494980 265804
rect 495032 265792 495038 265804
rect 575842 265792 575848 265804
rect 495032 265764 575848 265792
rect 495032 265752 495038 265764
rect 575842 265752 575848 265764
rect 575900 265752 575906 265804
rect 187694 265616 187700 265668
rect 187752 265656 187758 265668
rect 188246 265656 188252 265668
rect 187752 265628 188252 265656
rect 187752 265616 187758 265628
rect 188246 265616 188252 265628
rect 188304 265616 188310 265668
rect 247218 265616 247224 265668
rect 247276 265656 247282 265668
rect 247862 265656 247868 265668
rect 247276 265628 247868 265656
rect 247276 265616 247282 265628
rect 247862 265616 247868 265628
rect 247920 265616 247926 265668
rect 259546 265616 259552 265668
rect 259604 265656 259610 265668
rect 260374 265656 260380 265668
rect 259604 265628 260380 265656
rect 259604 265616 259610 265628
rect 260374 265616 260380 265628
rect 260432 265616 260438 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 480070 265616 480076 265668
rect 480128 265656 480134 265668
rect 554774 265656 554780 265668
rect 480128 265628 554780 265656
rect 480128 265616 480134 265628
rect 554774 265616 554780 265628
rect 554832 265616 554838 265668
rect 558178 265616 558184 265668
rect 558236 265656 558242 265668
rect 647234 265656 647240 265668
rect 558236 265628 647240 265656
rect 558236 265616 558242 265628
rect 647234 265616 647240 265628
rect 647292 265616 647298 265668
rect 533062 265072 533068 265124
rect 533120 265112 533126 265124
rect 536558 265112 536564 265124
rect 533120 265084 536564 265112
rect 533120 265072 533126 265084
rect 536558 265072 536564 265084
rect 536616 265072 536622 265124
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 567838 259468 567844 259480
rect 554372 259440 567844 259468
rect 554372 259428 554378 259440
rect 567838 259428 567844 259440
rect 567896 259428 567902 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 562318 256748 562324 256760
rect 554004 256720 562324 256748
rect 554004 256708 554010 256720
rect 562318 256708 562324 256720
rect 562376 256708 562382 256760
rect 554498 253376 554504 253428
rect 554556 253416 554562 253428
rect 559558 253416 559564 253428
rect 554556 253388 559564 253416
rect 554556 253376 554562 253388
rect 559558 253376 559564 253388
rect 559616 253376 559622 253428
rect 35802 252832 35808 252884
rect 35860 252872 35866 252884
rect 40678 252872 40684 252884
rect 35860 252844 40684 252872
rect 35860 252832 35866 252844
rect 40678 252832 40684 252844
rect 40736 252832 40742 252884
rect 35618 252696 35624 252748
rect 35676 252736 35682 252748
rect 41690 252736 41696 252748
rect 35676 252708 41696 252736
rect 35676 252696 35682 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35434 252560 35440 252612
rect 35492 252600 35498 252612
rect 41322 252600 41328 252612
rect 35492 252572 41328 252600
rect 35492 252560 35498 252572
rect 41322 252560 41328 252572
rect 41380 252560 41386 252612
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 675846 251540 675852 251592
rect 675904 251580 675910 251592
rect 678422 251580 678428 251592
rect 675904 251552 678428 251580
rect 675904 251540 675910 251552
rect 678422 251540 678428 251552
rect 678480 251540 678486 251592
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 36538 251240 36544 251252
rect 35860 251212 36544 251240
rect 35860 251200 35866 251212
rect 36538 251200 36544 251212
rect 36596 251200 36602 251252
rect 553486 251200 553492 251252
rect 553544 251240 553550 251252
rect 555418 251240 555424 251252
rect 553544 251212 555424 251240
rect 553544 251200 553550 251212
rect 555418 251200 555424 251212
rect 555476 251200 555482 251252
rect 553670 249024 553676 249076
rect 553728 249064 553734 249076
rect 571334 249064 571340 249076
rect 553728 249036 571340 249064
rect 553728 249024 553734 249036
rect 571334 249024 571340 249036
rect 571392 249024 571398 249076
rect 553854 246304 553860 246356
rect 553912 246344 553918 246356
rect 632698 246344 632704 246356
rect 553912 246316 632704 246344
rect 553912 246304 553918 246316
rect 632698 246304 632704 246316
rect 632756 246304 632762 246356
rect 554406 245624 554412 245676
rect 554464 245664 554470 245676
rect 591298 245664 591304 245676
rect 554464 245636 591304 245664
rect 554464 245624 554470 245636
rect 591298 245624 591304 245636
rect 591356 245624 591362 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 624418 244304 624424 244316
rect 554556 244276 624424 244304
rect 554556 244264 554562 244276
rect 624418 244264 624424 244276
rect 624476 244264 624482 244316
rect 36538 242836 36544 242888
rect 36596 242876 36602 242888
rect 41690 242876 41696 242888
rect 36596 242848 41696 242876
rect 36596 242836 36602 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553946 241476 553952 241528
rect 554004 241516 554010 241528
rect 628558 241516 628564 241528
rect 554004 241488 628564 241516
rect 554004 241476 554010 241488
rect 628558 241476 628564 241488
rect 628616 241476 628622 241528
rect 553854 240116 553860 240168
rect 553912 240156 553918 240168
rect 577498 240156 577504 240168
rect 553912 240128 577504 240156
rect 553912 240116 553918 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672166 237804 672172 237856
rect 672224 237844 672230 237856
rect 672756 237844 672784 238102
rect 672224 237816 672784 237844
rect 672224 237804 672230 237816
rect 671338 237600 671344 237652
rect 671396 237640 671402 237652
rect 672874 237640 672902 237898
rect 671396 237612 672902 237640
rect 671396 237600 671402 237612
rect 672966 237436 672994 237694
rect 672092 237408 672994 237436
rect 668762 237328 668768 237380
rect 668820 237368 668826 237380
rect 672092 237368 672120 237408
rect 668820 237340 672120 237368
rect 668820 237328 668826 237340
rect 671522 237192 671528 237244
rect 671580 237232 671586 237244
rect 673104 237232 673132 237490
rect 671580 237204 673132 237232
rect 671580 237192 671586 237204
rect 671614 236988 671620 237040
rect 671672 237028 671678 237040
rect 673196 237028 673224 237286
rect 671672 237000 673224 237028
rect 671672 236988 671678 237000
rect 673178 236716 673184 236768
rect 673236 236756 673242 236768
rect 673316 236756 673344 237082
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673236 236728 673344 236756
rect 673236 236716 673242 236728
rect 673528 236700 673580 236706
rect 673528 236642 673580 236648
rect 673644 236564 673696 236570
rect 673644 236506 673696 236512
rect 673362 236240 673368 236292
rect 673420 236280 673426 236292
rect 673420 236252 673778 236280
rect 673420 236240 673426 236252
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 673298 236036 673304 236088
rect 673356 236076 673362 236088
rect 673356 236048 673900 236076
rect 673356 236036 673362 236048
rect 670344 235912 673992 235940
rect 670344 235748 670372 235912
rect 670326 235696 670332 235748
rect 670384 235696 670390 235748
rect 672442 235696 672448 235748
rect 672500 235736 672506 235748
rect 672500 235708 674114 235736
rect 672500 235696 672506 235708
rect 673472 235504 674222 235532
rect 591298 235220 591304 235272
rect 591356 235260 591362 235272
rect 633618 235260 633624 235272
rect 591356 235232 633624 235260
rect 591356 235220 591362 235232
rect 633618 235220 633624 235232
rect 633676 235220 633682 235272
rect 673472 234784 673500 235504
rect 674190 234948 674196 235000
rect 674248 234988 674254 235000
rect 674324 234988 674352 235314
rect 674248 234960 674352 234988
rect 674248 234948 674254 234960
rect 674438 234796 674466 235110
rect 672644 234756 673500 234784
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 669774 234540 669780 234592
rect 669832 234580 669838 234592
rect 672644 234580 672672 234756
rect 674374 234744 674380 234796
rect 674432 234756 674466 234796
rect 674432 234744 674438 234756
rect 674548 234648 674576 234906
rect 669832 234552 672672 234580
rect 672736 234620 674576 234648
rect 669832 234540 669838 234552
rect 672258 234336 672264 234388
rect 672316 234376 672322 234388
rect 672736 234376 672764 234620
rect 674668 234444 674696 234702
rect 675846 234540 675852 234592
rect 675904 234580 675910 234592
rect 679618 234580 679624 234592
rect 675904 234552 679624 234580
rect 675904 234540 675910 234552
rect 679618 234540 679624 234552
rect 679676 234540 679682 234592
rect 672316 234348 672764 234376
rect 672828 234416 674696 234444
rect 672316 234336 672322 234348
rect 669590 234200 669596 234252
rect 669648 234240 669654 234252
rect 672828 234240 672856 234416
rect 669648 234212 672856 234240
rect 669648 234200 669654 234212
rect 674558 234200 674564 234252
rect 674616 234240 674622 234252
rect 674760 234240 674788 234498
rect 675846 234336 675852 234388
rect 675904 234376 675910 234388
rect 679986 234376 679992 234388
rect 675904 234348 679992 234376
rect 675904 234336 675910 234348
rect 679986 234336 679992 234348
rect 680044 234336 680050 234388
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674616 234212 674788 234240
rect 674616 234200 674622 234212
rect 675846 234200 675852 234252
rect 675904 234240 675910 234252
rect 679802 234240 679808 234252
rect 675904 234212 679808 234240
rect 675904 234200 675910 234212
rect 679802 234200 679808 234212
rect 679860 234200 679866 234252
rect 669130 234064 669136 234116
rect 669188 234104 669194 234116
rect 669188 234076 675004 234104
rect 669188 234064 669194 234076
rect 672994 233928 673000 233980
rect 673052 233968 673058 233980
rect 674926 233968 674932 233980
rect 673052 233940 674932 233968
rect 673052 233928 673058 233940
rect 674926 233928 674932 233940
rect 674984 233928 674990 233980
rect 675846 233928 675852 233980
rect 675904 233968 675910 233980
rect 683482 233968 683488 233980
rect 675904 233940 683488 233968
rect 675904 233928 675910 233940
rect 683482 233928 683488 233940
rect 683540 233928 683546 233980
rect 670786 233588 670792 233640
rect 670844 233628 670850 233640
rect 675108 233628 675136 233886
rect 675236 233708 675288 233714
rect 675236 233650 675288 233656
rect 670844 233600 675136 233628
rect 670844 233588 670850 233600
rect 675846 233520 675852 233572
rect 675904 233560 675910 233572
rect 677778 233560 677784 233572
rect 675904 233532 677784 233560
rect 675904 233520 675910 233532
rect 677778 233520 677784 233532
rect 677836 233520 677842 233572
rect 671062 233452 671068 233504
rect 671120 233492 671126 233504
rect 671120 233464 675372 233492
rect 671120 233452 671126 233464
rect 668302 233180 668308 233232
rect 668360 233220 668366 233232
rect 674190 233220 674196 233232
rect 668360 233192 674196 233220
rect 668360 233180 668366 233192
rect 674190 233180 674196 233192
rect 674248 233180 674254 233232
rect 670878 233044 670884 233096
rect 670936 233084 670942 233096
rect 674742 233084 674748 233096
rect 670936 233056 674748 233084
rect 670936 233044 670942 233056
rect 674742 233044 674748 233056
rect 674800 233044 674806 233096
rect 675478 232608 675484 232620
rect 659626 232580 675484 232608
rect 652018 232500 652024 232552
rect 652076 232540 652082 232552
rect 659626 232540 659654 232580
rect 675478 232568 675484 232580
rect 675536 232568 675542 232620
rect 652076 232512 659654 232540
rect 652076 232500 652082 232512
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 680170 232540 680176 232552
rect 675904 232512 680176 232540
rect 675904 232500 675910 232512
rect 680170 232500 680176 232512
rect 680228 232500 680234 232552
rect 662322 232296 662328 232348
rect 662380 232336 662386 232348
rect 675340 232336 675346 232348
rect 662380 232308 675346 232336
rect 662380 232296 662386 232308
rect 675340 232296 675346 232308
rect 675398 232296 675404 232348
rect 665082 232160 665088 232212
rect 665140 232200 665146 232212
rect 665140 232172 675556 232200
rect 665140 232160 665146 232172
rect 675346 232076 675398 232082
rect 675346 232018 675398 232024
rect 675180 231804 675232 231810
rect 675180 231746 675232 231752
rect 672258 231548 672264 231600
rect 672316 231588 672322 231600
rect 673362 231588 673368 231600
rect 672316 231560 673368 231588
rect 672316 231548 672322 231560
rect 673362 231548 673368 231560
rect 673420 231548 673426 231600
rect 675070 231532 675122 231538
rect 675070 231474 675122 231480
rect 674956 231328 675008 231334
rect 674956 231270 675008 231276
rect 675846 231208 675852 231260
rect 675904 231248 675910 231260
rect 677594 231248 677600 231260
rect 675904 231220 677600 231248
rect 675904 231208 675910 231220
rect 677594 231208 677600 231220
rect 677652 231208 677658 231260
rect 674840 231192 674892 231198
rect 674840 231134 674892 231140
rect 674732 230920 674784 230926
rect 674732 230862 674784 230868
rect 668118 230800 668124 230852
rect 668176 230840 668182 230852
rect 669406 230840 669412 230852
rect 668176 230812 669412 230840
rect 668176 230800 668182 230812
rect 669406 230800 669412 230812
rect 669464 230800 669470 230852
rect 673086 230800 673092 230852
rect 673144 230840 673150 230852
rect 673144 230812 674636 230840
rect 673144 230800 673150 230812
rect 158254 230704 158260 230716
rect 157306 230676 158260 230704
rect 144638 230528 144644 230580
rect 144696 230568 144702 230580
rect 150526 230568 150532 230580
rect 144696 230540 150532 230568
rect 144696 230528 144702 230540
rect 150526 230528 150532 230540
rect 150584 230528 150590 230580
rect 150894 230528 150900 230580
rect 150952 230568 150958 230580
rect 157306 230568 157334 230676
rect 158254 230664 158260 230676
rect 158312 230664 158318 230716
rect 150952 230540 157334 230568
rect 157536 230540 158760 230568
rect 150952 230528 150958 230540
rect 90358 230392 90364 230444
rect 90416 230432 90422 230444
rect 157536 230432 157564 230540
rect 90416 230404 157564 230432
rect 158732 230432 158760 230540
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 161106 230432 161112 230444
rect 158732 230404 161112 230432
rect 90416 230392 90422 230404
rect 161106 230392 161112 230404
rect 161164 230392 161170 230444
rect 161290 230392 161296 230444
rect 161348 230432 161354 230444
rect 215202 230432 215208 230444
rect 161348 230404 215208 230432
rect 161348 230392 161354 230404
rect 215202 230392 215208 230404
rect 215260 230392 215266 230444
rect 223390 230392 223396 230444
rect 223448 230432 223454 230444
rect 271874 230432 271880 230444
rect 223448 230404 271880 230432
rect 223448 230392 223454 230404
rect 271874 230392 271880 230404
rect 271932 230392 271938 230444
rect 274174 230392 274180 230444
rect 274232 230432 274238 230444
rect 307938 230432 307944 230444
rect 274232 230404 307944 230432
rect 274232 230392 274238 230404
rect 307938 230392 307944 230404
rect 307996 230392 308002 230444
rect 312538 230392 312544 230444
rect 312596 230432 312602 230444
rect 315666 230432 315672 230444
rect 312596 230404 315672 230432
rect 312596 230392 312602 230404
rect 315666 230392 315672 230404
rect 315724 230392 315730 230444
rect 377398 230392 377404 230444
rect 377456 230432 377462 230444
rect 378778 230432 378784 230444
rect 377456 230404 378784 230432
rect 377456 230392 377462 230404
rect 378778 230392 378784 230404
rect 378836 230392 378842 230444
rect 439516 230432 439544 230540
rect 674518 230512 674570 230518
rect 674518 230454 674570 230460
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 444466 230392 444472 230444
rect 444524 230432 444530 230444
rect 447594 230432 447600 230444
rect 444524 230404 447600 230432
rect 444524 230392 444530 230404
rect 447594 230392 447600 230404
rect 447652 230392 447658 230444
rect 528002 230392 528008 230444
rect 528060 230432 528066 230444
rect 529014 230432 529020 230444
rect 528060 230404 529020 230432
rect 528060 230392 528066 230404
rect 529014 230392 529020 230404
rect 529072 230392 529078 230444
rect 534626 230392 534632 230444
rect 534684 230432 534690 230444
rect 544194 230432 544200 230444
rect 534684 230404 544200 230432
rect 534684 230392 534690 230404
rect 544194 230392 544200 230404
rect 544252 230392 544258 230444
rect 671798 230392 671804 230444
rect 671856 230432 671862 230444
rect 671856 230404 674422 230432
rect 671856 230392 671862 230404
rect 404262 230324 404268 230376
rect 404320 230364 404326 230376
rect 412266 230364 412272 230376
rect 404320 230336 412272 230364
rect 404320 230324 404326 230336
rect 412266 230324 412272 230336
rect 412324 230324 412330 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 448330 230324 448336 230376
rect 448388 230364 448394 230376
rect 449158 230364 449164 230376
rect 448388 230336 449164 230364
rect 448388 230324 448394 230336
rect 449158 230324 449164 230336
rect 449216 230324 449222 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 475378 230324 475384 230376
rect 475436 230364 475442 230376
rect 478322 230364 478328 230376
rect 475436 230336 478328 230364
rect 475436 230324 475442 230336
rect 478322 230324 478328 230336
rect 478380 230324 478386 230376
rect 480530 230324 480536 230376
rect 480588 230364 480594 230376
rect 481542 230364 481548 230376
rect 480588 230336 481548 230364
rect 480588 230324 480594 230336
rect 481542 230324 481548 230336
rect 481600 230324 481606 230376
rect 492766 230324 492772 230376
rect 492824 230364 492830 230376
rect 493962 230364 493968 230376
rect 492824 230336 493968 230364
rect 492824 230324 492830 230336
rect 493962 230324 493968 230336
rect 494020 230324 494026 230376
rect 513374 230324 513380 230376
rect 513432 230364 513438 230376
rect 515398 230364 515404 230376
rect 513432 230336 515404 230364
rect 513432 230324 513438 230336
rect 515398 230324 515404 230336
rect 515456 230324 515462 230376
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521562 230364 521568 230376
rect 520516 230336 521568 230364
rect 520516 230324 520522 230336
rect 521562 230324 521568 230336
rect 521620 230324 521626 230376
rect 526898 230324 526904 230376
rect 526956 230364 526962 230376
rect 527818 230364 527824 230376
rect 526956 230336 527824 230364
rect 526956 230324 526962 230336
rect 527818 230324 527824 230336
rect 527876 230324 527882 230376
rect 118418 230256 118424 230308
rect 118476 230296 118482 230308
rect 189442 230296 189448 230308
rect 118476 230268 189448 230296
rect 118476 230256 118482 230268
rect 189442 230256 189448 230268
rect 189500 230256 189506 230308
rect 190914 230256 190920 230308
rect 190972 230296 190978 230308
rect 190972 230268 195974 230296
rect 190972 230256 190978 230268
rect 111058 230120 111064 230172
rect 111116 230160 111122 230172
rect 184290 230160 184296 230172
rect 111116 230132 184296 230160
rect 111116 230120 111122 230132
rect 184290 230120 184296 230132
rect 184348 230120 184354 230172
rect 191558 230160 191564 230172
rect 186286 230132 191564 230160
rect 88242 229984 88248 230036
rect 88300 230024 88306 230036
rect 166258 230024 166264 230036
rect 88300 229996 166264 230024
rect 88300 229984 88306 229996
rect 166258 229984 166264 229996
rect 166316 229984 166322 230036
rect 166626 229984 166632 230036
rect 166684 230024 166690 230036
rect 181714 230024 181720 230036
rect 166684 229996 181720 230024
rect 166684 229984 166690 229996
rect 181714 229984 181720 229996
rect 181772 229984 181778 230036
rect 184198 229984 184204 230036
rect 184256 230024 184262 230036
rect 186286 230024 186314 230132
rect 191558 230120 191564 230132
rect 191616 230120 191622 230172
rect 195946 230160 195974 230268
rect 196986 230256 196992 230308
rect 197044 230296 197050 230308
rect 197044 230268 204944 230296
rect 197044 230256 197050 230268
rect 202322 230160 202328 230172
rect 195946 230132 202328 230160
rect 202322 230120 202328 230132
rect 202380 230120 202386 230172
rect 204916 230160 204944 230268
rect 205358 230256 205364 230308
rect 205416 230296 205422 230308
rect 256418 230296 256424 230308
rect 205416 230268 256424 230296
rect 205416 230256 205422 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 276290 230256 276296 230308
rect 276348 230296 276354 230308
rect 313090 230296 313096 230308
rect 276348 230268 313096 230296
rect 276348 230256 276354 230268
rect 313090 230256 313096 230268
rect 313148 230256 313154 230308
rect 323394 230296 323400 230308
rect 313292 230268 323400 230296
rect 251266 230160 251272 230172
rect 204916 230132 251272 230160
rect 251266 230120 251272 230132
rect 251324 230120 251330 230172
rect 261386 230120 261392 230172
rect 261444 230160 261450 230172
rect 297634 230160 297640 230172
rect 261444 230132 297640 230160
rect 261444 230120 261450 230132
rect 297634 230120 297640 230132
rect 297692 230120 297698 230172
rect 308122 230120 308128 230172
rect 308180 230160 308186 230172
rect 313292 230160 313320 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 436094 230256 436100 230308
rect 436152 230296 436158 230308
rect 436830 230296 436836 230308
rect 436152 230268 436836 230296
rect 436152 230256 436158 230268
rect 436830 230256 436836 230268
rect 436888 230256 436894 230308
rect 497918 230256 497924 230308
rect 497976 230296 497982 230308
rect 504358 230296 504364 230308
rect 497976 230268 504364 230296
rect 497976 230256 497982 230268
rect 504358 230256 504364 230268
rect 504416 230256 504422 230308
rect 528830 230256 528836 230308
rect 528888 230296 528894 230308
rect 541618 230296 541624 230308
rect 528888 230268 541624 230296
rect 528888 230256 528894 230268
rect 541618 230256 541624 230268
rect 541676 230256 541682 230308
rect 408862 230188 408868 230240
rect 408920 230228 408926 230240
rect 410978 230228 410984 230240
rect 408920 230200 410984 230228
rect 408920 230188 408926 230200
rect 410978 230188 410984 230200
rect 411036 230188 411042 230240
rect 443822 230188 443828 230240
rect 443880 230228 443886 230240
rect 444650 230228 444656 230240
rect 443880 230200 444656 230228
rect 443880 230188 443886 230200
rect 444650 230188 444656 230200
rect 444708 230188 444714 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 454126 230188 454132 230240
rect 454184 230228 454190 230240
rect 455230 230228 455236 230240
rect 454184 230200 455236 230228
rect 454184 230188 454190 230200
rect 455230 230188 455236 230200
rect 455288 230188 455294 230240
rect 470870 230188 470876 230240
rect 470928 230228 470934 230240
rect 471882 230228 471888 230240
rect 470928 230200 471888 230228
rect 470928 230188 470934 230200
rect 471882 230188 471888 230200
rect 471940 230188 471946 230240
rect 476666 230188 476672 230240
rect 476724 230228 476730 230240
rect 479702 230228 479708 230240
rect 476724 230200 479708 230228
rect 476724 230188 476730 230200
rect 479702 230188 479708 230200
rect 479760 230188 479766 230240
rect 493410 230188 493416 230240
rect 493468 230228 493474 230240
rect 495158 230228 495164 230240
rect 493468 230200 495164 230228
rect 493468 230188 493474 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 516502 230228 516508 230240
rect 511500 230200 516508 230228
rect 511500 230188 511506 230200
rect 516502 230188 516508 230200
rect 516560 230188 516566 230240
rect 668118 230188 668124 230240
rect 668176 230228 668182 230240
rect 674098 230228 674104 230240
rect 668176 230200 674104 230228
rect 668176 230188 668182 230200
rect 674098 230188 674104 230200
rect 674156 230188 674162 230240
rect 308180 230132 313320 230160
rect 308180 230120 308186 230132
rect 315298 230120 315304 230172
rect 315356 230160 315362 230172
rect 340138 230160 340144 230172
rect 315356 230132 340144 230160
rect 315356 230120 315362 230132
rect 340138 230120 340144 230132
rect 340196 230120 340202 230172
rect 503254 230160 503260 230172
rect 499546 230132 503260 230160
rect 302878 230052 302884 230104
rect 302936 230092 302942 230104
rect 305362 230092 305368 230104
rect 302936 230064 305368 230092
rect 302936 230052 302942 230064
rect 305362 230052 305368 230064
rect 305420 230052 305426 230104
rect 345658 230052 345664 230104
rect 345716 230092 345722 230104
rect 353018 230092 353024 230104
rect 345716 230064 353024 230092
rect 345716 230052 345722 230064
rect 353018 230052 353024 230064
rect 353076 230052 353082 230104
rect 453482 230052 453488 230104
rect 453540 230092 453546 230104
rect 455782 230092 455788 230104
rect 453540 230064 455788 230092
rect 453540 230052 453546 230064
rect 455782 230052 455788 230064
rect 455840 230052 455846 230104
rect 476022 230052 476028 230104
rect 476080 230092 476086 230104
rect 479518 230092 479524 230104
rect 476080 230064 479524 230092
rect 476080 230052 476086 230064
rect 479518 230052 479524 230064
rect 479576 230052 479582 230104
rect 490834 230052 490840 230104
rect 490892 230092 490898 230104
rect 493778 230092 493784 230104
rect 490892 230064 493784 230092
rect 490892 230052 490898 230064
rect 493778 230052 493784 230064
rect 493836 230052 493842 230104
rect 494330 230052 494336 230104
rect 494388 230092 494394 230104
rect 499546 230092 499574 230132
rect 503254 230120 503260 230132
rect 503312 230120 503318 230172
rect 521102 230120 521108 230172
rect 521160 230160 521166 230172
rect 529934 230160 529940 230172
rect 521160 230132 529940 230160
rect 521160 230120 521166 230132
rect 529934 230120 529940 230132
rect 529992 230120 529998 230172
rect 536558 230120 536564 230172
rect 536616 230160 536622 230172
rect 549254 230160 549260 230172
rect 536616 230132 549260 230160
rect 536616 230120 536622 230132
rect 549254 230120 549260 230132
rect 549312 230120 549318 230172
rect 494388 230064 499574 230092
rect 494388 230052 494394 230064
rect 674282 230052 674288 230104
rect 674340 230052 674346 230104
rect 184256 229996 186314 230024
rect 184256 229984 184262 229996
rect 190178 229984 190184 230036
rect 190236 230024 190242 230036
rect 246114 230024 246120 230036
rect 190236 229996 246120 230024
rect 190236 229984 190242 229996
rect 246114 229984 246120 229996
rect 246172 229984 246178 230036
rect 251726 229984 251732 230036
rect 251784 230024 251790 230036
rect 292482 230024 292488 230036
rect 251784 229996 292488 230024
rect 251784 229984 251790 229996
rect 292482 229984 292488 229996
rect 292540 229984 292546 230036
rect 296990 229984 296996 230036
rect 297048 230024 297054 230036
rect 302510 230024 302516 230036
rect 297048 229996 302516 230024
rect 297048 229984 297054 229996
rect 302510 229984 302516 229996
rect 302568 229984 302574 230036
rect 305638 229984 305644 230036
rect 305696 230024 305702 230036
rect 334986 230024 334992 230036
rect 305696 229996 334992 230024
rect 305696 229984 305702 229996
rect 334986 229984 334992 229996
rect 335044 229984 335050 230036
rect 380434 229984 380440 230036
rect 380492 230024 380498 230036
rect 389082 230024 389088 230036
rect 380492 229996 389088 230024
rect 380492 229984 380498 229996
rect 389082 229984 389088 229996
rect 389140 229984 389146 230036
rect 410886 229984 410892 230036
rect 410944 230024 410950 230036
rect 417418 230024 417424 230036
rect 410944 229996 417424 230024
rect 410944 229984 410950 229996
rect 417418 229984 417424 229996
rect 417476 229984 417482 230036
rect 447042 229984 447048 230036
rect 447100 230024 447106 230036
rect 449894 230024 449900 230036
rect 447100 229996 449900 230024
rect 447100 229984 447106 229996
rect 449894 229984 449900 229996
rect 449952 229984 449958 230036
rect 467006 229984 467012 230036
rect 467064 230024 467070 230036
rect 473998 230024 474004 230036
rect 467064 229996 474004 230024
rect 467064 229984 467070 229996
rect 473998 229984 474004 229996
rect 474056 229984 474062 230036
rect 483106 229984 483112 230036
rect 483164 230024 483170 230036
rect 484302 230024 484308 230036
rect 483164 229996 484308 230024
rect 483164 229984 483170 229996
rect 484302 229984 484308 229996
rect 484360 229984 484366 230036
rect 484762 229984 484768 230036
rect 484820 230024 484826 230036
rect 490650 230024 490656 230036
rect 484820 229996 490656 230024
rect 484820 229984 484826 229996
rect 490650 229984 490656 229996
rect 490708 229984 490714 230036
rect 503714 229984 503720 230036
rect 503772 230024 503778 230036
rect 506934 230024 506940 230036
rect 503772 229996 506940 230024
rect 503772 229984 503778 229996
rect 506934 229984 506940 229996
rect 506992 229984 506998 230036
rect 509510 229984 509516 230036
rect 509568 230024 509574 230036
rect 518894 230024 518900 230036
rect 509568 229996 518900 230024
rect 509568 229984 509574 229996
rect 518894 229984 518900 229996
rect 518952 229984 518958 230036
rect 519170 229984 519176 230036
rect 519228 230024 519234 230036
rect 528002 230024 528008 230036
rect 519228 229996 528008 230024
rect 519228 229984 519234 229996
rect 528002 229984 528008 229996
rect 528060 229984 528066 230036
rect 530762 229984 530768 230036
rect 530820 230024 530826 230036
rect 547138 230024 547144 230036
rect 530820 229996 547144 230024
rect 530820 229984 530826 229996
rect 547138 229984 547144 229996
rect 547196 229984 547202 230036
rect 555418 229984 555424 230036
rect 555476 230024 555482 230036
rect 569954 230024 569960 230036
rect 555476 229996 569960 230024
rect 555476 229984 555482 229996
rect 569954 229984 569960 229996
rect 570012 229984 570018 230036
rect 675846 229984 675852 230036
rect 675904 230024 675910 230036
rect 676582 230024 676588 230036
rect 675904 229996 676588 230024
rect 675904 229984 675910 229996
rect 676582 229984 676588 229996
rect 676640 229984 676646 230036
rect 674172 229968 674224 229974
rect 674172 229910 674224 229916
rect 674058 229900 674110 229906
rect 74442 229848 74448 229900
rect 74500 229888 74506 229900
rect 155954 229888 155960 229900
rect 74500 229860 155960 229888
rect 74500 229848 74506 229860
rect 155954 229848 155960 229860
rect 156012 229848 156018 229900
rect 156322 229848 156328 229900
rect 156380 229888 156386 229900
rect 176562 229888 176568 229900
rect 156380 229860 176568 229888
rect 156380 229848 156386 229860
rect 176562 229848 176568 229860
rect 176620 229848 176626 229900
rect 177574 229848 177580 229900
rect 177632 229888 177638 229900
rect 177632 229860 191144 229888
rect 177632 229848 177638 229860
rect 67542 229712 67548 229764
rect 67600 229752 67606 229764
rect 144638 229752 144644 229764
rect 67600 229724 144644 229752
rect 67600 229712 67606 229724
rect 144638 229712 144644 229724
rect 144696 229712 144702 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 144880 229724 147168 229752
rect 144880 229712 144886 229724
rect 140038 229576 140044 229628
rect 140096 229616 140102 229628
rect 146938 229616 146944 229628
rect 140096 229588 146944 229616
rect 140096 229576 140102 229588
rect 146938 229576 146944 229588
rect 146996 229576 147002 229628
rect 147140 229616 147168 229724
rect 148594 229712 148600 229764
rect 148652 229752 148658 229764
rect 150894 229752 150900 229764
rect 148652 229724 150900 229752
rect 148652 229712 148658 229724
rect 150894 229712 150900 229724
rect 150952 229712 150958 229764
rect 151354 229712 151360 229764
rect 151412 229752 151418 229764
rect 190914 229752 190920 229764
rect 151412 229724 190920 229752
rect 151412 229712 151418 229724
rect 190914 229712 190920 229724
rect 190972 229712 190978 229764
rect 191116 229752 191144 229860
rect 191558 229848 191564 229900
rect 191616 229888 191622 229900
rect 240962 229888 240968 229900
rect 191616 229860 240968 229888
rect 191616 229848 191622 229860
rect 240962 229848 240968 229860
rect 241020 229848 241026 229900
rect 245654 229848 245660 229900
rect 245712 229888 245718 229900
rect 287330 229888 287336 229900
rect 245712 229860 287336 229888
rect 245712 229848 245718 229860
rect 287330 229848 287336 229860
rect 287388 229848 287394 229900
rect 300118 229848 300124 229900
rect 300176 229888 300182 229900
rect 329834 229888 329840 229900
rect 300176 229860 329840 229888
rect 300176 229848 300182 229860
rect 329834 229848 329840 229860
rect 329892 229848 329898 229900
rect 334250 229848 334256 229900
rect 334308 229888 334314 229900
rect 345290 229888 345296 229900
rect 334308 229860 345296 229888
rect 334308 229848 334314 229860
rect 345290 229848 345296 229860
rect 345348 229848 345354 229900
rect 352558 229848 352564 229900
rect 352616 229888 352622 229900
rect 358170 229888 358176 229900
rect 352616 229860 358176 229888
rect 352616 229848 352622 229860
rect 358170 229848 358176 229860
rect 358228 229848 358234 229900
rect 364150 229848 364156 229900
rect 364208 229888 364214 229900
rect 381354 229888 381360 229900
rect 364208 229860 381360 229888
rect 364208 229848 364214 229860
rect 381354 229848 381360 229860
rect 381412 229848 381418 229900
rect 384298 229848 384304 229900
rect 384356 229888 384362 229900
rect 394234 229888 394240 229900
rect 384356 229860 394240 229888
rect 384356 229848 384362 229860
rect 394234 229848 394240 229860
rect 394292 229848 394298 229900
rect 468938 229848 468944 229900
rect 468996 229888 469002 229900
rect 468996 229860 469444 229888
rect 468996 229848 469002 229860
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 235810 229752 235816 229764
rect 191116 229724 235816 229752
rect 235810 229712 235816 229724
rect 235868 229712 235874 229764
rect 236914 229712 236920 229764
rect 236972 229752 236978 229764
rect 282178 229752 282184 229764
rect 236972 229724 282184 229752
rect 236972 229712 236978 229724
rect 282178 229712 282184 229724
rect 282236 229712 282242 229764
rect 285306 229712 285312 229764
rect 285364 229752 285370 229764
rect 318242 229752 318248 229764
rect 285364 229724 318248 229752
rect 285364 229712 285370 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 324038 229712 324044 229764
rect 324096 229752 324102 229764
rect 350442 229752 350448 229764
rect 324096 229724 350448 229752
rect 324096 229712 324102 229724
rect 350442 229712 350448 229724
rect 350500 229712 350506 229764
rect 371050 229752 371056 229764
rect 354646 229724 371056 229752
rect 210050 229616 210056 229628
rect 147140 229588 210056 229616
rect 210050 229576 210056 229588
rect 210108 229576 210114 229628
rect 210234 229576 210240 229628
rect 210292 229616 210298 229628
rect 261570 229616 261576 229628
rect 210292 229588 261576 229616
rect 210292 229576 210298 229588
rect 261570 229576 261576 229588
rect 261628 229576 261634 229628
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 354646 229616 354674 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 386506 229752 386512 229764
rect 373966 229724 386512 229752
rect 350592 229588 354674 229616
rect 350592 229576 350598 229588
rect 370958 229576 370964 229628
rect 371016 229616 371022 229628
rect 373966 229616 373994 229724
rect 386506 229712 386512 229724
rect 386564 229712 386570 229764
rect 386966 229712 386972 229764
rect 387024 229752 387030 229764
rect 396810 229752 396816 229764
rect 387024 229724 396816 229752
rect 387024 229712 387030 229724
rect 396810 229712 396816 229724
rect 396868 229712 396874 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 412450 229712 412456 229764
rect 412508 229752 412514 229764
rect 419350 229752 419356 229764
rect 412508 229724 419356 229752
rect 412508 229712 412514 229724
rect 419350 229712 419356 229724
rect 419408 229712 419414 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 468294 229712 468300 229764
rect 468352 229752 468358 229764
rect 469122 229752 469128 229764
rect 468352 229724 469128 229752
rect 468352 229712 468358 229724
rect 469122 229712 469128 229724
rect 469180 229712 469186 229764
rect 469416 229752 469444 229860
rect 469582 229848 469588 229900
rect 469640 229888 469646 229900
rect 476758 229888 476764 229900
rect 469640 229860 476764 229888
rect 469640 229848 469646 229860
rect 476758 229848 476764 229860
rect 476816 229848 476822 229900
rect 479242 229848 479248 229900
rect 479300 229888 479306 229900
rect 484026 229888 484032 229900
rect 479300 229860 484032 229888
rect 479300 229848 479306 229860
rect 484026 229848 484032 229860
rect 484084 229848 484090 229900
rect 486326 229848 486332 229900
rect 486384 229888 486390 229900
rect 500218 229888 500224 229900
rect 486384 229860 500224 229888
rect 486384 229848 486390 229860
rect 500218 229848 500224 229860
rect 500276 229848 500282 229900
rect 505646 229848 505652 229900
rect 505704 229888 505710 229900
rect 516042 229888 516048 229900
rect 505704 229860 516048 229888
rect 505704 229848 505710 229860
rect 516042 229848 516048 229860
rect 516100 229848 516106 229900
rect 517422 229848 517428 229900
rect 517480 229888 517486 229900
rect 522298 229888 522304 229900
rect 517480 229860 522304 229888
rect 517480 229848 517486 229860
rect 522298 229848 522304 229860
rect 522356 229848 522362 229900
rect 523034 229848 523040 229900
rect 523092 229888 523098 229900
rect 534718 229888 534724 229900
rect 523092 229860 534724 229888
rect 523092 229848 523098 229860
rect 534718 229848 534724 229860
rect 534776 229848 534782 229900
rect 538490 229848 538496 229900
rect 538548 229888 538554 229900
rect 556798 229888 556804 229900
rect 538548 229860 556804 229888
rect 538548 229848 538554 229860
rect 556798 229848 556804 229860
rect 556856 229848 556862 229900
rect 675846 229848 675852 229900
rect 675904 229888 675910 229900
rect 677226 229888 677232 229900
rect 675904 229860 677232 229888
rect 675904 229848 675910 229860
rect 677226 229848 677232 229860
rect 677284 229848 677290 229900
rect 674058 229842 674110 229848
rect 475378 229752 475384 229764
rect 469416 229724 475384 229752
rect 475378 229712 475384 229724
rect 475436 229712 475442 229764
rect 481818 229712 481824 229764
rect 481876 229752 481882 229764
rect 489914 229752 489920 229764
rect 481876 229724 489920 229752
rect 481876 229712 481882 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 495986 229712 495992 229764
rect 496044 229752 496050 229764
rect 509234 229752 509240 229764
rect 496044 229724 509240 229752
rect 496044 229712 496050 229724
rect 509234 229712 509240 229724
rect 509292 229712 509298 229764
rect 515674 229712 515680 229764
rect 515732 229752 515738 229764
rect 525518 229752 525524 229764
rect 515732 229724 525524 229752
rect 515732 229712 515738 229724
rect 525518 229712 525524 229724
rect 525576 229712 525582 229764
rect 532694 229712 532700 229764
rect 532752 229752 532758 229764
rect 555602 229752 555608 229764
rect 532752 229724 555608 229752
rect 532752 229712 532758 229724
rect 555602 229712 555608 229724
rect 555660 229712 555666 229764
rect 675846 229712 675852 229764
rect 675904 229752 675910 229764
rect 676950 229752 676956 229764
rect 675904 229724 676956 229752
rect 675904 229712 675910 229724
rect 676950 229712 676956 229724
rect 677008 229712 677014 229764
rect 371016 229588 373994 229616
rect 371016 229576 371022 229588
rect 455414 229576 455420 229628
rect 455472 229616 455478 229628
rect 457162 229616 457168 229628
rect 455472 229588 457168 229616
rect 455472 229576 455478 229588
rect 457162 229576 457168 229588
rect 457220 229576 457226 229628
rect 490650 229576 490656 229628
rect 490708 229616 490714 229628
rect 497458 229616 497464 229628
rect 490708 229588 497464 229616
rect 490708 229576 490714 229588
rect 497458 229576 497464 229588
rect 497516 229576 497522 229628
rect 524966 229576 524972 229628
rect 525024 229616 525030 229628
rect 532418 229616 532424 229628
rect 525024 229588 532424 229616
rect 525024 229576 525030 229588
rect 532418 229576 532424 229588
rect 532476 229576 532482 229628
rect 673948 229560 674000 229566
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451366 229548 451372 229560
rect 449032 229520 451372 229548
rect 449032 229508 449038 229520
rect 451366 229508 451372 229520
rect 451424 229508 451430 229560
rect 673948 229502 674000 229508
rect 131114 229440 131120 229492
rect 131172 229480 131178 229492
rect 197170 229480 197176 229492
rect 131172 229452 197176 229480
rect 131172 229440 131178 229452
rect 197170 229440 197176 229452
rect 197228 229440 197234 229492
rect 203886 229440 203892 229492
rect 203944 229480 203950 229492
rect 205358 229480 205364 229492
rect 203944 229452 205364 229480
rect 203944 229440 203950 229452
rect 205358 229440 205364 229452
rect 205416 229440 205422 229492
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 277026 229480 277032 229492
rect 231176 229452 277032 229480
rect 231176 229440 231182 229452
rect 277026 229440 277032 229452
rect 277084 229440 277090 229492
rect 499850 229440 499856 229492
rect 499908 229480 499914 229492
rect 501322 229480 501328 229492
rect 499908 229452 501328 229480
rect 499908 229440 499914 229452
rect 501322 229440 501328 229452
rect 501380 229440 501386 229492
rect 673454 229440 673460 229492
rect 673512 229480 673518 229492
rect 673512 229452 673854 229480
rect 673512 229440 673518 229452
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448606 229412 448612 229424
rect 446456 229384 448612 229412
rect 446456 229372 446462 229384
rect 448606 229372 448612 229384
rect 448664 229372 448670 229424
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 453022 229412 453028 229424
rect 450964 229384 453028 229412
rect 450964 229372 450970 229384
rect 453022 229372 453028 229384
rect 453080 229372 453086 229424
rect 501782 229372 501788 229424
rect 501840 229412 501846 229424
rect 507118 229412 507124 229424
rect 501840 229384 507124 229412
rect 501840 229372 501846 229384
rect 507118 229372 507124 229384
rect 507176 229372 507182 229424
rect 92474 229304 92480 229356
rect 92532 229344 92538 229356
rect 146294 229344 146300 229356
rect 92532 229316 146300 229344
rect 92532 229304 92538 229316
rect 146294 229304 146300 229316
rect 146352 229304 146358 229356
rect 146938 229304 146944 229356
rect 146996 229344 147002 229356
rect 153378 229344 153384 229356
rect 146996 229316 153384 229344
rect 146996 229304 147002 229316
rect 153378 229304 153384 229316
rect 153436 229304 153442 229356
rect 153838 229304 153844 229356
rect 153896 229344 153902 229356
rect 163682 229344 163688 229356
rect 153896 229316 163688 229344
rect 153896 229304 153902 229316
rect 163682 229304 163688 229316
rect 163740 229304 163746 229356
rect 163866 229304 163872 229356
rect 163924 229344 163930 229356
rect 166626 229344 166632 229356
rect 163924 229316 166632 229344
rect 163924 229304 163930 229316
rect 166626 229304 166632 229316
rect 166684 229304 166690 229356
rect 167638 229304 167644 229356
rect 167696 229344 167702 229356
rect 220354 229344 220360 229356
rect 167696 229316 220360 229344
rect 167696 229304 167702 229316
rect 220354 229304 220360 229316
rect 220412 229304 220418 229356
rect 494698 229304 494704 229356
rect 494756 229344 494762 229356
rect 496354 229344 496360 229356
rect 494756 229316 496360 229344
rect 494756 229304 494762 229316
rect 496354 229304 496360 229316
rect 496412 229304 496418 229356
rect 673086 229304 673092 229356
rect 673144 229344 673150 229356
rect 673144 229316 673428 229344
rect 673144 229304 673150 229316
rect 358078 229236 358084 229288
rect 358136 229276 358142 229288
rect 360746 229276 360752 229288
rect 358136 229248 360752 229276
rect 358136 229236 358142 229248
rect 360746 229236 360752 229248
rect 360804 229236 360810 229288
rect 360930 229236 360936 229288
rect 360988 229276 360994 229288
rect 363322 229276 363328 229288
rect 360988 229248 363328 229276
rect 360988 229236 360994 229248
rect 363322 229236 363328 229248
rect 363380 229236 363386 229288
rect 419442 229236 419448 229288
rect 419500 229276 419506 229288
rect 424502 229276 424508 229288
rect 419500 229248 424508 229276
rect 419500 229236 419506 229248
rect 424502 229236 424508 229248
rect 424560 229236 424566 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451826 229276 451832 229288
rect 450320 229248 451832 229276
rect 450320 229236 450326 229248
rect 451826 229236 451832 229248
rect 451884 229236 451890 229288
rect 479886 229236 479892 229288
rect 479944 229276 479950 229288
rect 482278 229276 482284 229288
rect 479944 229248 482284 229276
rect 479944 229236 479950 229248
rect 482278 229236 482284 229248
rect 482336 229236 482342 229288
rect 483750 229236 483756 229288
rect 483808 229276 483814 229288
rect 486786 229276 486792 229288
rect 483808 229248 486792 229276
rect 483808 229236 483814 229248
rect 486786 229236 486792 229248
rect 486844 229236 486850 229288
rect 673400 229276 673428 229316
rect 673400 229248 673762 229276
rect 115750 229168 115756 229220
rect 115808 229208 115814 229220
rect 115808 229180 115934 229208
rect 115808 229168 115814 229180
rect 106182 229032 106188 229084
rect 106240 229072 106246 229084
rect 115906 229072 115934 229180
rect 122926 229168 122932 229220
rect 122984 229208 122990 229220
rect 179138 229208 179144 229220
rect 122984 229180 179144 229208
rect 122984 229168 122990 229180
rect 179138 229168 179144 229180
rect 179196 229168 179202 229220
rect 181622 229168 181628 229220
rect 181680 229208 181686 229220
rect 230658 229208 230664 229220
rect 181680 229180 230664 229208
rect 181680 229168 181686 229180
rect 230658 229168 230664 229180
rect 230716 229168 230722 229220
rect 669314 229168 669320 229220
rect 669372 229208 669378 229220
rect 673270 229208 673276 229220
rect 669372 229180 673276 229208
rect 669372 229168 669378 229180
rect 673270 229168 673276 229180
rect 673328 229168 673334 229220
rect 675846 229168 675852 229220
rect 675904 229208 675910 229220
rect 675904 229180 677456 229208
rect 675904 229168 675910 229180
rect 378962 229100 378968 229152
rect 379020 229140 379026 229152
rect 383930 229140 383936 229152
rect 379020 229112 383936 229140
rect 379020 229100 379026 229112
rect 383930 229100 383936 229112
rect 383988 229100 383994 229152
rect 419994 229140 420000 229152
rect 418126 229112 420000 229140
rect 116026 229072 116032 229084
rect 106240 229044 115796 229072
rect 115906 229044 116032 229072
rect 106240 229032 106246 229044
rect 97902 228896 97908 228948
rect 97960 228936 97966 228948
rect 97960 228908 106872 228936
rect 97960 228896 97966 228908
rect 106642 228800 106648 228812
rect 84166 228772 106648 228800
rect 82078 228624 82084 228676
rect 82136 228664 82142 228676
rect 84166 228664 84194 228772
rect 106642 228760 106648 228772
rect 106700 228760 106706 228812
rect 106844 228800 106872 228908
rect 107010 228896 107016 228948
rect 107068 228936 107074 228948
rect 115566 228936 115572 228948
rect 107068 228908 115572 228936
rect 107068 228896 107074 228908
rect 115566 228896 115572 228908
rect 115624 228896 115630 228948
rect 115768 228936 115796 229044
rect 116026 229032 116032 229044
rect 116084 229032 116090 229084
rect 179782 229072 179788 229084
rect 116228 229044 179788 229072
rect 116228 228936 116256 229044
rect 179782 229032 179788 229044
rect 179840 229032 179846 229084
rect 180610 229032 180616 229084
rect 180668 229072 180674 229084
rect 180668 229044 185164 229072
rect 180668 229032 180674 229044
rect 115768 228908 116256 228936
rect 116394 228896 116400 228948
rect 116452 228936 116458 228948
rect 184934 228936 184940 228948
rect 116452 228908 184940 228936
rect 116452 228896 116458 228908
rect 184934 228896 184940 228908
rect 184992 228896 184998 228948
rect 185136 228936 185164 229044
rect 185670 229032 185676 229084
rect 185728 229072 185734 229084
rect 185728 229044 190224 229072
rect 185728 229032 185734 229044
rect 190196 228936 190224 229044
rect 190362 229032 190368 229084
rect 190420 229072 190426 229084
rect 194594 229072 194600 229084
rect 190420 229044 194600 229072
rect 190420 229032 190426 229044
rect 194594 229032 194600 229044
rect 194652 229032 194658 229084
rect 195698 229032 195704 229084
rect 195756 229072 195762 229084
rect 250622 229072 250628 229084
rect 195756 229044 250628 229072
rect 195756 229032 195762 229044
rect 250622 229032 250628 229044
rect 250680 229032 250686 229084
rect 259270 229032 259276 229084
rect 259328 229072 259334 229084
rect 298278 229072 298284 229084
rect 259328 229044 298284 229072
rect 259328 229032 259334 229044
rect 298278 229032 298284 229044
rect 298336 229032 298342 229084
rect 413830 229032 413836 229084
rect 413888 229072 413894 229084
rect 418126 229072 418154 229112
rect 419994 229100 420000 229112
rect 420052 229100 420058 229152
rect 420178 229100 420184 229152
rect 420236 229140 420242 229152
rect 421926 229140 421932 229152
rect 420236 229112 421932 229140
rect 420236 229100 420242 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 424318 229100 424324 229152
rect 424376 229140 424382 229152
rect 427722 229140 427728 229152
rect 424376 229112 427728 229140
rect 424376 229100 424382 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 507578 229100 507584 229152
rect 507636 229140 507642 229152
rect 511258 229140 511264 229152
rect 507636 229112 511264 229140
rect 507636 229100 507642 229112
rect 511258 229100 511264 229112
rect 511316 229100 511322 229152
rect 677428 229084 677456 229180
rect 413888 229044 418154 229072
rect 413888 229032 413894 229044
rect 517882 229032 517888 229084
rect 517940 229072 517946 229084
rect 540238 229072 540244 229084
rect 517940 229044 540244 229072
rect 517940 229032 517946 229044
rect 540238 229032 540244 229044
rect 540296 229032 540302 229084
rect 673454 229032 673460 229084
rect 673512 229072 673518 229084
rect 673512 229044 673624 229072
rect 673512 229032 673518 229044
rect 675846 229032 675852 229084
rect 675904 229072 675910 229084
rect 677042 229072 677048 229084
rect 675904 229044 677048 229072
rect 675904 229032 675910 229044
rect 677042 229032 677048 229044
rect 677100 229032 677106 229084
rect 677410 229032 677416 229084
rect 677468 229032 677474 229084
rect 241606 228936 241612 228948
rect 185136 228908 190132 228936
rect 190196 228908 241612 228936
rect 173986 228800 173992 228812
rect 106844 228772 173992 228800
rect 173986 228760 173992 228772
rect 174044 228760 174050 228812
rect 174170 228760 174176 228812
rect 174228 228800 174234 228812
rect 174228 228772 175596 228800
rect 174228 228760 174234 228772
rect 82136 228636 84194 228664
rect 82136 228624 82142 228636
rect 96246 228624 96252 228676
rect 96304 228664 96310 228676
rect 172054 228664 172060 228676
rect 96304 228636 172060 228664
rect 96304 228624 96310 228636
rect 172054 228624 172060 228636
rect 172112 228624 172118 228676
rect 172238 228624 172244 228676
rect 172296 228664 172302 228676
rect 175274 228664 175280 228676
rect 172296 228636 175280 228664
rect 172296 228624 172302 228636
rect 175274 228624 175280 228636
rect 175332 228624 175338 228676
rect 175568 228664 175596 228772
rect 175734 228760 175740 228812
rect 175792 228800 175798 228812
rect 188338 228800 188344 228812
rect 175792 228772 188344 228800
rect 175792 228760 175798 228772
rect 188338 228760 188344 228772
rect 188396 228760 188402 228812
rect 190104 228800 190132 228908
rect 241606 228896 241612 228908
rect 241664 228896 241670 228948
rect 251082 228896 251088 228948
rect 251140 228936 251146 228948
rect 291194 228936 291200 228948
rect 251140 228908 291200 228936
rect 251140 228896 251146 228908
rect 291194 228896 291200 228908
rect 291252 228896 291258 228948
rect 319806 228896 319812 228948
rect 319864 228936 319870 228948
rect 345934 228936 345940 228948
rect 319864 228908 345940 228936
rect 319864 228896 319870 228908
rect 345934 228896 345940 228908
rect 345992 228896 345998 228948
rect 350166 228896 350172 228948
rect 350224 228936 350230 228948
rect 369118 228936 369124 228948
rect 350224 228908 369124 228936
rect 350224 228896 350230 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 507118 228896 507124 228948
rect 507176 228936 507182 228948
rect 520182 228936 520188 228948
rect 507176 228908 520188 228936
rect 507176 228896 507182 228908
rect 520182 228896 520188 228908
rect 520240 228896 520246 228948
rect 526254 228896 526260 228948
rect 526312 228936 526318 228948
rect 551646 228936 551652 228948
rect 526312 228908 551652 228936
rect 526312 228896 526318 228908
rect 551646 228896 551652 228908
rect 551704 228896 551710 228948
rect 673506 228880 673558 228886
rect 673506 228822 673558 228828
rect 204714 228800 204720 228812
rect 190104 228772 204720 228800
rect 204714 228760 204720 228772
rect 204772 228760 204778 228812
rect 204898 228760 204904 228812
rect 204956 228800 204962 228812
rect 210694 228800 210700 228812
rect 204956 228772 210700 228800
rect 204956 228760 204962 228772
rect 210694 228760 210700 228772
rect 210752 228760 210758 228812
rect 214098 228760 214104 228812
rect 214156 228800 214162 228812
rect 218422 228800 218428 228812
rect 214156 228772 218428 228800
rect 214156 228760 214162 228772
rect 218422 228760 218428 228772
rect 218480 228760 218486 228812
rect 219342 228760 219348 228812
rect 219400 228800 219406 228812
rect 224034 228800 224040 228812
rect 219400 228772 224040 228800
rect 219400 228760 219406 228772
rect 224034 228760 224040 228772
rect 224092 228760 224098 228812
rect 231302 228800 231308 228812
rect 224236 228772 231308 228800
rect 224236 228664 224264 228772
rect 231302 228760 231308 228772
rect 231360 228760 231366 228812
rect 246298 228760 246304 228812
rect 246356 228800 246362 228812
rect 253842 228800 253848 228812
rect 246356 228772 253848 228800
rect 246356 228760 246362 228772
rect 253842 228760 253848 228772
rect 253900 228760 253906 228812
rect 255130 228760 255136 228812
rect 255188 228800 255194 228812
rect 295702 228800 295708 228812
rect 255188 228772 295708 228800
rect 255188 228760 255194 228772
rect 295702 228760 295708 228772
rect 295760 228760 295766 228812
rect 317966 228760 317972 228812
rect 318024 228800 318030 228812
rect 344646 228800 344652 228812
rect 318024 228772 344652 228800
rect 318024 228760 318030 228772
rect 344646 228760 344652 228772
rect 344704 228760 344710 228812
rect 346210 228760 346216 228812
rect 346268 228800 346274 228812
rect 366542 228800 366548 228812
rect 346268 228772 366548 228800
rect 346268 228760 346274 228772
rect 366542 228760 366548 228772
rect 366600 228760 366606 228812
rect 376570 228760 376576 228812
rect 376628 228800 376634 228812
rect 389726 228800 389732 228812
rect 376628 228772 389732 228800
rect 376628 228760 376634 228772
rect 389726 228760 389732 228772
rect 389784 228760 389790 228812
rect 401410 228760 401416 228812
rect 401468 228800 401474 228812
rect 408402 228800 408408 228812
rect 401468 228772 408408 228800
rect 401468 228760 401474 228772
rect 408402 228760 408408 228772
rect 408460 228760 408466 228812
rect 493778 228760 493784 228812
rect 493836 228800 493842 228812
rect 506014 228800 506020 228812
rect 493836 228772 506020 228800
rect 493836 228760 493842 228772
rect 506014 228760 506020 228772
rect 506072 228760 506078 228812
rect 519814 228760 519820 228812
rect 519872 228800 519878 228812
rect 543182 228800 543188 228812
rect 519872 228772 543188 228800
rect 519872 228760 519878 228772
rect 543182 228760 543188 228772
rect 543240 228760 543246 228812
rect 675846 228760 675852 228812
rect 675904 228800 675910 228812
rect 676214 228800 676220 228812
rect 675904 228772 676220 228800
rect 675904 228760 675910 228772
rect 676214 228760 676220 228772
rect 676272 228760 676278 228812
rect 237098 228664 237104 228676
rect 175568 228636 224264 228664
rect 224328 228636 237104 228664
rect 62758 228488 62764 228540
rect 62816 228528 62822 228540
rect 140774 228528 140780 228540
rect 62816 228500 140780 228528
rect 62816 228488 62822 228500
rect 140774 228488 140780 228500
rect 140832 228488 140838 228540
rect 140958 228488 140964 228540
rect 141016 228528 141022 228540
rect 141016 228500 149744 228528
rect 141016 228488 141022 228500
rect 66162 228352 66168 228404
rect 66220 228392 66226 228404
rect 147628 228392 147634 228404
rect 66220 228364 147634 228392
rect 66220 228352 66226 228364
rect 147628 228352 147634 228364
rect 147686 228352 147692 228404
rect 149716 228392 149744 228500
rect 153286 228488 153292 228540
rect 153344 228528 153350 228540
rect 204898 228528 204904 228540
rect 153344 228500 204904 228528
rect 153344 228488 153350 228500
rect 204898 228488 204904 228500
rect 204956 228488 204962 228540
rect 205082 228488 205088 228540
rect 205140 228528 205146 228540
rect 224328 228528 224356 228636
rect 237098 228624 237104 228636
rect 237156 228624 237162 228676
rect 239398 228624 239404 228676
rect 239456 228664 239462 228676
rect 284110 228664 284116 228676
rect 239456 228636 284116 228664
rect 239456 228624 239462 228636
rect 284110 228624 284116 228636
rect 284168 228624 284174 228676
rect 292390 228624 292396 228676
rect 292448 228664 292454 228676
rect 326614 228664 326620 228676
rect 292448 228636 326620 228664
rect 292448 228624 292454 228636
rect 326614 228624 326620 228636
rect 326672 228624 326678 228676
rect 333238 228624 333244 228676
rect 333296 228664 333302 228676
rect 355594 228664 355600 228676
rect 333296 228636 355600 228664
rect 333296 228624 333302 228636
rect 355594 228624 355600 228636
rect 355652 228624 355658 228676
rect 369762 228664 369768 228676
rect 359016 228636 369768 228664
rect 267366 228528 267372 228540
rect 205140 228500 224356 228528
rect 224420 228500 267372 228528
rect 205140 228488 205146 228500
rect 157426 228392 157432 228404
rect 149716 228364 157432 228392
rect 157426 228352 157432 228364
rect 157484 228352 157490 228404
rect 157794 228352 157800 228404
rect 157852 228392 157858 228404
rect 214098 228392 214104 228404
rect 157852 228364 214104 228392
rect 157852 228352 157858 228364
rect 214098 228352 214104 228364
rect 214156 228352 214162 228404
rect 222746 228392 222752 228404
rect 214576 228364 222752 228392
rect 102042 228216 102048 228268
rect 102100 228256 102106 228268
rect 171042 228256 171048 228268
rect 102100 228228 171048 228256
rect 102100 228216 102106 228228
rect 171042 228216 171048 228228
rect 171100 228216 171106 228268
rect 171226 228216 171232 228268
rect 171284 228256 171290 228268
rect 214576 228256 214604 228364
rect 222746 228352 222752 228364
rect 222804 228352 222810 228404
rect 224034 228352 224040 228404
rect 224092 228392 224098 228404
rect 224420 228392 224448 228500
rect 267366 228488 267372 228500
rect 267424 228488 267430 228540
rect 267550 228488 267556 228540
rect 267608 228528 267614 228540
rect 307294 228528 307300 228540
rect 267608 228500 307300 228528
rect 267608 228488 267614 228500
rect 307294 228488 307300 228500
rect 307352 228488 307358 228540
rect 307662 228488 307668 228540
rect 307720 228528 307726 228540
rect 335630 228528 335636 228540
rect 307720 228500 335636 228528
rect 307720 228488 307726 228500
rect 335630 228488 335636 228500
rect 335688 228488 335694 228540
rect 336642 228488 336648 228540
rect 336700 228528 336706 228540
rect 358814 228528 358820 228540
rect 336700 228500 358820 228528
rect 336700 228488 336706 228500
rect 358814 228488 358820 228500
rect 358872 228488 358878 228540
rect 224092 228364 224448 228392
rect 224092 228352 224098 228364
rect 225690 228352 225696 228404
rect 225748 228392 225754 228404
rect 273806 228392 273812 228404
rect 225748 228364 273812 228392
rect 225748 228352 225754 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 284110 228352 284116 228404
rect 284168 228392 284174 228404
rect 320174 228392 320180 228404
rect 284168 228364 320180 228392
rect 284168 228352 284174 228364
rect 320174 228352 320180 228364
rect 320232 228352 320238 228404
rect 326890 228352 326896 228404
rect 326948 228392 326954 228404
rect 351086 228392 351092 228404
rect 326948 228364 351092 228392
rect 326948 228352 326954 228364
rect 351086 228352 351092 228364
rect 351144 228352 351150 228404
rect 355226 228352 355232 228404
rect 355284 228392 355290 228404
rect 359016 228392 359044 228636
rect 369762 228624 369768 228636
rect 369820 228624 369826 228676
rect 373810 228624 373816 228676
rect 373868 228664 373874 228676
rect 387242 228664 387248 228676
rect 373868 228636 387248 228664
rect 373868 228624 373874 228636
rect 387242 228624 387248 228636
rect 387300 228624 387306 228676
rect 390278 228624 390284 228676
rect 390336 228664 390342 228676
rect 400030 228664 400036 228676
rect 390336 228636 400036 228664
rect 390336 228624 390342 228636
rect 400030 228624 400036 228636
rect 400088 228624 400094 228676
rect 410886 228624 410892 228676
rect 410944 228664 410950 228676
rect 416130 228664 416136 228676
rect 410944 228636 416136 228664
rect 410944 228624 410950 228636
rect 416130 228624 416136 228636
rect 416188 228624 416194 228676
rect 478782 228624 478788 228676
rect 478840 228664 478846 228676
rect 483566 228664 483572 228676
rect 478840 228636 483572 228664
rect 478840 228624 478846 228636
rect 483566 228624 483572 228636
rect 483624 228624 483630 228676
rect 495342 228624 495348 228676
rect 495400 228664 495406 228676
rect 511810 228664 511816 228676
rect 495400 228636 511816 228664
rect 495400 228624 495406 228636
rect 511810 228624 511816 228636
rect 511868 228624 511874 228676
rect 512086 228624 512092 228676
rect 512144 228664 512150 228676
rect 512144 228636 528554 228664
rect 512144 228624 512150 228636
rect 366910 228488 366916 228540
rect 366968 228528 366974 228540
rect 381998 228528 382004 228540
rect 366968 228500 382004 228528
rect 366968 228488 366974 228500
rect 381998 228488 382004 228500
rect 382056 228488 382062 228540
rect 392946 228528 392952 228540
rect 383626 228500 392952 228528
rect 355284 228364 359044 228392
rect 355284 228352 355290 228364
rect 362862 228352 362868 228404
rect 362920 228392 362926 228404
rect 379422 228392 379428 228404
rect 362920 228364 379428 228392
rect 362920 228352 362926 228364
rect 379422 228352 379428 228364
rect 379480 228352 379486 228404
rect 381722 228352 381728 228404
rect 381780 228392 381786 228404
rect 383626 228392 383654 228500
rect 392946 228488 392952 228500
rect 393004 228488 393010 228540
rect 393222 228488 393228 228540
rect 393280 228528 393286 228540
rect 393280 228500 397960 228528
rect 393280 228488 393286 228500
rect 381780 228364 383654 228392
rect 381780 228352 381786 228364
rect 391842 228352 391848 228404
rect 391900 228392 391906 228404
rect 397932 228392 397960 228500
rect 400122 228488 400128 228540
rect 400180 228528 400186 228540
rect 407758 228528 407764 228540
rect 400180 228500 407764 228528
rect 400180 228488 400186 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 482462 228488 482468 228540
rect 482520 228528 482526 228540
rect 494606 228528 494612 228540
rect 482520 228500 494612 228528
rect 482520 228488 482526 228500
rect 494606 228488 494612 228500
rect 494664 228488 494670 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 520918 228528 520924 228540
rect 502484 228500 520924 228528
rect 502484 228488 502490 228500
rect 520918 228488 520924 228500
rect 520976 228488 520982 228540
rect 402606 228392 402612 228404
rect 391900 228364 393314 228392
rect 397932 228364 402612 228392
rect 391900 228352 391906 228364
rect 171284 228228 214604 228256
rect 171284 228216 171290 228228
rect 214742 228216 214748 228268
rect 214800 228256 214806 228268
rect 257062 228256 257068 228268
rect 214800 228228 257068 228256
rect 214800 228216 214806 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 277210 228216 277216 228268
rect 277268 228256 277274 228268
rect 311802 228256 311808 228268
rect 277268 228228 311808 228256
rect 277268 228216 277274 228228
rect 311802 228216 311808 228228
rect 311860 228216 311866 228268
rect 393286 228256 393314 228364
rect 402606 228352 402612 228364
rect 402664 228352 402670 228404
rect 409782 228352 409788 228404
rect 409840 228392 409846 228404
rect 415486 228392 415492 228404
rect 409840 228364 415492 228392
rect 409840 228352 409846 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 487614 228352 487620 228404
rect 487672 228392 487678 228404
rect 501506 228392 501512 228404
rect 487672 228364 501512 228392
rect 487672 228352 487678 228364
rect 501506 228352 501512 228364
rect 501564 228352 501570 228404
rect 506290 228352 506296 228404
rect 506348 228392 506354 228404
rect 525886 228392 525892 228404
rect 506348 228364 525892 228392
rect 506348 228352 506354 228364
rect 525886 228352 525892 228364
rect 525944 228352 525950 228404
rect 528526 228392 528554 228636
rect 533982 228624 533988 228676
rect 534040 228664 534046 228676
rect 561582 228664 561588 228676
rect 534040 228636 561588 228664
rect 534040 228624 534046 228636
rect 561582 228624 561588 228636
rect 561640 228624 561646 228676
rect 673388 228540 673440 228546
rect 531406 228488 531412 228540
rect 531464 228528 531470 228540
rect 558178 228528 558184 228540
rect 531464 228500 558184 228528
rect 531464 228488 531470 228500
rect 558178 228488 558184 228500
rect 558236 228488 558242 228540
rect 673388 228482 673440 228488
rect 672166 228420 672172 228472
rect 672224 228460 672230 228472
rect 672224 228432 673302 228460
rect 672224 228420 672230 228432
rect 533890 228392 533896 228404
rect 528526 228364 533896 228392
rect 533890 228352 533896 228364
rect 533948 228352 533954 228404
rect 537846 228352 537852 228404
rect 537904 228392 537910 228404
rect 566366 228392 566372 228404
rect 537904 228364 566372 228392
rect 537904 228352 537910 228364
rect 566366 228352 566372 228364
rect 566424 228352 566430 228404
rect 403894 228256 403900 228268
rect 393286 228228 403900 228256
rect 403894 228216 403900 228228
rect 403952 228216 403958 228268
rect 479702 228216 479708 228268
rect 479760 228256 479766 228268
rect 487798 228256 487804 228268
rect 479760 228228 487804 228256
rect 479760 228216 479766 228228
rect 487798 228216 487804 228228
rect 487856 228216 487862 228268
rect 671798 228216 671804 228268
rect 671856 228256 671862 228268
rect 671856 228228 673190 228256
rect 671856 228216 671862 228228
rect 112990 228080 112996 228132
rect 113048 228120 113054 228132
rect 115750 228120 115756 228132
rect 113048 228092 115756 228120
rect 113048 228080 113054 228092
rect 115750 228080 115756 228092
rect 115808 228080 115814 228132
rect 140958 228120 140964 228132
rect 115952 228092 140964 228120
rect 115566 227944 115572 227996
rect 115624 227984 115630 227996
rect 115952 227984 115980 228092
rect 140958 228080 140964 228092
rect 141016 228080 141022 228132
rect 141142 228080 141148 228132
rect 141200 228120 141206 228132
rect 201034 228120 201040 228132
rect 141200 228092 201040 228120
rect 141200 228080 141206 228092
rect 201034 228080 201040 228092
rect 201092 228080 201098 228132
rect 201402 228080 201408 228132
rect 201460 228120 201466 228132
rect 252554 228120 252560 228132
rect 201460 228092 252560 228120
rect 201460 228080 201466 228092
rect 252554 228080 252560 228092
rect 252612 228080 252618 228132
rect 288158 228080 288164 228132
rect 288216 228120 288222 228132
rect 321462 228120 321468 228132
rect 288216 228092 321468 228120
rect 288216 228080 288222 228092
rect 321462 228080 321468 228092
rect 321520 228080 321526 228132
rect 484026 228080 484032 228132
rect 484084 228120 484090 228132
rect 490558 228120 490564 228132
rect 484084 228092 490564 228120
rect 484084 228080 484090 228092
rect 490558 228080 490564 228092
rect 490616 228080 490622 228132
rect 115624 227956 115980 227984
rect 115624 227944 115630 227956
rect 122742 227944 122748 227996
rect 122800 227984 122806 227996
rect 192662 227984 192668 227996
rect 122800 227956 192668 227984
rect 122800 227944 122806 227956
rect 192662 227944 192668 227956
rect 192720 227944 192726 227996
rect 197906 227944 197912 227996
rect 197964 227984 197970 227996
rect 204530 227984 204536 227996
rect 197964 227956 204536 227984
rect 197964 227944 197970 227956
rect 204530 227944 204536 227956
rect 204588 227944 204594 227996
rect 205450 227944 205456 227996
rect 205508 227984 205514 227996
rect 214742 227984 214748 227996
rect 205508 227956 214748 227984
rect 205508 227944 205514 227956
rect 214742 227944 214748 227956
rect 214800 227944 214806 227996
rect 222746 227944 222752 227996
rect 222804 227984 222810 227996
rect 226150 227984 226156 227996
rect 222804 227956 226156 227984
rect 222804 227944 222810 227956
rect 226150 227944 226156 227956
rect 226208 227944 226214 227996
rect 272518 227984 272524 227996
rect 229066 227956 272524 227984
rect 134610 227808 134616 227860
rect 134668 227848 134674 227860
rect 141142 227848 141148 227860
rect 134668 227820 141148 227848
rect 134668 227808 134674 227820
rect 141142 227808 141148 227820
rect 141200 227808 141206 227860
rect 141326 227808 141332 227860
rect 141384 227848 141390 227860
rect 200390 227848 200396 227860
rect 141384 227820 200396 227848
rect 141384 227808 141390 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 226150 227808 226156 227860
rect 226208 227848 226214 227860
rect 229066 227848 229094 227956
rect 272518 227944 272524 227956
rect 272576 227944 272582 227996
rect 673046 227928 673098 227934
rect 369118 227876 369124 227928
rect 369176 227916 369182 227928
rect 375558 227916 375564 227928
rect 369176 227888 375564 227916
rect 369176 227876 369182 227888
rect 375558 227876 375564 227888
rect 375616 227876 375622 227928
rect 407758 227876 407764 227928
rect 407816 227916 407822 227928
rect 411622 227916 411628 227928
rect 407816 227888 411628 227916
rect 407816 227876 407822 227888
rect 411622 227876 411628 227888
rect 411680 227876 411686 227928
rect 471514 227876 471520 227928
rect 471572 227916 471578 227928
rect 479334 227916 479340 227928
rect 471572 227888 479340 227916
rect 471572 227876 471578 227888
rect 479334 227876 479340 227888
rect 479392 227876 479398 227928
rect 673046 227870 673098 227876
rect 226208 227820 229094 227848
rect 226208 227808 226214 227820
rect 242710 227740 242716 227792
rect 242768 227780 242774 227792
rect 245654 227780 245660 227792
rect 242768 227752 245660 227780
rect 242768 227740 242774 227752
rect 245654 227740 245660 227752
rect 245712 227740 245718 227792
rect 255958 227740 255964 227792
rect 256016 227780 256022 227792
rect 258994 227780 259000 227792
rect 256016 227752 259000 227780
rect 256016 227740 256022 227752
rect 258994 227740 259000 227752
rect 259052 227740 259058 227792
rect 366358 227740 366364 227792
rect 366416 227780 366422 227792
rect 372982 227780 372988 227792
rect 366416 227752 372988 227780
rect 366416 227740 366422 227752
rect 372982 227740 372988 227752
rect 373040 227740 373046 227792
rect 393958 227740 393964 227792
rect 394016 227780 394022 227792
rect 395522 227780 395528 227792
rect 394016 227752 395528 227780
rect 394016 227740 394022 227752
rect 395522 227740 395528 227752
rect 395580 227740 395586 227792
rect 396626 227740 396632 227792
rect 396684 227780 396690 227792
rect 397454 227780 397460 227792
rect 396684 227752 397460 227780
rect 396684 227740 396690 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 402238 227740 402244 227792
rect 402296 227780 402302 227792
rect 403250 227780 403256 227792
rect 402296 227752 403256 227780
rect 402296 227740 402302 227752
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 404078 227740 404084 227792
rect 404136 227780 404142 227792
rect 408862 227780 408868 227792
rect 404136 227752 408868 227780
rect 404136 227740 404142 227752
rect 408862 227740 408868 227752
rect 408920 227740 408926 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416682 227740 416688 227792
rect 416740 227780 416746 227792
rect 420638 227780 420644 227792
rect 416740 227752 420644 227780
rect 416740 227740 416746 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 475010 227740 475016 227792
rect 475068 227780 475074 227792
rect 482922 227780 482928 227792
rect 475068 227752 482928 227780
rect 475068 227740 475074 227752
rect 482922 227740 482928 227752
rect 482980 227740 482986 227792
rect 672954 227724 673006 227730
rect 110138 227672 110144 227724
rect 110196 227712 110202 227724
rect 182358 227712 182364 227724
rect 110196 227684 182364 227712
rect 110196 227672 110202 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 186682 227672 186688 227724
rect 186740 227712 186746 227724
rect 187234 227712 187240 227724
rect 186740 227684 187240 227712
rect 186740 227672 186746 227684
rect 187234 227672 187240 227684
rect 187292 227672 187298 227724
rect 191558 227672 191564 227724
rect 191616 227712 191622 227724
rect 191616 227684 238754 227712
rect 191616 227672 191622 227684
rect 238726 227644 238754 227684
rect 270126 227672 270132 227724
rect 270184 227712 270190 227724
rect 306650 227712 306656 227724
rect 270184 227684 306656 227712
rect 270184 227672 270190 227684
rect 306650 227672 306656 227684
rect 306708 227672 306714 227724
rect 321370 227672 321376 227724
rect 321428 227712 321434 227724
rect 346578 227712 346584 227724
rect 321428 227684 346584 227712
rect 321428 227672 321434 227684
rect 346578 227672 346584 227684
rect 346636 227672 346642 227724
rect 525518 227672 525524 227724
rect 525576 227712 525582 227724
rect 537570 227712 537576 227724
rect 525576 227684 537576 227712
rect 525576 227672 525582 227684
rect 537570 227672 537576 227684
rect 537628 227672 537634 227724
rect 672954 227666 673006 227672
rect 248046 227644 248052 227656
rect 238726 227616 248052 227644
rect 248046 227604 248052 227616
rect 248104 227604 248110 227656
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 100662 227536 100668 227588
rect 100720 227576 100726 227588
rect 174630 227576 174636 227588
rect 100720 227548 174636 227576
rect 100720 227536 100726 227548
rect 174630 227536 174636 227548
rect 174688 227536 174694 227588
rect 179046 227536 179052 227588
rect 179104 227576 179110 227588
rect 236454 227576 236460 227588
rect 179104 227548 236460 227576
rect 179104 227536 179110 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 252462 227536 252468 227588
rect 252520 227576 252526 227588
rect 293126 227576 293132 227588
rect 252520 227548 293132 227576
rect 252520 227536 252526 227548
rect 293126 227536 293132 227548
rect 293184 227536 293190 227588
rect 299290 227536 299296 227588
rect 299348 227576 299354 227588
rect 328546 227576 328552 227588
rect 299348 227548 328552 227576
rect 299348 227536 299354 227548
rect 328546 227536 328552 227548
rect 328604 227536 328610 227588
rect 359366 227536 359372 227588
rect 359424 227576 359430 227588
rect 374914 227576 374920 227588
rect 359424 227548 374920 227576
rect 359424 227536 359430 227548
rect 374914 227536 374920 227548
rect 374972 227536 374978 227588
rect 515858 227536 515864 227588
rect 515916 227576 515922 227588
rect 538858 227576 538864 227588
rect 515916 227548 538864 227576
rect 515916 227536 515922 227548
rect 538858 227536 538864 227548
rect 538916 227536 538922 227588
rect 663702 227536 663708 227588
rect 663760 227576 663766 227588
rect 665542 227576 665548 227588
rect 663760 227548 665548 227576
rect 663760 227536 663766 227548
rect 665542 227536 665548 227548
rect 665600 227536 665606 227588
rect 672816 227520 672868 227526
rect 672816 227462 672868 227468
rect 89622 227400 89628 227452
rect 89680 227440 89686 227452
rect 159634 227440 159640 227452
rect 89680 227412 159640 227440
rect 89680 227400 89686 227412
rect 159634 227400 159640 227412
rect 159692 227400 159698 227452
rect 160002 227400 160008 227452
rect 160060 227440 160066 227452
rect 166902 227440 166908 227452
rect 160060 227412 166908 227440
rect 160060 227400 160066 227412
rect 166902 227400 166908 227412
rect 166960 227400 166966 227452
rect 171106 227412 173756 227440
rect 86862 227264 86868 227316
rect 86920 227304 86926 227316
rect 151906 227304 151912 227316
rect 86920 227276 151912 227304
rect 86920 227264 86926 227276
rect 151906 227264 151912 227276
rect 151964 227264 151970 227316
rect 152918 227264 152924 227316
rect 152976 227304 152982 227316
rect 164326 227304 164332 227316
rect 152976 227276 164332 227304
rect 152976 227264 152982 227276
rect 164326 227264 164332 227276
rect 164384 227264 164390 227316
rect 165430 227264 165436 227316
rect 165488 227304 165494 227316
rect 171106 227304 171134 227412
rect 165488 227276 171134 227304
rect 173728 227304 173756 227412
rect 175182 227400 175188 227452
rect 175240 227440 175246 227452
rect 231946 227440 231952 227452
rect 175240 227412 231952 227440
rect 175240 227400 175246 227412
rect 231946 227400 231952 227412
rect 232004 227400 232010 227452
rect 248230 227400 248236 227452
rect 248288 227440 248294 227452
rect 291838 227440 291844 227452
rect 248288 227412 291844 227440
rect 248288 227400 248294 227412
rect 291838 227400 291844 227412
rect 291896 227400 291902 227452
rect 293770 227400 293776 227452
rect 293828 227440 293834 227452
rect 325326 227440 325332 227452
rect 293828 227412 325332 227440
rect 293828 227400 293834 227412
rect 325326 227400 325332 227412
rect 325384 227400 325390 227452
rect 340598 227400 340604 227452
rect 340656 227440 340662 227452
rect 361390 227440 361396 227452
rect 340656 227412 361396 227440
rect 340656 227400 340662 227412
rect 361390 227400 361396 227412
rect 361448 227400 361454 227452
rect 377214 227440 377220 227452
rect 361592 227412 377220 227440
rect 227438 227304 227444 227316
rect 173728 227276 227444 227304
rect 165488 227264 165494 227276
rect 227438 227264 227444 227276
rect 227496 227264 227502 227316
rect 233234 227304 233240 227316
rect 228928 227276 233240 227304
rect 75822 227128 75828 227180
rect 75880 227168 75886 227180
rect 150158 227168 150164 227180
rect 75880 227140 150164 227168
rect 75880 227128 75886 227140
rect 150158 227128 150164 227140
rect 150216 227128 150222 227180
rect 150342 227128 150348 227180
rect 150400 227168 150406 227180
rect 150400 227140 152136 227168
rect 150400 227128 150406 227140
rect 57882 226992 57888 227044
rect 57940 227032 57946 227044
rect 135254 227032 135260 227044
rect 57940 227004 135260 227032
rect 57940 226992 57946 227004
rect 135254 226992 135260 227004
rect 135312 226992 135318 227044
rect 135438 226992 135444 227044
rect 135496 227032 135502 227044
rect 151906 227032 151912 227044
rect 135496 227004 151912 227032
rect 135496 226992 135502 227004
rect 151906 226992 151912 227004
rect 151964 226992 151970 227044
rect 152108 227032 152136 227140
rect 152274 227128 152280 227180
rect 152332 227168 152338 227180
rect 168834 227168 168840 227180
rect 152332 227140 168840 227168
rect 152332 227128 152338 227140
rect 168834 227128 168840 227140
rect 168892 227128 168898 227180
rect 169570 227128 169576 227180
rect 169628 227168 169634 227180
rect 228726 227168 228732 227180
rect 169628 227140 228732 227168
rect 169628 227128 169634 227140
rect 228726 227128 228732 227140
rect 228784 227128 228790 227180
rect 213270 227032 213276 227044
rect 152108 227004 213276 227032
rect 213270 226992 213276 227004
rect 213328 226992 213334 227044
rect 226886 226992 226892 227044
rect 226944 227032 226950 227044
rect 228928 227032 228956 227276
rect 233234 227264 233240 227276
rect 233292 227264 233298 227316
rect 234522 227264 234528 227316
rect 234580 227304 234586 227316
rect 278314 227304 278320 227316
rect 234580 227276 278320 227304
rect 234580 227264 234586 227276
rect 278314 227264 278320 227276
rect 278372 227264 278378 227316
rect 280706 227264 280712 227316
rect 280764 227304 280770 227316
rect 312078 227304 312084 227316
rect 280764 227276 312084 227304
rect 280764 227264 280770 227276
rect 312078 227264 312084 227276
rect 312136 227264 312142 227316
rect 326338 227264 326344 227316
rect 326396 227304 326402 227316
rect 352374 227304 352380 227316
rect 326396 227276 352380 227304
rect 326396 227264 326402 227276
rect 352374 227264 352380 227276
rect 352432 227264 352438 227316
rect 361206 227264 361212 227316
rect 361264 227304 361270 227316
rect 361592 227304 361620 227412
rect 377214 227400 377220 227412
rect 377272 227400 377278 227452
rect 383286 227440 383292 227452
rect 378612 227412 383292 227440
rect 361264 227276 361620 227304
rect 361264 227264 361270 227276
rect 361758 227264 361764 227316
rect 361816 227304 361822 227316
rect 372338 227304 372344 227316
rect 361816 227276 372344 227304
rect 361816 227264 361822 227276
rect 372338 227264 372344 227276
rect 372396 227264 372402 227316
rect 373258 227264 373264 227316
rect 373316 227304 373322 227316
rect 378612 227304 378640 227412
rect 383286 227400 383292 227412
rect 383344 227400 383350 227452
rect 524322 227400 524328 227452
rect 524380 227440 524386 227452
rect 547874 227440 547880 227452
rect 524380 227412 547880 227440
rect 524380 227400 524386 227412
rect 547874 227400 547880 227412
rect 547932 227400 547938 227452
rect 672724 227316 672776 227322
rect 373316 227276 378640 227304
rect 373316 227264 373322 227276
rect 382918 227264 382924 227316
rect 382976 227304 382982 227316
rect 391658 227304 391664 227316
rect 382976 227276 391664 227304
rect 382976 227264 382982 227276
rect 391658 227264 391664 227276
rect 391716 227264 391722 227316
rect 395982 227264 395988 227316
rect 396040 227304 396046 227316
rect 406470 227304 406476 227316
rect 396040 227276 406476 227304
rect 396040 227264 396046 227276
rect 406470 227264 406476 227276
rect 406528 227264 406534 227316
rect 485038 227264 485044 227316
rect 485096 227304 485102 227316
rect 498746 227304 498752 227316
rect 485096 227276 498752 227304
rect 485096 227264 485102 227276
rect 498746 227264 498752 227276
rect 498804 227264 498810 227316
rect 501322 227264 501328 227316
rect 501380 227304 501386 227316
rect 517698 227304 517704 227316
rect 501380 227276 517704 227304
rect 501380 227264 501386 227276
rect 517698 227264 517704 227276
rect 517756 227264 517762 227316
rect 521746 227264 521752 227316
rect 521804 227304 521810 227316
rect 545758 227304 545764 227316
rect 521804 227276 545764 227304
rect 521804 227264 521810 227276
rect 545758 227264 545764 227276
rect 545816 227264 545822 227316
rect 672724 227258 672776 227264
rect 672258 227196 672264 227248
rect 672316 227236 672322 227248
rect 672316 227208 672630 227236
rect 672316 227196 672322 227208
rect 235902 227128 235908 227180
rect 235960 227168 235966 227180
rect 280246 227168 280252 227180
rect 235960 227140 280252 227168
rect 235960 227128 235966 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 296438 227128 296444 227180
rect 296496 227168 296502 227180
rect 329190 227168 329196 227180
rect 296496 227140 329196 227168
rect 296496 227128 296502 227140
rect 329190 227128 329196 227140
rect 329248 227128 329254 227180
rect 329742 227128 329748 227180
rect 329800 227168 329806 227180
rect 353662 227168 353668 227180
rect 329800 227140 353668 227168
rect 329800 227128 329806 227140
rect 353662 227128 353668 227140
rect 353720 227128 353726 227180
rect 354582 227128 354588 227180
rect 354640 227168 354646 227180
rect 373626 227168 373632 227180
rect 354640 227140 373632 227168
rect 354640 227128 354646 227140
rect 373626 227128 373632 227140
rect 373684 227128 373690 227180
rect 381906 227128 381912 227180
rect 381964 227168 381970 227180
rect 396166 227168 396172 227180
rect 381964 227140 396172 227168
rect 381964 227128 381970 227140
rect 396166 227128 396172 227140
rect 396224 227128 396230 227180
rect 481174 227128 481180 227180
rect 481232 227168 481238 227180
rect 492950 227168 492956 227180
rect 481232 227140 492956 227168
rect 481232 227128 481238 227140
rect 492950 227128 492956 227140
rect 493008 227128 493014 227180
rect 498562 227128 498568 227180
rect 498620 227168 498626 227180
rect 515858 227168 515864 227180
rect 498620 227140 515864 227168
rect 498620 227128 498626 227140
rect 515858 227128 515864 227140
rect 515916 227128 515922 227180
rect 516042 227128 516048 227180
rect 516100 227168 516106 227180
rect 525058 227168 525064 227180
rect 516100 227140 525064 227168
rect 516100 227128 516106 227140
rect 525058 227128 525064 227140
rect 525116 227128 525122 227180
rect 535914 227128 535920 227180
rect 535972 227168 535978 227180
rect 564066 227168 564072 227180
rect 535972 227140 564072 227168
rect 535972 227128 535978 227140
rect 564066 227128 564072 227140
rect 564124 227128 564130 227180
rect 226944 227004 228956 227032
rect 226944 226992 226950 227004
rect 229048 226992 229054 227044
rect 229106 227032 229112 227044
rect 271230 227032 271236 227044
rect 229106 227004 271236 227032
rect 229106 226992 229112 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 308766 226992 308772 227044
rect 308824 227032 308830 227044
rect 336274 227032 336280 227044
rect 308824 227004 336280 227032
rect 308824 226992 308830 227004
rect 336274 226992 336280 227004
rect 336332 226992 336338 227044
rect 336458 226992 336464 227044
rect 336516 227032 336522 227044
rect 360102 227032 360108 227044
rect 336516 227004 360108 227032
rect 336516 226992 336522 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 369762 226992 369768 227044
rect 369820 227032 369826 227044
rect 385862 227032 385868 227044
rect 369820 227004 385868 227032
rect 369820 226992 369826 227004
rect 385862 226992 385868 227004
rect 385920 226992 385926 227044
rect 386322 226992 386328 227044
rect 386380 227032 386386 227044
rect 398742 227032 398748 227044
rect 386380 227004 398748 227032
rect 386380 226992 386386 227004
rect 398742 226992 398748 227004
rect 398800 226992 398806 227044
rect 472158 226992 472164 227044
rect 472216 227032 472222 227044
rect 481174 227032 481180 227044
rect 472216 227004 481180 227032
rect 472216 226992 472222 227004
rect 481174 226992 481180 227004
rect 481232 226992 481238 227044
rect 497274 226992 497280 227044
rect 497332 227032 497338 227044
rect 497332 227004 509234 227032
rect 497332 226992 497338 227004
rect 106918 226856 106924 226908
rect 106976 226896 106982 226908
rect 125778 226896 125784 226908
rect 106976 226868 125784 226896
rect 106976 226856 106982 226868
rect 125778 226856 125784 226868
rect 125836 226856 125842 226908
rect 190730 226896 190736 226908
rect 125980 226868 190736 226896
rect 121086 226720 121092 226772
rect 121144 226760 121150 226772
rect 125980 226760 126008 226868
rect 190730 226856 190736 226868
rect 190788 226856 190794 226908
rect 200022 226856 200028 226908
rect 200080 226896 200086 226908
rect 251910 226896 251916 226908
rect 200080 226868 251916 226896
rect 200080 226856 200086 226868
rect 251910 226856 251916 226868
rect 251968 226856 251974 226908
rect 272426 226856 272432 226908
rect 272484 226896 272490 226908
rect 284754 226896 284760 226908
rect 272484 226868 284760 226896
rect 272484 226856 272490 226868
rect 284754 226856 284760 226868
rect 284812 226856 284818 226908
rect 355502 226856 355508 226908
rect 355560 226896 355566 226908
rect 361758 226896 361764 226908
rect 355560 226868 361764 226896
rect 355560 226856 355566 226868
rect 361758 226856 361764 226868
rect 361816 226856 361822 226908
rect 398466 226856 398472 226908
rect 398524 226896 398530 226908
rect 408678 226896 408684 226908
rect 398524 226868 408684 226896
rect 398524 226856 398530 226868
rect 408678 226856 408684 226868
rect 408736 226856 408742 226908
rect 509206 226896 509234 227004
rect 514018 226992 514024 227044
rect 514076 227032 514082 227044
rect 536006 227032 536012 227044
rect 514076 227004 536012 227032
rect 514076 226992 514082 227004
rect 536006 226992 536012 227004
rect 536064 226992 536070 227044
rect 537202 226992 537208 227044
rect 537260 227032 537266 227044
rect 565722 227032 565728 227044
rect 537260 227004 565728 227032
rect 537260 226992 537266 227004
rect 565722 226992 565728 227004
rect 565780 226992 565786 227044
rect 671062 226992 671068 227044
rect 671120 227032 671126 227044
rect 671120 227004 672520 227032
rect 671120 226992 671126 227004
rect 514294 226896 514300 226908
rect 509206 226868 514300 226896
rect 514294 226856 514300 226868
rect 514352 226856 514358 226908
rect 672258 226856 672264 226908
rect 672316 226896 672322 226908
rect 672316 226868 672406 226896
rect 672316 226856 672322 226868
rect 189718 226760 189724 226772
rect 121144 226732 126008 226760
rect 126072 226732 189724 226760
rect 121144 226720 121150 226732
rect 119982 226584 119988 226636
rect 120040 226624 120046 226636
rect 126072 226624 126100 226732
rect 189718 226720 189724 226732
rect 189776 226720 189782 226772
rect 195882 226720 195888 226772
rect 195940 226760 195946 226772
rect 199286 226760 199292 226772
rect 195940 226732 199292 226760
rect 195940 226720 195946 226732
rect 199286 226720 199292 226732
rect 199344 226720 199350 226772
rect 212166 226720 212172 226772
rect 212224 226760 212230 226772
rect 262214 226760 262220 226772
rect 212224 226732 262220 226760
rect 212224 226720 212230 226732
rect 262214 226720 262220 226732
rect 262272 226720 262278 226772
rect 135438 226624 135444 226636
rect 120040 226596 126100 226624
rect 126164 226596 135444 226624
rect 120040 226584 120046 226596
rect 125778 226448 125784 226500
rect 125836 226488 125842 226500
rect 126164 226488 126192 226596
rect 135438 226584 135444 226596
rect 135496 226584 135502 226636
rect 135622 226584 135628 226636
rect 135680 226624 135686 226636
rect 135680 226596 137416 226624
rect 135680 226584 135686 226596
rect 125836 226460 126192 226488
rect 125836 226448 125842 226460
rect 129366 226448 129372 226500
rect 129424 226488 129430 226500
rect 137186 226488 137192 226500
rect 129424 226460 137192 226488
rect 129424 226448 129430 226460
rect 137186 226448 137192 226460
rect 137244 226448 137250 226500
rect 137388 226488 137416 226596
rect 137554 226584 137560 226636
rect 137612 226624 137618 226636
rect 197354 226624 197360 226636
rect 137612 226596 197360 226624
rect 137612 226584 137618 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 222010 226584 222016 226636
rect 222068 226624 222074 226636
rect 269942 226624 269948 226636
rect 222068 226596 269948 226624
rect 222068 226584 222074 226596
rect 269942 226584 269948 226596
rect 270000 226584 270006 226636
rect 669406 226584 669412 226636
rect 669464 226624 669470 226636
rect 669464 226596 672290 226624
rect 669464 226584 669470 226596
rect 142108 226488 142114 226500
rect 137388 226460 142114 226488
rect 142108 226448 142114 226460
rect 142166 226448 142172 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 205266 226488 205272 226500
rect 142304 226460 205272 226488
rect 142304 226448 142310 226460
rect 205266 226448 205272 226460
rect 205324 226448 205330 226500
rect 213178 226448 213184 226500
rect 213236 226488 213242 226500
rect 217778 226488 217784 226500
rect 213236 226460 217784 226488
rect 213236 226448 213242 226460
rect 217778 226448 217784 226460
rect 217836 226448 217842 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 229002 226488 229008 226500
rect 221884 226460 229008 226488
rect 221884 226448 221890 226460
rect 229002 226448 229008 226460
rect 229060 226448 229066 226500
rect 232498 226448 232504 226500
rect 232556 226488 232562 226500
rect 266722 226488 266728 226500
rect 232556 226460 266728 226488
rect 232556 226448 232562 226460
rect 266722 226448 266728 226460
rect 266780 226448 266786 226500
rect 666830 226448 666836 226500
rect 666888 226488 666894 226500
rect 666888 226460 672182 226488
rect 666888 226448 666894 226460
rect 291838 226380 291844 226432
rect 291896 226420 291902 226432
rect 295058 226420 295064 226432
rect 291896 226392 295064 226420
rect 291896 226380 291902 226392
rect 295058 226380 295064 226392
rect 295116 226380 295122 226432
rect 152200 226324 152688 226352
rect 83458 226244 83464 226296
rect 83516 226284 83522 226296
rect 152200 226284 152228 226324
rect 83516 226256 152228 226284
rect 83516 226244 83522 226256
rect 69566 226108 69572 226160
rect 69624 226148 69630 226160
rect 143534 226148 143540 226160
rect 69624 226120 143540 226148
rect 69624 226108 69630 226120
rect 143534 226108 143540 226120
rect 143592 226108 143598 226160
rect 152660 226148 152688 226324
rect 166948 226312 166954 226364
rect 167006 226352 167012 226364
rect 220998 226352 221004 226364
rect 167006 226324 221004 226352
rect 167006 226312 167012 226324
rect 220998 226312 221004 226324
rect 221056 226312 221062 226364
rect 152826 226244 152832 226296
rect 152884 226284 152890 226296
rect 161934 226284 161940 226296
rect 152884 226256 161940 226284
rect 152884 226244 152890 226256
rect 161934 226244 161940 226256
rect 161992 226244 161998 226296
rect 162302 226244 162308 226296
rect 162360 226284 162366 226296
rect 166810 226284 166816 226296
rect 162360 226256 166816 226284
rect 162360 226244 162366 226256
rect 166810 226244 166816 226256
rect 166868 226244 166874 226296
rect 222470 226244 222476 226296
rect 222528 226284 222534 226296
rect 225506 226284 225512 226296
rect 222528 226256 225512 226284
rect 222528 226244 222534 226256
rect 225506 226244 225512 226256
rect 225564 226244 225570 226296
rect 228726 226244 228732 226296
rect 228784 226284 228790 226296
rect 275094 226284 275100 226296
rect 228784 226256 275100 226284
rect 228784 226244 228790 226256
rect 275094 226244 275100 226256
rect 275152 226244 275158 226296
rect 278498 226244 278504 226296
rect 278556 226284 278562 226296
rect 315022 226284 315028 226296
rect 278556 226256 315028 226284
rect 278556 226244 278562 226256
rect 315022 226244 315028 226256
rect 315080 226244 315086 226296
rect 317322 226244 317328 226296
rect 317380 226284 317386 226296
rect 334250 226284 334256 226296
rect 317380 226256 334256 226284
rect 317380 226244 317386 226256
rect 334250 226244 334256 226256
rect 334308 226244 334314 226296
rect 503254 226244 503260 226296
rect 503312 226284 503318 226296
rect 510154 226284 510160 226296
rect 503312 226256 510160 226284
rect 503312 226244 503318 226256
rect 510154 226244 510160 226256
rect 510212 226244 510218 226296
rect 529934 226244 529940 226296
rect 529992 226284 529998 226296
rect 544930 226284 544936 226296
rect 529992 226256 544936 226284
rect 529992 226244 529998 226256
rect 544930 226244 544936 226256
rect 544988 226244 544994 226296
rect 562318 226244 562324 226296
rect 562376 226284 562382 226296
rect 568390 226284 568396 226296
rect 562376 226256 568396 226284
rect 562376 226244 562382 226256
rect 568390 226244 568396 226256
rect 568448 226244 568454 226296
rect 671062 226244 671068 226296
rect 671120 226284 671126 226296
rect 671120 226256 672060 226284
rect 671120 226244 671126 226256
rect 157426 226148 157432 226160
rect 152660 226120 157432 226148
rect 157426 226108 157432 226120
rect 157484 226108 157490 226160
rect 157610 226108 157616 226160
rect 157668 226148 157674 226160
rect 215846 226148 215852 226160
rect 157668 226120 215852 226148
rect 157668 226108 157674 226120
rect 215846 226108 215852 226120
rect 215904 226108 215910 226160
rect 216490 226108 216496 226160
rect 216548 226148 216554 226160
rect 264790 226148 264796 226160
rect 216548 226120 264796 226148
rect 216548 226108 216554 226120
rect 264790 226108 264796 226120
rect 264848 226108 264854 226160
rect 266262 226108 266268 226160
rect 266320 226148 266326 226160
rect 303430 226148 303436 226160
rect 266320 226120 303436 226148
rect 266320 226108 266326 226120
rect 303430 226108 303436 226120
rect 303488 226108 303494 226160
rect 325418 226108 325424 226160
rect 325476 226148 325482 226160
rect 349154 226148 349160 226160
rect 325476 226120 349160 226148
rect 325476 226108 325482 226120
rect 349154 226108 349160 226120
rect 349212 226108 349218 226160
rect 510798 226108 510804 226160
rect 510856 226148 510862 226160
rect 531682 226148 531688 226160
rect 510856 226120 531688 226148
rect 510856 226108 510862 226120
rect 531682 226108 531688 226120
rect 531740 226108 531746 226160
rect 667014 226040 667020 226092
rect 667072 226080 667078 226092
rect 667072 226052 671968 226080
rect 667072 226040 667078 226052
rect 93762 225972 93768 226024
rect 93820 226012 93826 226024
rect 161566 226012 161572 226024
rect 93820 225984 161572 226012
rect 93820 225972 93826 225984
rect 161566 225972 161572 225984
rect 161624 225972 161630 226024
rect 161934 225972 161940 226024
rect 161992 226012 161998 226024
rect 171042 226012 171048 226024
rect 161992 225984 171048 226012
rect 161992 225972 161998 225984
rect 171042 225972 171048 225984
rect 171100 225972 171106 226024
rect 171226 225972 171232 226024
rect 171284 226012 171290 226024
rect 186268 226012 186274 226024
rect 171284 225984 186274 226012
rect 171284 225972 171290 225984
rect 186268 225972 186274 225984
rect 186326 225972 186332 226024
rect 186406 225972 186412 226024
rect 186464 226012 186470 226024
rect 224218 226012 224224 226024
rect 186464 225984 224224 226012
rect 186464 225972 186470 225984
rect 224218 225972 224224 225984
rect 224276 225972 224282 226024
rect 233878 226012 233884 226024
rect 229066 225984 233884 226012
rect 95142 225836 95148 225888
rect 95200 225876 95206 225888
rect 166810 225876 166816 225888
rect 95200 225848 166816 225876
rect 95200 225836 95206 225848
rect 166810 225836 166816 225848
rect 166868 225836 166874 225888
rect 166948 225836 166954 225888
rect 167006 225876 167012 225888
rect 167006 225848 176148 225876
rect 167006 225836 167012 225848
rect 64782 225700 64788 225752
rect 64840 225740 64846 225752
rect 92474 225740 92480 225752
rect 64840 225712 92480 225740
rect 64840 225700 64846 225712
rect 92474 225700 92480 225712
rect 92532 225700 92538 225752
rect 108298 225700 108304 225752
rect 108356 225740 108362 225752
rect 171042 225740 171048 225752
rect 108356 225712 171048 225740
rect 108356 225700 108362 225712
rect 171042 225700 171048 225712
rect 171100 225700 171106 225752
rect 171226 225700 171232 225752
rect 171284 225740 171290 225752
rect 175918 225740 175924 225752
rect 171284 225712 175924 225740
rect 171284 225700 171290 225712
rect 175918 225700 175924 225712
rect 175976 225700 175982 225752
rect 176120 225740 176148 225848
rect 176286 225836 176292 225888
rect 176344 225876 176350 225888
rect 176608 225876 176614 225888
rect 176344 225848 176614 225876
rect 176344 225836 176350 225848
rect 176608 225836 176614 225848
rect 176666 225836 176672 225888
rect 176746 225836 176752 225888
rect 176804 225876 176810 225888
rect 181070 225876 181076 225888
rect 176804 225848 181076 225876
rect 176804 225836 176810 225848
rect 181070 225836 181076 225848
rect 181128 225836 181134 225888
rect 185946 225876 185952 225888
rect 181272 225848 185952 225876
rect 181272 225740 181300 225848
rect 185946 225836 185952 225848
rect 186004 225836 186010 225888
rect 186130 225836 186136 225888
rect 186188 225876 186194 225888
rect 229066 225876 229094 225984
rect 233878 225972 233884 225984
rect 233936 225972 233942 226024
rect 243446 225972 243452 226024
rect 243504 226012 243510 226024
rect 248690 226012 248696 226024
rect 243504 225984 248696 226012
rect 243504 225972 243510 225984
rect 248690 225972 248696 225984
rect 248748 225972 248754 226024
rect 267688 225972 267694 226024
rect 267746 226012 267752 226024
rect 304074 226012 304080 226024
rect 267746 225984 304080 226012
rect 267746 225972 267752 225984
rect 304074 225972 304080 225984
rect 304132 225972 304138 226024
rect 313090 225972 313096 226024
rect 313148 226012 313154 226024
rect 340782 226012 340788 226024
rect 313148 225984 340788 226012
rect 313148 225972 313154 225984
rect 340782 225972 340788 225984
rect 340840 225972 340846 226024
rect 347866 226012 347872 226024
rect 344986 225984 347872 226012
rect 239030 225876 239036 225888
rect 186188 225848 229094 225876
rect 232700 225848 239036 225876
rect 186188 225836 186194 225848
rect 176120 225712 181300 225740
rect 181438 225700 181444 225752
rect 181496 225740 181502 225752
rect 186682 225740 186688 225752
rect 181496 225712 186688 225740
rect 181496 225700 181502 225712
rect 186682 225700 186688 225712
rect 186740 225700 186746 225752
rect 186866 225700 186872 225752
rect 186924 225740 186930 225752
rect 232700 225740 232728 225848
rect 239030 225836 239036 225848
rect 239088 225836 239094 225888
rect 249702 225836 249708 225888
rect 249760 225876 249766 225888
rect 290550 225876 290556 225888
rect 249760 225848 290556 225876
rect 249760 225836 249766 225848
rect 290550 225836 290556 225848
rect 290608 225836 290614 225888
rect 294966 225836 294972 225888
rect 295024 225876 295030 225888
rect 325970 225876 325976 225888
rect 295024 225848 325976 225876
rect 295024 225836 295030 225848
rect 325970 225836 325976 225848
rect 326028 225836 326034 225888
rect 340138 225836 340144 225888
rect 340196 225876 340202 225888
rect 344986 225876 345014 225984
rect 347866 225972 347872 225984
rect 347924 225972 347930 226024
rect 349062 225972 349068 226024
rect 349120 226012 349126 226024
rect 367186 226012 367192 226024
rect 349120 225984 367192 226012
rect 349120 225972 349126 225984
rect 367186 225972 367192 225984
rect 367244 225972 367250 226024
rect 518526 225972 518532 226024
rect 518584 226012 518590 226024
rect 541434 226012 541440 226024
rect 518584 225984 541440 226012
rect 518584 225972 518590 225984
rect 541434 225972 541440 225984
rect 541492 225972 541498 226024
rect 544194 225972 544200 226024
rect 544252 226012 544258 226024
rect 561950 226012 561956 226024
rect 544252 225984 561956 226012
rect 544252 225972 544258 225984
rect 561950 225972 561956 225984
rect 562008 225972 562014 226024
rect 340196 225848 345014 225876
rect 340196 225836 340202 225848
rect 347038 225836 347044 225888
rect 347096 225876 347102 225888
rect 365898 225876 365904 225888
rect 347096 225848 365904 225876
rect 347096 225836 347102 225848
rect 365898 225836 365904 225848
rect 365956 225836 365962 225888
rect 367646 225836 367652 225888
rect 367704 225876 367710 225888
rect 379606 225876 379612 225888
rect 367704 225848 379612 225876
rect 367704 225836 367710 225848
rect 379606 225836 379612 225848
rect 379664 225836 379670 225888
rect 488902 225836 488908 225888
rect 488960 225876 488966 225888
rect 503070 225876 503076 225888
rect 488960 225848 503076 225876
rect 488960 225836 488966 225848
rect 503070 225836 503076 225848
rect 503128 225836 503134 225888
rect 528186 225836 528192 225888
rect 528244 225876 528250 225888
rect 554038 225876 554044 225888
rect 528244 225848 554044 225876
rect 528244 225836 528250 225848
rect 554038 225836 554044 225848
rect 554096 225836 554102 225888
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 671820 225752 671872 225758
rect 242894 225740 242900 225752
rect 186924 225712 232728 225740
rect 232792 225712 242900 225740
rect 186924 225700 186930 225712
rect 61286 225564 61292 225616
rect 61344 225604 61350 225616
rect 136818 225604 136824 225616
rect 61344 225576 136824 225604
rect 61344 225564 61350 225576
rect 136818 225564 136824 225576
rect 136876 225564 136882 225616
rect 137002 225564 137008 225616
rect 137060 225604 137066 225616
rect 147030 225604 147036 225616
rect 137060 225576 147036 225604
rect 137060 225564 137066 225576
rect 147030 225564 147036 225576
rect 147088 225564 147094 225616
rect 147398 225564 147404 225616
rect 147456 225604 147462 225616
rect 203886 225604 203892 225616
rect 147456 225576 186544 225604
rect 147456 225564 147462 225576
rect 186516 225536 186544 225576
rect 186792 225576 203892 225604
rect 186792 225536 186820 225576
rect 203886 225564 203892 225576
rect 203944 225564 203950 225616
rect 204898 225564 204904 225616
rect 204956 225604 204962 225616
rect 222470 225604 222476 225616
rect 204956 225576 222476 225604
rect 204956 225564 204962 225576
rect 222470 225564 222476 225576
rect 222528 225564 222534 225616
rect 224218 225564 224224 225616
rect 224276 225604 224282 225616
rect 232792 225604 232820 225712
rect 242894 225700 242900 225712
rect 242952 225700 242958 225752
rect 257706 225700 257712 225752
rect 257764 225740 257770 225752
rect 299566 225740 299572 225752
rect 257764 225712 299572 225740
rect 257764 225700 257770 225712
rect 299566 225700 299572 225712
rect 299624 225700 299630 225752
rect 304902 225700 304908 225752
rect 304960 225740 304966 225752
rect 333698 225740 333704 225752
rect 304960 225712 333704 225740
rect 304960 225700 304966 225712
rect 333698 225700 333704 225712
rect 333756 225700 333762 225752
rect 335262 225700 335268 225752
rect 335320 225740 335326 225752
rect 356882 225740 356888 225752
rect 335320 225712 356888 225740
rect 335320 225700 335326 225712
rect 356882 225700 356888 225712
rect 356940 225700 356946 225752
rect 379330 225700 379336 225752
rect 379388 225740 379394 225752
rect 393590 225740 393596 225752
rect 379388 225712 393596 225740
rect 379388 225700 379394 225712
rect 393590 225700 393596 225712
rect 393648 225700 393654 225752
rect 394602 225700 394608 225752
rect 394660 225740 394666 225752
rect 404538 225740 404544 225752
rect 394660 225712 404544 225740
rect 394660 225700 394666 225712
rect 404538 225700 404544 225712
rect 404596 225700 404602 225752
rect 491478 225700 491484 225752
rect 491536 225740 491542 225752
rect 506842 225740 506848 225752
rect 491536 225712 506848 225740
rect 491536 225700 491542 225712
rect 506842 225700 506848 225712
rect 506900 225700 506906 225752
rect 507302 225700 507308 225752
rect 507360 225740 507366 225752
rect 526346 225740 526352 225752
rect 507360 225712 526352 225740
rect 507360 225700 507366 225712
rect 526346 225700 526352 225712
rect 526404 225700 526410 225752
rect 527542 225700 527548 225752
rect 527600 225740 527606 225752
rect 553302 225740 553308 225752
rect 527600 225712 553308 225740
rect 527600 225700 527606 225712
rect 553302 225700 553308 225712
rect 553360 225700 553366 225752
rect 671820 225694 671872 225700
rect 224276 225576 232820 225604
rect 224276 225564 224282 225576
rect 234338 225564 234344 225616
rect 234396 225604 234402 225616
rect 281534 225604 281540 225616
rect 234396 225576 281540 225604
rect 234396 225564 234402 225576
rect 281534 225564 281540 225576
rect 281592 225564 281598 225616
rect 285490 225564 285496 225616
rect 285548 225604 285554 225616
rect 318886 225604 318892 225616
rect 285548 225576 318892 225604
rect 285548 225564 285554 225576
rect 318886 225564 318892 225576
rect 318944 225564 318950 225616
rect 322842 225564 322848 225616
rect 322900 225604 322906 225616
rect 349798 225604 349804 225616
rect 322900 225576 349804 225604
rect 322900 225564 322906 225576
rect 349798 225564 349804 225576
rect 349856 225564 349862 225616
rect 351178 225564 351184 225616
rect 351236 225604 351242 225616
rect 370406 225604 370412 225616
rect 351236 225576 370412 225604
rect 351236 225564 351242 225576
rect 370406 225564 370412 225576
rect 370464 225564 370470 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 388070 225604 388076 225616
rect 372580 225576 388076 225604
rect 372580 225564 372586 225576
rect 388070 225564 388076 225576
rect 388128 225564 388134 225616
rect 388438 225564 388444 225616
rect 388496 225604 388502 225616
rect 399386 225604 399392 225616
rect 388496 225576 399392 225604
rect 388496 225564 388502 225576
rect 399386 225564 399392 225576
rect 399444 225564 399450 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 489178 225604 489184 225616
rect 477368 225576 489184 225604
rect 477368 225564 477374 225576
rect 489178 225564 489184 225576
rect 489236 225564 489242 225616
rect 495158 225564 495164 225616
rect 495216 225604 495222 225616
rect 509694 225604 509700 225616
rect 495216 225576 509700 225604
rect 495216 225564 495222 225576
rect 509694 225564 509700 225576
rect 509752 225564 509758 225616
rect 510338 225564 510344 225616
rect 510396 225604 510402 225616
rect 530946 225604 530952 225616
rect 510396 225576 530952 225604
rect 510396 225564 510402 225576
rect 530946 225564 530952 225576
rect 531004 225564 531010 225616
rect 532050 225564 532056 225616
rect 532108 225604 532114 225616
rect 558914 225604 558920 225616
rect 532108 225576 558920 225604
rect 532108 225564 532114 225576
rect 558914 225564 558920 225576
rect 558972 225564 558978 225616
rect 186516 225508 186820 225536
rect 671712 225548 671764 225554
rect 671712 225490 671764 225496
rect 103422 225428 103428 225480
rect 103480 225468 103486 225480
rect 108298 225468 108304 225480
rect 103480 225440 108304 225468
rect 103480 225428 103486 225440
rect 108298 225428 108304 225440
rect 108356 225428 108362 225480
rect 127434 225468 127440 225480
rect 113146 225440 127440 225468
rect 105998 225292 106004 225344
rect 106056 225332 106062 225344
rect 113146 225332 113174 225440
rect 127434 225428 127440 225440
rect 127492 225428 127498 225480
rect 181438 225468 181444 225480
rect 127636 225440 181444 225468
rect 106056 225304 113174 225332
rect 106056 225292 106062 225304
rect 117222 225292 117228 225344
rect 117280 225332 117286 225344
rect 127636 225332 127664 225440
rect 181438 225428 181444 225440
rect 181496 225428 181502 225480
rect 183278 225428 183284 225480
rect 183336 225468 183342 225480
rect 185670 225468 185676 225480
rect 183336 225440 185676 225468
rect 183336 225428 183342 225440
rect 185670 225428 185676 225440
rect 185728 225428 185734 225480
rect 190730 225428 190736 225480
rect 190788 225468 190794 225480
rect 242250 225468 242256 225480
rect 190788 225440 242256 225468
rect 190788 225428 190794 225440
rect 242250 225428 242256 225440
rect 242308 225428 242314 225480
rect 668394 225428 668400 225480
rect 668452 225468 668458 225480
rect 668452 225440 671622 225468
rect 668452 225428 668458 225440
rect 185872 225372 187188 225400
rect 137002 225332 137008 225344
rect 117280 225304 127664 225332
rect 127728 225304 137008 225332
rect 117280 225292 117286 225304
rect 127434 225156 127440 225208
rect 127492 225196 127498 225208
rect 127728 225196 127756 225304
rect 137002 225292 137008 225304
rect 137060 225292 137066 225344
rect 142108 225332 142114 225344
rect 137204 225304 142114 225332
rect 127492 225168 127756 225196
rect 127492 225156 127498 225168
rect 128262 225156 128268 225208
rect 128320 225196 128326 225208
rect 137204 225196 137232 225304
rect 142108 225292 142114 225304
rect 142166 225292 142172 225344
rect 142246 225292 142252 225344
rect 142304 225332 142310 225344
rect 185872 225332 185900 225372
rect 142304 225304 185900 225332
rect 187160 225332 187188 225372
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 203150 225332 203156 225344
rect 187160 225304 203156 225332
rect 142304 225292 142310 225304
rect 203150 225292 203156 225304
rect 203208 225292 203214 225344
rect 203886 225292 203892 225344
rect 203944 225332 203950 225344
rect 207750 225332 207756 225344
rect 203944 225304 207756 225332
rect 203944 225292 203950 225304
rect 207750 225292 207756 225304
rect 207808 225292 207814 225344
rect 208026 225292 208032 225344
rect 208084 225332 208090 225344
rect 260926 225332 260932 225344
rect 208084 225304 260932 225332
rect 208084 225292 208090 225304
rect 260926 225292 260932 225304
rect 260984 225292 260990 225344
rect 671062 225224 671068 225276
rect 671120 225264 671126 225276
rect 671120 225236 671508 225264
rect 671120 225224 671126 225236
rect 186866 225196 186872 225208
rect 128320 225168 137232 225196
rect 137296 225168 186872 225196
rect 128320 225156 128326 225168
rect 126882 225020 126888 225072
rect 126940 225060 126946 225072
rect 137296 225060 137324 225168
rect 186866 225156 186872 225168
rect 186924 225156 186930 225208
rect 187234 225156 187240 225208
rect 187292 225196 187298 225208
rect 195882 225196 195888 225208
rect 187292 225168 195888 225196
rect 187292 225156 187298 225168
rect 195882 225156 195888 225168
rect 195940 225156 195946 225208
rect 199378 225156 199384 225208
rect 199436 225196 199442 225208
rect 204898 225196 204904 225208
rect 199436 225168 204904 225196
rect 199436 225156 199442 225168
rect 204898 225156 204904 225168
rect 204956 225156 204962 225208
rect 205082 225156 205088 225208
rect 205140 225196 205146 225208
rect 254486 225196 254492 225208
rect 205140 225168 254492 225196
rect 205140 225156 205146 225168
rect 254486 225156 254492 225168
rect 254544 225156 254550 225208
rect 126940 225032 137324 225060
rect 126940 225020 126946 225032
rect 137462 225020 137468 225072
rect 137520 225060 137526 225072
rect 141510 225060 141516 225072
rect 137520 225032 141516 225060
rect 137520 225020 137526 225032
rect 141510 225020 141516 225032
rect 141568 225020 141574 225072
rect 141786 225020 141792 225072
rect 141844 225060 141850 225072
rect 141844 225032 142292 225060
rect 141844 225020 141850 225032
rect 116762 224884 116768 224936
rect 116820 224924 116826 224936
rect 122926 224924 122932 224936
rect 116820 224896 122932 224924
rect 116820 224884 116826 224896
rect 122926 224884 122932 224896
rect 122984 224884 122990 224936
rect 123478 224884 123484 224936
rect 123536 224924 123542 224936
rect 142062 224924 142068 224936
rect 123536 224896 142068 224924
rect 123536 224884 123542 224896
rect 142062 224884 142068 224896
rect 142120 224884 142126 224936
rect 142264 224924 142292 225032
rect 142430 225020 142436 225072
rect 142488 225060 142494 225072
rect 162302 225060 162308 225072
rect 142488 225032 162308 225060
rect 142488 225020 142494 225032
rect 162302 225020 162308 225032
rect 162360 225020 162366 225072
rect 162486 225020 162492 225072
rect 162544 225060 162550 225072
rect 166534 225060 166540 225072
rect 162544 225032 166540 225060
rect 162544 225020 162550 225032
rect 166534 225020 166540 225032
rect 166592 225020 166598 225072
rect 166718 225020 166724 225072
rect 166776 225060 166782 225072
rect 169018 225060 169024 225072
rect 166776 225032 169024 225060
rect 166776 225020 166782 225032
rect 169018 225020 169024 225032
rect 169076 225020 169082 225072
rect 169202 225020 169208 225072
rect 169260 225060 169266 225072
rect 170858 225060 170864 225072
rect 169260 225032 170864 225060
rect 169260 225020 169266 225032
rect 170858 225020 170864 225032
rect 170916 225020 170922 225072
rect 171042 225020 171048 225072
rect 171100 225060 171106 225072
rect 223574 225060 223580 225072
rect 171100 225032 223580 225060
rect 171100 225020 171106 225032
rect 223574 225020 223580 225032
rect 223632 225020 223638 225072
rect 224862 225020 224868 225072
rect 224920 225060 224926 225072
rect 270586 225060 270592 225072
rect 224920 225032 270592 225060
rect 224920 225020 224926 225032
rect 270586 225020 270592 225032
rect 270644 225020 270650 225072
rect 669406 225020 669412 225072
rect 669464 225060 669470 225072
rect 669464 225032 671398 225060
rect 669464 225020 669470 225032
rect 275830 224952 275836 225004
rect 275888 224992 275894 225004
rect 276290 224992 276296 225004
rect 275888 224964 276296 224992
rect 275888 224952 275894 224964
rect 276290 224952 276296 224964
rect 276348 224952 276354 225004
rect 282730 224952 282736 225004
rect 282788 224992 282794 225004
rect 285306 224992 285312 225004
rect 282788 224964 285312 224992
rect 282788 224952 282794 224964
rect 285306 224952 285312 224964
rect 285364 224952 285370 225004
rect 489914 224952 489920 225004
rect 489972 224992 489978 225004
rect 494790 224992 494796 225004
rect 489972 224964 494796 224992
rect 489972 224952 489978 224964
rect 494790 224952 494796 224964
rect 494848 224952 494854 225004
rect 509234 224952 509240 225004
rect 509292 224992 509298 225004
rect 512638 224992 512644 225004
rect 509292 224964 512644 224992
rect 509292 224952 509298 224964
rect 512638 224952 512644 224964
rect 512696 224952 512702 225004
rect 209406 224924 209412 224936
rect 142264 224896 209412 224924
rect 209406 224884 209412 224896
rect 209464 224884 209470 224936
rect 209682 224884 209688 224936
rect 209740 224924 209746 224936
rect 259638 224924 259644 224936
rect 209740 224896 259644 224924
rect 209740 224884 209746 224896
rect 259638 224884 259644 224896
rect 259696 224884 259702 224936
rect 264146 224884 264152 224936
rect 264204 224924 264210 224936
rect 269298 224924 269304 224936
rect 264204 224896 269304 224924
rect 264204 224884 264210 224896
rect 269298 224884 269304 224896
rect 269356 224884 269362 224936
rect 288342 224884 288348 224936
rect 288400 224924 288406 224936
rect 322382 224924 322388 224936
rect 288400 224896 322388 224924
rect 288400 224884 288406 224896
rect 322382 224884 322388 224896
rect 322440 224884 322446 224936
rect 406746 224884 406752 224936
rect 406804 224924 406810 224936
rect 414842 224924 414848 224936
rect 406804 224896 414848 224924
rect 406804 224884 406810 224896
rect 414842 224884 414848 224896
rect 414900 224884 414906 224936
rect 516502 224884 516508 224936
rect 516560 224924 516566 224936
rect 531314 224924 531320 224936
rect 516560 224896 531320 224924
rect 516560 224884 516566 224896
rect 531314 224884 531320 224896
rect 531372 224884 531378 224936
rect 669406 224816 669412 224868
rect 669464 224856 669470 224868
rect 669464 224828 671278 224856
rect 669464 224816 669470 224828
rect 118602 224748 118608 224800
rect 118660 224788 118666 224800
rect 177206 224788 177212 224800
rect 118660 224760 177212 224788
rect 118660 224748 118666 224760
rect 177206 224748 177212 224760
rect 177264 224748 177270 224800
rect 177390 224748 177396 224800
rect 177448 224788 177454 224800
rect 181254 224788 181260 224800
rect 177448 224760 181260 224788
rect 177448 224748 177454 224760
rect 181254 224748 181260 224760
rect 181312 224748 181318 224800
rect 187050 224788 187056 224800
rect 181456 224760 187056 224788
rect 115750 224612 115756 224664
rect 115808 224652 115814 224664
rect 181456 224652 181484 224760
rect 187050 224748 187056 224760
rect 187108 224748 187114 224800
rect 187326 224748 187332 224800
rect 187384 224788 187390 224800
rect 190730 224788 190736 224800
rect 187384 224760 190736 224788
rect 187384 224748 187390 224760
rect 190730 224748 190736 224760
rect 190788 224748 190794 224800
rect 194502 224748 194508 224800
rect 194560 224788 194566 224800
rect 247402 224788 247408 224800
rect 194560 224760 247408 224788
rect 194560 224748 194566 224760
rect 247402 224748 247408 224760
rect 247460 224748 247466 224800
rect 282546 224748 282552 224800
rect 282604 224788 282610 224800
rect 316310 224788 316316 224800
rect 282604 224760 316316 224788
rect 282604 224748 282610 224760
rect 316310 224748 316316 224760
rect 316368 224748 316374 224800
rect 532418 224748 532424 224800
rect 532476 224788 532482 224800
rect 550450 224788 550456 224800
rect 532476 224760 550456 224788
rect 532476 224748 532482 224760
rect 550450 224748 550456 224760
rect 550508 224748 550514 224800
rect 460566 224680 460572 224732
rect 460624 224720 460630 224732
rect 463142 224720 463148 224732
rect 460624 224692 463148 224720
rect 460624 224680 460630 224692
rect 463142 224680 463148 224692
rect 463200 224680 463206 224732
rect 191374 224652 191380 224664
rect 115808 224624 181484 224652
rect 181548 224624 191380 224652
rect 115808 224612 115814 224624
rect 60642 224476 60648 224528
rect 60700 224516 60706 224528
rect 103606 224516 103612 224528
rect 60700 224488 103612 224516
rect 60700 224476 60706 224488
rect 103606 224476 103612 224488
rect 103664 224476 103670 224528
rect 108666 224476 108672 224528
rect 108724 224516 108730 224528
rect 177022 224516 177028 224528
rect 108724 224488 177028 224516
rect 108724 224476 108730 224488
rect 177022 224476 177028 224488
rect 177080 224476 177086 224528
rect 177206 224476 177212 224528
rect 177264 224516 177270 224528
rect 181548 224516 181576 224624
rect 191374 224612 191380 224624
rect 191432 224612 191438 224664
rect 192754 224612 192760 224664
rect 192812 224652 192818 224664
rect 194318 224652 194324 224664
rect 192812 224624 194324 224652
rect 192812 224612 192818 224624
rect 194318 224612 194324 224624
rect 194376 224612 194382 224664
rect 195606 224612 195612 224664
rect 195664 224652 195670 224664
rect 248874 224652 248880 224664
rect 195664 224624 248880 224652
rect 195664 224612 195670 224624
rect 248874 224612 248880 224624
rect 248932 224612 248938 224664
rect 249058 224612 249064 224664
rect 249116 224652 249122 224664
rect 263870 224652 263876 224664
rect 249116 224624 263876 224652
rect 249116 224612 249122 224624
rect 263870 224612 263876 224624
rect 263928 224612 263934 224664
rect 271598 224612 271604 224664
rect 271656 224652 271662 224664
rect 309870 224652 309876 224664
rect 271656 224624 309876 224652
rect 271656 224612 271662 224624
rect 309870 224612 309876 224624
rect 309928 224612 309934 224664
rect 315850 224612 315856 224664
rect 315908 224652 315914 224664
rect 341426 224652 341432 224664
rect 315908 224624 341432 224652
rect 315908 224612 315914 224624
rect 341426 224612 341432 224624
rect 341484 224612 341490 224664
rect 344646 224612 344652 224664
rect 344704 224652 344710 224664
rect 364610 224652 364616 224664
rect 344704 224624 364616 224652
rect 344704 224612 344710 224624
rect 364610 224612 364616 224624
rect 364668 224612 364674 224664
rect 514662 224612 514668 224664
rect 514720 224652 514726 224664
rect 536650 224652 536656 224664
rect 514720 224624 536656 224652
rect 514720 224612 514726 224624
rect 536650 224612 536656 224624
rect 536708 224612 536714 224664
rect 668394 224612 668400 224664
rect 668452 224652 668458 224664
rect 668452 224624 671186 224652
rect 668452 224612 668458 224624
rect 456058 224544 456064 224596
rect 456116 224584 456122 224596
rect 459646 224584 459652 224596
rect 456116 224556 459652 224584
rect 456116 224544 456122 224556
rect 459646 224544 459652 224556
rect 459704 224544 459710 224596
rect 177264 224488 181576 224516
rect 177264 224476 177270 224488
rect 181714 224476 181720 224528
rect 181772 224516 181778 224528
rect 183830 224516 183836 224528
rect 181772 224488 183836 224516
rect 181772 224476 181778 224488
rect 183830 224476 183836 224488
rect 183888 224476 183894 224528
rect 184014 224476 184020 224528
rect 184072 224516 184078 224528
rect 233694 224516 233700 224528
rect 184072 224488 233700 224516
rect 184072 224476 184078 224488
rect 233694 224476 233700 224488
rect 233752 224476 233758 224528
rect 233878 224476 233884 224528
rect 233936 224516 233942 224528
rect 246758 224516 246764 224528
rect 233936 224488 246764 224516
rect 233936 224476 233942 224488
rect 246758 224476 246764 224488
rect 246816 224476 246822 224528
rect 247678 224476 247684 224528
rect 247736 224516 247742 224528
rect 289262 224516 289268 224528
rect 247736 224488 289268 224516
rect 247736 224476 247742 224488
rect 289262 224476 289268 224488
rect 289320 224476 289326 224528
rect 319990 224476 319996 224528
rect 320048 224516 320054 224528
rect 347222 224516 347228 224528
rect 320048 224488 347228 224516
rect 320048 224476 320054 224488
rect 347222 224476 347228 224488
rect 347280 224476 347286 224528
rect 479518 224476 479524 224528
rect 479576 224516 479582 224528
rect 486602 224516 486608 224528
rect 479576 224488 486608 224516
rect 479576 224476 479582 224488
rect 486602 224476 486608 224488
rect 486660 224476 486666 224528
rect 508222 224476 508228 224528
rect 508280 224516 508286 224528
rect 528370 224516 528376 224528
rect 508280 224488 528376 224516
rect 508280 224476 508286 224488
rect 528370 224476 528376 224488
rect 528428 224476 528434 224528
rect 530118 224476 530124 224528
rect 530176 224516 530182 224528
rect 556522 224516 556528 224528
rect 530176 224488 556528 224516
rect 530176 224476 530182 224488
rect 556522 224476 556528 224488
rect 556580 224476 556586 224528
rect 670712 224420 671048 224448
rect 82722 224340 82728 224392
rect 82780 224380 82786 224392
rect 123478 224380 123484 224392
rect 82780 224352 123484 224380
rect 82780 224340 82786 224352
rect 123478 224340 123484 224352
rect 123536 224340 123542 224392
rect 131298 224340 131304 224392
rect 131356 224380 131362 224392
rect 193950 224380 193956 224392
rect 131356 224352 193956 224380
rect 131356 224340 131362 224352
rect 193950 224340 193956 224352
rect 194008 224340 194014 224392
rect 194134 224340 194140 224392
rect 194192 224380 194198 224392
rect 204898 224380 204904 224392
rect 194192 224352 204904 224380
rect 194192 224340 194198 224352
rect 204898 224340 204904 224352
rect 204956 224340 204962 224392
rect 205082 224340 205088 224392
rect 205140 224380 205146 224392
rect 255774 224380 255780 224392
rect 205140 224352 255780 224380
rect 205140 224340 205146 224352
rect 255774 224340 255780 224352
rect 255832 224340 255838 224392
rect 261846 224340 261852 224392
rect 261904 224380 261910 224392
rect 300854 224380 300860 224392
rect 261904 224352 300860 224380
rect 261904 224340 261910 224352
rect 300854 224340 300860 224352
rect 300912 224340 300918 224392
rect 303246 224340 303252 224392
rect 303304 224380 303310 224392
rect 333054 224380 333060 224392
rect 303304 224352 333060 224380
rect 303304 224340 303310 224352
rect 333054 224340 333060 224352
rect 333112 224340 333118 224392
rect 333882 224340 333888 224392
rect 333940 224380 333946 224392
rect 356238 224380 356244 224392
rect 333940 224352 356244 224380
rect 333940 224340 333946 224352
rect 356238 224340 356244 224352
rect 356296 224340 356302 224392
rect 357342 224340 357348 224392
rect 357400 224380 357406 224392
rect 374270 224380 374276 224392
rect 357400 224352 374276 224380
rect 357400 224340 357406 224352
rect 374270 224340 374276 224352
rect 374328 224340 374334 224392
rect 375282 224340 375288 224392
rect 375340 224380 375346 224392
rect 387794 224380 387800 224392
rect 375340 224352 387800 224380
rect 375340 224340 375346 224352
rect 387794 224340 387800 224352
rect 387852 224340 387858 224392
rect 462498 224340 462504 224392
rect 462556 224380 462562 224392
rect 469306 224380 469312 224392
rect 462556 224352 469312 224380
rect 462556 224340 462562 224352
rect 469306 224340 469312 224352
rect 469364 224340 469370 224392
rect 470226 224340 470232 224392
rect 470284 224380 470290 224392
rect 479702 224380 479708 224392
rect 470284 224352 479708 224380
rect 470284 224340 470290 224352
rect 479702 224340 479708 224352
rect 479760 224340 479766 224392
rect 486786 224340 486792 224392
rect 486844 224380 486850 224392
rect 496906 224380 496912 224392
rect 486844 224352 496912 224380
rect 486844 224340 486850 224352
rect 496906 224340 496912 224352
rect 496964 224340 496970 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525702 224340 525708 224392
rect 525760 224380 525766 224392
rect 550634 224380 550640 224392
rect 525760 224352 550640 224380
rect 525760 224340 525766 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 58986 224204 58992 224256
rect 59044 224244 59050 224256
rect 145190 224244 145196 224256
rect 59044 224216 145196 224244
rect 59044 224204 59050 224216
rect 145190 224204 145196 224216
rect 145248 224204 145254 224256
rect 145374 224204 145380 224256
rect 145432 224244 145438 224256
rect 147214 224244 147220 224256
rect 145432 224216 147220 224244
rect 145432 224204 145438 224216
rect 147214 224204 147220 224216
rect 147272 224204 147278 224256
rect 147766 224204 147772 224256
rect 147824 224244 147830 224256
rect 156690 224244 156696 224256
rect 147824 224216 156696 224244
rect 147824 224204 147830 224216
rect 156690 224204 156696 224216
rect 156748 224204 156754 224256
rect 157426 224204 157432 224256
rect 157484 224244 157490 224256
rect 170950 224244 170956 224256
rect 157484 224216 170956 224244
rect 157484 224204 157490 224216
rect 170950 224204 170956 224216
rect 171008 224204 171014 224256
rect 171088 224204 171094 224256
rect 171146 224244 171152 224256
rect 186866 224244 186872 224256
rect 171146 224216 186872 224244
rect 171146 224204 171152 224216
rect 186866 224204 186872 224216
rect 186924 224204 186930 224256
rect 187050 224204 187056 224256
rect 187108 224244 187114 224256
rect 188798 224244 188804 224256
rect 187108 224216 188804 224244
rect 187108 224204 187114 224216
rect 188798 224204 188804 224216
rect 188856 224204 188862 224256
rect 188982 224204 188988 224256
rect 189040 224244 189046 224256
rect 243814 224244 243820 224256
rect 189040 224216 243820 224244
rect 189040 224204 189046 224216
rect 243814 224204 243820 224216
rect 243872 224204 243878 224256
rect 246942 224204 246948 224256
rect 247000 224244 247006 224256
rect 288618 224244 288624 224256
rect 247000 224216 288624 224244
rect 247000 224204 247006 224216
rect 288618 224204 288624 224216
rect 288676 224204 288682 224256
rect 289630 224204 289636 224256
rect 289688 224244 289694 224256
rect 308122 224244 308128 224256
rect 289688 224216 308128 224244
rect 289688 224204 289694 224216
rect 308122 224204 308128 224216
rect 308180 224204 308186 224256
rect 308950 224204 308956 224256
rect 309008 224244 309014 224256
rect 339494 224244 339500 224256
rect 309008 224216 339500 224244
rect 309008 224204 309014 224216
rect 339494 224204 339500 224216
rect 339552 224204 339558 224256
rect 342070 224204 342076 224256
rect 342128 224244 342134 224256
rect 364794 224244 364800 224256
rect 342128 224216 364800 224244
rect 342128 224204 342134 224216
rect 364794 224204 364800 224216
rect 364852 224204 364858 224256
rect 364978 224204 364984 224256
rect 365036 224244 365042 224256
rect 378134 224244 378140 224256
rect 365036 224216 378140 224244
rect 365036 224204 365042 224216
rect 378134 224204 378140 224216
rect 378192 224204 378198 224256
rect 389082 224204 389088 224256
rect 389140 224244 389146 224256
rect 400950 224244 400956 224256
rect 389140 224216 400956 224244
rect 389140 224204 389146 224216
rect 400950 224204 400956 224216
rect 401008 224204 401014 224256
rect 416498 224204 416504 224256
rect 416556 224244 416562 224256
rect 422202 224244 422208 224256
rect 416556 224216 422208 224244
rect 416556 224204 416562 224216
rect 422202 224204 422208 224216
rect 422260 224204 422266 224256
rect 423306 224204 423312 224256
rect 423364 224244 423370 224256
rect 424318 224244 424324 224256
rect 423364 224216 424324 224244
rect 423364 224204 423370 224216
rect 424318 224204 424324 224216
rect 424376 224204 424382 224256
rect 451366 224204 451372 224256
rect 451424 224244 451430 224256
rect 452194 224244 452200 224256
rect 451424 224216 452200 224244
rect 451424 224204 451430 224216
rect 452194 224204 452200 224216
rect 452252 224204 452258 224256
rect 474734 224204 474740 224256
rect 474792 224244 474798 224256
rect 484578 224244 484584 224256
rect 474792 224216 484584 224244
rect 474792 224204 474798 224216
rect 484578 224204 484584 224216
rect 484636 224204 484642 224256
rect 485682 224204 485688 224256
rect 485740 224244 485746 224256
rect 499390 224244 499396 224256
rect 485740 224216 499396 224244
rect 485740 224204 485746 224216
rect 499390 224204 499396 224216
rect 499448 224204 499454 224256
rect 508866 224204 508872 224256
rect 508924 224244 508930 224256
rect 529198 224244 529204 224256
rect 508924 224216 529204 224244
rect 508924 224204 508930 224216
rect 529198 224204 529204 224216
rect 529256 224204 529262 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 563698 224244 563704 224256
rect 535328 224216 563704 224244
rect 535328 224204 535334 224216
rect 563698 224204 563704 224216
rect 563756 224204 563762 224256
rect 104802 224068 104808 224120
rect 104860 224108 104866 224120
rect 116762 224108 116768 224120
rect 104860 224080 116768 224108
rect 104860 224068 104866 224080
rect 116762 224068 116768 224080
rect 116820 224068 116826 224120
rect 116946 224068 116952 224120
rect 117004 224108 117010 224120
rect 118418 224108 118424 224120
rect 117004 224080 118424 224108
rect 117004 224068 117010 224080
rect 118418 224068 118424 224080
rect 118476 224068 118482 224120
rect 121914 224068 121920 224120
rect 121972 224108 121978 224120
rect 131298 224108 131304 224120
rect 121972 224080 131304 224108
rect 121972 224068 121978 224080
rect 131298 224068 131304 224080
rect 131356 224068 131362 224120
rect 131482 224068 131488 224120
rect 131540 224108 131546 224120
rect 192754 224108 192760 224120
rect 131540 224080 192760 224108
rect 131540 224068 131546 224080
rect 192754 224068 192760 224080
rect 192812 224068 192818 224120
rect 192938 224068 192944 224120
rect 192996 224108 193002 224120
rect 194134 224108 194140 224120
rect 192996 224080 194140 224108
rect 192996 224068 193002 224080
rect 194134 224068 194140 224080
rect 194192 224068 194198 224120
rect 194318 224068 194324 224120
rect 194376 224108 194382 224120
rect 196526 224108 196532 224120
rect 194376 224080 196532 224108
rect 194376 224068 194382 224080
rect 196526 224068 196532 224080
rect 196584 224068 196590 224120
rect 201218 224068 201224 224120
rect 201276 224108 201282 224120
rect 204714 224108 204720 224120
rect 201276 224080 204720 224108
rect 201276 224068 201282 224080
rect 204714 224068 204720 224080
rect 204772 224068 204778 224120
rect 204898 224068 204904 224120
rect 204956 224108 204962 224120
rect 233878 224108 233884 224120
rect 204956 224080 233884 224108
rect 204956 224068 204962 224080
rect 233878 224068 233884 224080
rect 233936 224068 233942 224120
rect 278958 224108 278964 224120
rect 235276 224080 278964 224108
rect 76558 223932 76564 223984
rect 76616 223972 76622 223984
rect 140958 223972 140964 223984
rect 76616 223944 140964 223972
rect 76616 223932 76622 223944
rect 140958 223932 140964 223944
rect 141016 223932 141022 223984
rect 142062 223932 142068 223984
rect 142120 223972 142126 223984
rect 157058 223972 157064 223984
rect 142120 223944 157064 223972
rect 142120 223932 142126 223944
rect 157058 223932 157064 223944
rect 157116 223932 157122 223984
rect 157242 223932 157248 223984
rect 157300 223972 157306 223984
rect 217134 223972 217140 223984
rect 157300 223944 217140 223972
rect 157300 223932 157306 223944
rect 217134 223932 217140 223944
rect 217192 223932 217198 223984
rect 217318 223932 217324 223984
rect 217376 223972 217382 223984
rect 228082 223972 228088 223984
rect 217376 223944 228088 223972
rect 217376 223932 217382 223944
rect 228082 223932 228088 223944
rect 228140 223932 228146 223984
rect 231670 223932 231676 223984
rect 231728 223972 231734 223984
rect 235276 223972 235304 224080
rect 278958 224068 278964 224080
rect 279016 224068 279022 224120
rect 286686 224068 286692 224120
rect 286744 224108 286750 224120
rect 319530 224108 319536 224120
rect 286744 224080 319536 224108
rect 286744 224068 286750 224080
rect 319530 224068 319536 224080
rect 319588 224068 319594 224120
rect 670712 223984 670740 224420
rect 670930 224324 670982 224330
rect 670930 224266 670982 224272
rect 231728 223944 235304 223972
rect 231728 223932 231734 223944
rect 238662 223932 238668 223984
rect 238720 223972 238726 223984
rect 282362 223972 282368 223984
rect 238720 223944 282368 223972
rect 238720 223932 238726 223944
rect 282362 223932 282368 223944
rect 282420 223932 282426 223984
rect 670694 223932 670700 223984
rect 670752 223932 670758 223984
rect 125226 223796 125232 223848
rect 125284 223836 125290 223848
rect 131482 223836 131488 223848
rect 125284 223808 131488 223836
rect 125284 223796 125290 223808
rect 131482 223796 131488 223808
rect 131540 223796 131546 223848
rect 134426 223796 134432 223848
rect 134484 223836 134490 223848
rect 204254 223836 204260 223848
rect 134484 223808 204260 223836
rect 134484 223796 134490 223808
rect 204254 223796 204260 223808
rect 204312 223796 204318 223848
rect 205266 223796 205272 223848
rect 205324 223836 205330 223848
rect 212626 223836 212632 223848
rect 205324 223808 212632 223836
rect 205324 223796 205330 223808
rect 212626 223796 212632 223808
rect 212684 223796 212690 223848
rect 215938 223796 215944 223848
rect 215996 223836 216002 223848
rect 222930 223836 222936 223848
rect 215996 223808 222936 223836
rect 215996 223796 216002 223808
rect 222930 223796 222936 223808
rect 222988 223796 222994 223848
rect 233694 223796 233700 223848
rect 233752 223836 233758 223848
rect 239674 223836 239680 223848
rect 233752 223808 239680 223836
rect 233752 223796 233758 223808
rect 239674 223796 239680 223808
rect 239732 223796 239738 223848
rect 241974 223796 241980 223848
rect 242032 223836 242038 223848
rect 285030 223836 285036 223848
rect 242032 223808 285036 223836
rect 242032 223796 242038 223808
rect 285030 223796 285036 223808
rect 285088 223796 285094 223848
rect 126698 223660 126704 223712
rect 126756 223700 126762 223712
rect 131114 223700 131120 223712
rect 126756 223672 131120 223700
rect 126756 223660 126762 223672
rect 131114 223660 131120 223672
rect 131172 223660 131178 223712
rect 132402 223660 132408 223712
rect 132460 223700 132466 223712
rect 201678 223700 201684 223712
rect 132460 223672 201684 223700
rect 132460 223660 132466 223672
rect 201678 223660 201684 223672
rect 201736 223660 201742 223712
rect 297836 223672 300348 223700
rect 87966 223524 87972 223576
rect 88024 223564 88030 223576
rect 88024 223536 161152 223564
rect 88024 223524 88030 223536
rect 81342 223388 81348 223440
rect 81400 223428 81406 223440
rect 157242 223428 157248 223440
rect 81400 223400 157248 223428
rect 81400 223388 81406 223400
rect 157242 223388 157248 223400
rect 157300 223388 157306 223440
rect 157426 223388 157432 223440
rect 157484 223428 157490 223440
rect 159818 223428 159824 223440
rect 157484 223400 159824 223428
rect 157484 223388 157490 223400
rect 159818 223388 159824 223400
rect 159876 223388 159882 223440
rect 161124 223428 161152 223536
rect 161934 223524 161940 223576
rect 161992 223564 161998 223576
rect 167822 223564 167828 223576
rect 161992 223536 167828 223564
rect 161992 223524 161998 223536
rect 167822 223524 167828 223536
rect 167880 223524 167886 223576
rect 168282 223524 168288 223576
rect 168340 223564 168346 223576
rect 226702 223564 226708 223576
rect 168340 223536 226708 223564
rect 168340 223524 168346 223536
rect 226702 223524 226708 223536
rect 226760 223524 226766 223576
rect 269022 223524 269028 223576
rect 269080 223564 269086 223576
rect 297836 223564 297864 223672
rect 269080 223536 297864 223564
rect 269080 223524 269086 223536
rect 298002 223524 298008 223576
rect 298060 223564 298066 223576
rect 300118 223564 300124 223576
rect 298060 223536 300124 223564
rect 298060 223524 298066 223536
rect 300118 223524 300124 223536
rect 300176 223524 300182 223576
rect 300320 223564 300348 223672
rect 426434 223592 426440 223644
rect 426492 223632 426498 223644
rect 426986 223632 426992 223644
rect 426492 223604 426992 223632
rect 426492 223592 426498 223604
rect 426986 223592 426992 223604
rect 427044 223592 427050 223644
rect 306006 223564 306012 223576
rect 300320 223536 306012 223564
rect 306006 223524 306012 223536
rect 306064 223524 306070 223576
rect 329098 223524 329104 223576
rect 329156 223564 329162 223576
rect 342714 223564 342720 223576
rect 329156 223536 342720 223564
rect 329156 223524 329162 223536
rect 342714 223524 342720 223536
rect 342772 223524 342778 223576
rect 457990 223524 457996 223576
rect 458048 223564 458054 223576
rect 460198 223564 460204 223576
rect 458048 223536 460204 223564
rect 458048 223524 458054 223536
rect 460198 223524 460204 223536
rect 460256 223524 460262 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 679250 223524 679256 223576
rect 679308 223564 679314 223576
rect 680170 223564 680176 223576
rect 679308 223536 680176 223564
rect 679308 223524 679314 223536
rect 680170 223524 680176 223536
rect 680228 223524 680234 223576
rect 164970 223428 164976 223440
rect 161124 223400 164976 223428
rect 164970 223388 164976 223400
rect 165028 223388 165034 223440
rect 165246 223388 165252 223440
rect 165304 223428 165310 223440
rect 224034 223428 224040 223440
rect 165304 223400 224040 223428
rect 165304 223388 165310 223400
rect 224034 223388 224040 223400
rect 224092 223388 224098 223440
rect 260098 223388 260104 223440
rect 260156 223428 260162 223440
rect 298922 223428 298928 223440
rect 260156 223400 298928 223428
rect 260156 223388 260162 223400
rect 298922 223388 298928 223400
rect 298980 223388 298986 223440
rect 302142 223388 302148 223440
rect 302200 223428 302206 223440
rect 331122 223428 331128 223440
rect 302200 223400 331128 223428
rect 302200 223388 302206 223400
rect 331122 223388 331128 223400
rect 331180 223388 331186 223440
rect 518894 223388 518900 223440
rect 518952 223428 518958 223440
rect 530026 223428 530032 223440
rect 518952 223400 530032 223428
rect 518952 223388 518958 223400
rect 530026 223388 530032 223400
rect 530084 223388 530090 223440
rect 92106 223252 92112 223304
rect 92164 223292 92170 223304
rect 166810 223292 166816 223304
rect 92164 223264 166816 223292
rect 92164 223252 92170 223264
rect 166810 223252 166816 223264
rect 166868 223252 166874 223304
rect 166948 223252 166954 223304
rect 167006 223292 167012 223304
rect 176102 223292 176108 223304
rect 167006 223264 176108 223292
rect 167006 223252 167012 223264
rect 176102 223252 176108 223264
rect 176160 223252 176166 223304
rect 176286 223252 176292 223304
rect 176344 223292 176350 223304
rect 181438 223292 181444 223304
rect 176344 223264 181444 223292
rect 176344 223252 176350 223264
rect 181438 223252 181444 223264
rect 181496 223252 181502 223304
rect 181622 223252 181628 223304
rect 181680 223292 181686 223304
rect 192018 223292 192024 223304
rect 181680 223264 192024 223292
rect 181680 223252 181686 223264
rect 192018 223252 192024 223264
rect 192076 223252 192082 223304
rect 203886 223252 203892 223304
rect 203944 223292 203950 223304
rect 254854 223292 254860 223304
rect 203944 223264 254860 223292
rect 203944 223252 203950 223264
rect 254854 223252 254860 223264
rect 254912 223252 254918 223304
rect 264790 223252 264796 223304
rect 264848 223292 264854 223304
rect 304718 223292 304724 223304
rect 264848 223264 304724 223292
rect 264848 223252 264854 223264
rect 304718 223252 304724 223264
rect 304776 223252 304782 223304
rect 306282 223252 306288 223304
rect 306340 223292 306346 223304
rect 336918 223292 336924 223304
rect 306340 223264 336924 223292
rect 306340 223252 306346 223264
rect 336918 223252 336924 223264
rect 336976 223252 336982 223304
rect 343542 223252 343548 223304
rect 343600 223292 343606 223304
rect 363966 223292 363972 223304
rect 343600 223264 363972 223292
rect 343600 223252 343606 223264
rect 363966 223252 363972 223264
rect 364024 223252 364030 223304
rect 489546 223252 489552 223304
rect 489604 223292 489610 223304
rect 504358 223292 504364 223304
rect 489604 223264 504364 223292
rect 489604 223252 489610 223264
rect 504358 223252 504364 223264
rect 504416 223252 504422 223304
rect 505094 223252 505100 223304
rect 505152 223292 505158 223304
rect 524230 223292 524236 223304
rect 505152 223264 524236 223292
rect 505152 223252 505158 223264
rect 524230 223252 524236 223264
rect 524288 223252 524294 223304
rect 529014 223252 529020 223304
rect 529072 223292 529078 223304
rect 542446 223292 542452 223304
rect 529072 223264 542452 223292
rect 529072 223252 529078 223264
rect 542446 223252 542452 223264
rect 542504 223252 542510 223304
rect 78582 223116 78588 223168
rect 78640 223156 78646 223168
rect 156874 223156 156880 223168
rect 78640 223128 156880 223156
rect 78640 223116 78646 223128
rect 156874 223116 156880 223128
rect 156932 223116 156938 223168
rect 157058 223116 157064 223168
rect 157116 223156 157122 223168
rect 162118 223156 162124 223168
rect 157116 223128 162124 223156
rect 157116 223116 157122 223128
rect 162118 223116 162124 223128
rect 162176 223116 162182 223168
rect 164142 223116 164148 223168
rect 164200 223156 164206 223168
rect 165246 223156 165252 223168
rect 164200 223128 165252 223156
rect 164200 223116 164206 223128
rect 165246 223116 165252 223128
rect 165304 223116 165310 223168
rect 165798 223116 165804 223168
rect 165856 223156 165862 223168
rect 222286 223156 222292 223168
rect 165856 223128 222292 223156
rect 165856 223116 165862 223128
rect 222286 223116 222292 223128
rect 222344 223116 222350 223168
rect 224218 223116 224224 223168
rect 224276 223156 224282 223168
rect 238386 223156 238392 223168
rect 224276 223128 238392 223156
rect 224276 223116 224282 223128
rect 238386 223116 238392 223128
rect 238444 223116 238450 223168
rect 245286 223116 245292 223168
rect 245344 223156 245350 223168
rect 287606 223156 287612 223168
rect 245344 223128 287612 223156
rect 245344 223116 245350 223128
rect 287606 223116 287612 223128
rect 287664 223116 287670 223168
rect 290826 223116 290832 223168
rect 290884 223156 290890 223168
rect 323670 223156 323676 223168
rect 290884 223128 323676 223156
rect 290884 223116 290890 223128
rect 323670 223116 323676 223128
rect 323728 223116 323734 223168
rect 330478 223116 330484 223168
rect 330536 223156 330542 223168
rect 354950 223156 354956 223168
rect 330536 223128 354956 223156
rect 330536 223116 330542 223128
rect 354950 223116 354956 223128
rect 355008 223116 355014 223168
rect 357066 223116 357072 223168
rect 357124 223156 357130 223168
rect 376202 223156 376208 223168
rect 357124 223128 376208 223156
rect 357124 223116 357130 223128
rect 376202 223116 376208 223128
rect 376260 223116 376266 223168
rect 490190 223116 490196 223168
rect 490248 223156 490254 223168
rect 505646 223156 505652 223168
rect 490248 223128 505652 223156
rect 490248 223116 490254 223128
rect 505646 223116 505652 223128
rect 505704 223116 505710 223168
rect 513098 223116 513104 223168
rect 513156 223156 513162 223168
rect 534166 223156 534172 223168
rect 513156 223128 534172 223156
rect 513156 223116 513162 223128
rect 534166 223116 534172 223128
rect 534224 223116 534230 223168
rect 534718 223116 534724 223168
rect 534776 223156 534782 223168
rect 547414 223156 547420 223168
rect 534776 223128 547420 223156
rect 534776 223116 534782 223128
rect 547414 223116 547420 223128
rect 547472 223116 547478 223168
rect 89438 222980 89444 223032
rect 89496 223020 89502 223032
rect 161934 223020 161940 223032
rect 89496 222992 161940 223020
rect 89496 222980 89502 222992
rect 161934 222980 161940 222992
rect 161992 222980 161998 223032
rect 180886 223020 180892 223032
rect 162136 222992 180892 223020
rect 112806 222844 112812 222896
rect 112864 222884 112870 222896
rect 162136 222884 162164 222992
rect 180886 222980 180892 222992
rect 180944 222980 180950 223032
rect 181438 222980 181444 223032
rect 181496 223020 181502 223032
rect 234798 223020 234804 223032
rect 181496 222992 234804 223020
rect 181496 222980 181502 222992
rect 234798 222980 234804 222992
rect 234856 222980 234862 223032
rect 235166 222980 235172 223032
rect 235224 223020 235230 223032
rect 243262 223020 243268 223032
rect 235224 222992 243268 223020
rect 235224 222980 235230 222992
rect 243262 222980 243268 222992
rect 243320 222980 243326 223032
rect 250898 222980 250904 223032
rect 250956 223020 250962 223032
rect 294414 223020 294420 223032
rect 250956 222992 294420 223020
rect 250956 222980 250962 222992
rect 294414 222980 294420 222992
rect 294472 222980 294478 223032
rect 300302 222980 300308 223032
rect 300360 223020 300366 223032
rect 331766 223020 331772 223032
rect 300360 222992 331772 223020
rect 300360 222980 300366 222992
rect 331766 222980 331772 222992
rect 331824 222980 331830 223032
rect 337930 222980 337936 223032
rect 337988 223020 337994 223032
rect 359182 223020 359188 223032
rect 337988 222992 359188 223020
rect 337988 222980 337994 222992
rect 359182 222980 359188 222992
rect 359240 222980 359246 223032
rect 370498 222980 370504 223032
rect 370556 223020 370562 223032
rect 384574 223020 384580 223032
rect 370556 222992 384580 223020
rect 370556 222980 370562 222992
rect 384574 222980 384580 222992
rect 384632 222980 384638 223032
rect 387702 222980 387708 223032
rect 387760 223020 387766 223032
rect 398098 223020 398104 223032
rect 387760 222992 398104 223020
rect 387760 222980 387766 222992
rect 398098 222980 398104 222992
rect 398156 222980 398162 223032
rect 501138 222980 501144 223032
rect 501196 223020 501202 223032
rect 519262 223020 519268 223032
rect 501196 222992 519268 223020
rect 501196 222980 501202 222992
rect 519262 222980 519268 222992
rect 519320 222980 519326 223032
rect 523678 222980 523684 223032
rect 523736 223020 523742 223032
rect 548058 223020 548064 223032
rect 523736 222992 548064 223020
rect 523736 222980 523742 222992
rect 548058 222980 548064 222992
rect 548116 222980 548122 223032
rect 549254 222980 549260 223032
rect 549312 223020 549318 223032
rect 564802 223020 564808 223032
rect 549312 222992 564808 223020
rect 549312 222980 549318 222992
rect 564802 222980 564808 222992
rect 564860 222980 564866 223032
rect 112864 222856 162164 222884
rect 112864 222844 112870 222856
rect 162302 222844 162308 222896
rect 162360 222884 162366 222896
rect 221642 222884 221648 222896
rect 162360 222856 221648 222884
rect 162360 222844 162366 222856
rect 221642 222844 221648 222856
rect 221700 222844 221706 222896
rect 233142 222844 233148 222896
rect 233200 222884 233206 222896
rect 277670 222884 277676 222896
rect 233200 222856 277676 222884
rect 233200 222844 233206 222856
rect 277670 222844 277676 222856
rect 277728 222844 277734 222896
rect 283374 222844 283380 222896
rect 283432 222884 283438 222896
rect 316954 222884 316960 222896
rect 283432 222856 316960 222884
rect 283432 222844 283438 222856
rect 316954 222844 316960 222856
rect 317012 222844 317018 222896
rect 317138 222844 317144 222896
rect 317196 222884 317202 222896
rect 343358 222884 343364 222896
rect 317196 222856 343364 222884
rect 317196 222844 317202 222856
rect 343358 222844 343364 222856
rect 343416 222844 343422 222896
rect 347590 222844 347596 222896
rect 347648 222884 347654 222896
rect 368474 222884 368480 222896
rect 347648 222856 368480 222884
rect 347648 222844 347654 222856
rect 368474 222844 368480 222856
rect 368532 222844 368538 222896
rect 375098 222844 375104 222896
rect 375156 222884 375162 222896
rect 391014 222884 391020 222896
rect 375156 222856 391020 222884
rect 375156 222844 375162 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 397362 222844 397368 222896
rect 397420 222884 397426 222896
rect 407114 222884 407120 222896
rect 397420 222856 407120 222884
rect 397420 222844 397426 222856
rect 407114 222844 407120 222856
rect 407172 222844 407178 222896
rect 408402 222844 408408 222896
rect 408460 222884 408466 222896
rect 416866 222884 416872 222896
rect 408460 222856 416872 222884
rect 408460 222844 408466 222856
rect 416866 222844 416872 222856
rect 416924 222844 416930 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 478322 222844 478328 222896
rect 478380 222884 478386 222896
rect 486142 222884 486148 222896
rect 478380 222856 486148 222884
rect 478380 222844 478386 222856
rect 486142 222844 486148 222856
rect 486200 222844 486206 222896
rect 486970 222844 486976 222896
rect 487028 222884 487034 222896
rect 501046 222884 501052 222896
rect 487028 222856 501052 222884
rect 487028 222844 487034 222856
rect 501046 222844 501052 222856
rect 501104 222844 501110 222896
rect 504634 222844 504640 222896
rect 504692 222884 504698 222896
rect 523402 222884 523408 222896
rect 504692 222856 523408 222884
rect 504692 222844 504698 222856
rect 523402 222844 523408 222856
rect 523460 222844 523466 222896
rect 533706 222844 533712 222896
rect 533764 222884 533770 222896
rect 560754 222884 560760 222896
rect 533764 222856 560760 222884
rect 533764 222844 533770 222856
rect 560754 222844 560760 222856
rect 560812 222884 560818 222896
rect 562962 222884 562968 222896
rect 560812 222856 562968 222884
rect 560812 222844 560818 222856
rect 562962 222844 562968 222856
rect 563020 222844 563026 222896
rect 564618 222776 564624 222828
rect 564676 222816 564682 222828
rect 569310 222816 569316 222828
rect 564676 222788 569316 222816
rect 564676 222776 564682 222788
rect 569310 222776 569316 222788
rect 569368 222776 569374 222828
rect 85482 222708 85488 222760
rect 85540 222748 85546 222760
rect 161750 222748 161756 222760
rect 85540 222720 161756 222748
rect 85540 222708 85546 222720
rect 161750 222708 161756 222720
rect 161808 222708 161814 222760
rect 162118 222708 162124 222760
rect 162176 222748 162182 222760
rect 162176 222720 175964 222748
rect 162176 222708 162182 222720
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 175550 222612 175556 222624
rect 99340 222584 175556 222612
rect 99340 222572 99346 222584
rect 175550 222572 175556 222584
rect 175608 222572 175614 222624
rect 175936 222612 175964 222720
rect 176102 222708 176108 222760
rect 176160 222748 176166 222760
rect 181622 222748 181628 222760
rect 176160 222720 181628 222748
rect 176160 222708 176166 222720
rect 181622 222708 181628 222720
rect 181680 222708 181686 222760
rect 192110 222708 192116 222760
rect 192168 222748 192174 222760
rect 207474 222748 207480 222760
rect 192168 222720 207480 222748
rect 192168 222708 192174 222720
rect 207474 222708 207480 222720
rect 207532 222708 207538 222760
rect 209498 222708 209504 222760
rect 209556 222748 209562 222760
rect 210234 222748 210240 222760
rect 209556 222720 210240 222748
rect 209556 222708 209562 222720
rect 210234 222708 210240 222720
rect 210292 222708 210298 222760
rect 213822 222708 213828 222760
rect 213880 222748 213886 222760
rect 262858 222748 262864 222760
rect 213880 222720 262864 222748
rect 213880 222708 213886 222720
rect 262858 222708 262864 222720
rect 262916 222708 262922 222760
rect 263502 222708 263508 222760
rect 263560 222748 263566 222760
rect 296990 222748 296996 222760
rect 263560 222720 296996 222748
rect 263560 222708 263566 222720
rect 296990 222708 296996 222720
rect 297048 222708 297054 222760
rect 564802 222640 564808 222692
rect 564860 222680 564866 222692
rect 572162 222680 572168 222692
rect 564860 222652 572168 222680
rect 564860 222640 564866 222652
rect 572162 222640 572168 222652
rect 572220 222640 572226 222692
rect 175936 222584 214604 222612
rect 133506 222436 133512 222488
rect 133564 222476 133570 222488
rect 151354 222476 151360 222488
rect 133564 222448 151360 222476
rect 133564 222436 133570 222448
rect 151354 222436 151360 222448
rect 151412 222436 151418 222488
rect 154206 222436 154212 222488
rect 154264 222476 154270 222488
rect 214374 222476 214380 222488
rect 154264 222448 214380 222476
rect 154264 222436 154270 222448
rect 214374 222436 214380 222448
rect 214432 222436 214438 222488
rect 214576 222476 214604 222584
rect 214742 222572 214748 222624
rect 214800 222612 214806 222624
rect 260282 222612 260288 222624
rect 214800 222584 260288 222612
rect 214800 222572 214806 222584
rect 260282 222572 260288 222584
rect 260340 222572 260346 222624
rect 562410 222504 562416 222556
rect 562468 222544 562474 222556
rect 569126 222544 569132 222556
rect 562468 222516 569132 222544
rect 562468 222504 562474 222516
rect 569126 222504 569132 222516
rect 569184 222504 569190 222556
rect 219710 222476 219716 222488
rect 214576 222448 219716 222476
rect 219710 222436 219716 222448
rect 219768 222436 219774 222488
rect 220078 222436 220084 222488
rect 220136 222476 220142 222488
rect 268654 222476 268660 222488
rect 220136 222448 268660 222476
rect 220136 222436 220142 222448
rect 268654 222436 268660 222448
rect 268712 222436 268718 222488
rect 557350 222368 557356 222420
rect 557408 222408 557414 222420
rect 562778 222408 562784 222420
rect 557408 222380 562784 222408
rect 557408 222368 557414 222380
rect 562778 222368 562784 222380
rect 562836 222368 562842 222420
rect 563422 222368 563428 222420
rect 563480 222408 563486 222420
rect 571426 222408 571432 222420
rect 563480 222380 571432 222408
rect 563480 222368 563486 222380
rect 571426 222368 571432 222380
rect 571484 222368 571490 222420
rect 572346 222368 572352 222420
rect 572404 222408 572410 222420
rect 573174 222408 573180 222420
rect 572404 222380 573180 222408
rect 572404 222368 572410 222380
rect 573174 222368 573180 222380
rect 573232 222368 573238 222420
rect 56502 222300 56508 222352
rect 56560 222340 56566 222352
rect 142614 222340 142620 222352
rect 56560 222312 142620 222340
rect 56560 222300 56566 222312
rect 142614 222300 142620 222312
rect 142672 222300 142678 222352
rect 145006 222300 145012 222352
rect 145064 222340 145070 222352
rect 208762 222340 208768 222352
rect 145064 222312 208768 222340
rect 145064 222300 145070 222312
rect 208762 222300 208768 222312
rect 208820 222300 208826 222352
rect 210970 222300 210976 222352
rect 211028 222340 211034 222352
rect 214742 222340 214748 222352
rect 211028 222312 214748 222340
rect 211028 222300 211034 222312
rect 214742 222300 214748 222312
rect 214800 222300 214806 222352
rect 220446 222300 220452 222352
rect 220504 222340 220510 222352
rect 268010 222340 268016 222352
rect 220504 222312 268016 222340
rect 220504 222300 220510 222312
rect 268010 222300 268016 222312
rect 268068 222300 268074 222352
rect 143442 222232 143448 222284
rect 143500 222272 143506 222284
rect 144822 222272 144828 222284
rect 143500 222244 144828 222272
rect 143500 222232 143506 222244
rect 144822 222232 144828 222244
rect 144880 222232 144886 222284
rect 214926 222232 214932 222284
rect 214984 222272 214990 222284
rect 216214 222272 216220 222284
rect 214984 222244 216220 222272
rect 214984 222232 214990 222244
rect 216214 222232 216220 222244
rect 216272 222232 216278 222284
rect 593966 222272 593972 222284
rect 543706 222244 593972 222272
rect 171244 222176 171456 222204
rect 117774 222136 117780 222148
rect 103486 222108 117780 222136
rect 95418 221960 95424 222012
rect 95476 222000 95482 222012
rect 103486 222000 103514 222108
rect 117774 222096 117780 222108
rect 117832 222096 117838 222148
rect 117958 222096 117964 222148
rect 118016 222136 118022 222148
rect 171042 222136 171048 222148
rect 118016 222108 171048 222136
rect 118016 222096 118022 222108
rect 171042 222096 171048 222108
rect 171100 222096 171106 222148
rect 95476 221972 103514 222000
rect 95476 221960 95482 221972
rect 104526 221960 104532 222012
rect 104584 222000 104590 222012
rect 171244 222000 171272 222176
rect 171428 222136 171456 222176
rect 173084 222176 173204 222204
rect 173084 222136 173112 222176
rect 171428 222108 173112 222136
rect 173176 222068 173204 222176
rect 174906 222164 174912 222216
rect 174964 222204 174970 222216
rect 176286 222204 176292 222216
rect 174964 222176 176292 222204
rect 174964 222164 174970 222176
rect 176286 222164 176292 222176
rect 176344 222164 176350 222216
rect 180886 222164 180892 222216
rect 180944 222204 180950 222216
rect 185210 222204 185216 222216
rect 180944 222176 185216 222204
rect 180944 222164 180950 222176
rect 185210 222164 185216 222176
rect 185268 222164 185274 222216
rect 482922 222164 482928 222216
rect 482980 222204 482986 222216
rect 543706 222204 543734 222244
rect 593966 222232 593972 222244
rect 594024 222232 594030 222284
rect 482980 222176 543734 222204
rect 482980 222164 482986 222176
rect 176654 222096 176660 222148
rect 176712 222136 176718 222148
rect 179966 222136 179972 222148
rect 176712 222108 179972 222136
rect 176712 222096 176718 222108
rect 179966 222096 179972 222108
rect 180024 222096 180030 222148
rect 240134 222136 240140 222148
rect 185412 222108 240140 222136
rect 176102 222068 176108 222080
rect 173176 222040 176108 222068
rect 176102 222028 176108 222040
rect 176160 222028 176166 222080
rect 181622 222028 181628 222080
rect 181680 222068 181686 222080
rect 185412 222068 185440 222108
rect 240134 222096 240140 222108
rect 240192 222096 240198 222148
rect 261018 222096 261024 222148
rect 261076 222136 261082 222148
rect 301682 222136 301688 222148
rect 261076 222108 301688 222136
rect 261076 222096 261082 222108
rect 301682 222096 301688 222108
rect 301740 222096 301746 222148
rect 311526 222096 311532 222148
rect 311584 222136 311590 222148
rect 338390 222136 338396 222148
rect 311584 222108 338396 222136
rect 311584 222096 311590 222108
rect 338390 222096 338396 222108
rect 338448 222096 338454 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 553210 222096 553216 222148
rect 553268 222136 553274 222148
rect 558178 222136 558184 222148
rect 553268 222108 558184 222136
rect 553268 222096 553274 222108
rect 558178 222096 558184 222108
rect 558236 222096 558242 222148
rect 558362 222096 558368 222148
rect 558420 222136 558426 222148
rect 562410 222136 562416 222148
rect 558420 222108 562416 222136
rect 558420 222096 558426 222108
rect 562410 222096 562416 222108
rect 562468 222096 562474 222148
rect 562962 222096 562968 222148
rect 563020 222136 563026 222148
rect 567562 222136 567568 222148
rect 563020 222108 567568 222136
rect 563020 222096 563026 222108
rect 567562 222096 567568 222108
rect 567620 222096 567626 222148
rect 567746 222096 567752 222148
rect 567804 222136 567810 222148
rect 572346 222136 572352 222148
rect 567804 222108 572352 222136
rect 567804 222096 567810 222108
rect 572346 222096 572352 222108
rect 572404 222096 572410 222148
rect 572622 222096 572628 222148
rect 572680 222136 572686 222148
rect 572680 222108 600820 222136
rect 572680 222096 572686 222108
rect 181680 222040 185440 222068
rect 181680 222028 181686 222040
rect 172974 222000 172980 222012
rect 104584 221972 171272 222000
rect 171336 221972 172980 222000
rect 104584 221960 104590 221972
rect 71406 221824 71412 221876
rect 71464 221864 71470 221876
rect 142798 221864 142804 221876
rect 71464 221836 142804 221864
rect 71464 221824 71470 221836
rect 142798 221824 142804 221836
rect 142856 221824 142862 221876
rect 142982 221824 142988 221876
rect 143040 221864 143046 221876
rect 171336 221864 171364 221972
rect 172974 221960 172980 221972
rect 173032 221960 173038 222012
rect 176286 221960 176292 222012
rect 176344 222000 176350 222012
rect 181438 222000 181444 222012
rect 176344 221972 181444 222000
rect 176344 221960 176350 221972
rect 181438 221960 181444 221972
rect 181496 221960 181502 222012
rect 185854 221960 185860 222012
rect 185912 222000 185918 222012
rect 237558 222000 237564 222012
rect 185912 221972 237564 222000
rect 185912 221960 185918 221972
rect 237558 221960 237564 221972
rect 237616 221960 237622 222012
rect 243630 221960 243636 222012
rect 243688 222000 243694 222012
rect 285950 222000 285956 222012
rect 243688 221972 285956 222000
rect 243688 221960 243694 221972
rect 285950 221960 285956 221972
rect 286008 221960 286014 222012
rect 309870 221960 309876 222012
rect 309928 222000 309934 222012
rect 338206 222000 338212 222012
rect 309928 221972 338212 222000
rect 309928 221960 309934 221972
rect 338206 221960 338212 221972
rect 338264 221960 338270 222012
rect 500034 221960 500040 222012
rect 500092 222000 500098 222012
rect 518434 222000 518440 222012
rect 500092 221972 518440 222000
rect 500092 221960 500098 221972
rect 518434 221960 518440 221972
rect 518492 221960 518498 222012
rect 525886 221960 525892 222012
rect 525944 222000 525950 222012
rect 597462 222000 597468 222012
rect 525944 221972 597468 222000
rect 525944 221960 525950 221972
rect 597462 221960 597468 221972
rect 597520 221960 597526 222012
rect 600590 222000 600596 222012
rect 597664 221972 600596 222000
rect 340874 221892 340880 221944
rect 340932 221932 340938 221944
rect 341610 221932 341616 221944
rect 340932 221904 341616 221932
rect 340932 221892 340938 221904
rect 341610 221892 341616 221904
rect 341668 221892 341674 221944
rect 143040 221836 171364 221864
rect 143040 221824 143046 221836
rect 171502 221824 171508 221876
rect 171560 221864 171566 221876
rect 229646 221864 229652 221876
rect 171560 221836 229652 221864
rect 171560 221824 171566 221836
rect 229646 221824 229652 221836
rect 229704 221824 229710 221876
rect 230382 221824 230388 221876
rect 230440 221864 230446 221876
rect 258718 221864 258724 221876
rect 230440 221836 258724 221864
rect 230440 221824 230446 221836
rect 258718 221824 258724 221836
rect 258776 221824 258782 221876
rect 267826 221824 267832 221876
rect 267884 221864 267890 221876
rect 273990 221864 273996 221876
rect 267884 221836 273996 221864
rect 267884 221824 267890 221836
rect 273990 221824 273996 221836
rect 274048 221824 274054 221876
rect 285674 221824 285680 221876
rect 285732 221864 285738 221876
rect 286318 221864 286324 221876
rect 285732 221836 286324 221864
rect 285732 221824 285738 221836
rect 286318 221824 286324 221836
rect 286376 221824 286382 221876
rect 304626 221824 304632 221876
rect 304684 221864 304690 221876
rect 334066 221864 334072 221876
rect 304684 221836 334072 221864
rect 304684 221824 304690 221836
rect 334066 221824 334072 221836
rect 334124 221824 334130 221876
rect 515398 221824 515404 221876
rect 515456 221864 515462 221876
rect 534994 221864 535000 221876
rect 515456 221836 535000 221864
rect 515456 221824 515462 221836
rect 534994 221824 535000 221836
rect 535052 221824 535058 221876
rect 542722 221824 542728 221876
rect 542780 221864 542786 221876
rect 543182 221864 543188 221876
rect 542780 221836 543188 221864
rect 542780 221824 542786 221836
rect 543182 221824 543188 221836
rect 543240 221864 543246 221876
rect 597664 221864 597692 221972
rect 600590 221960 600596 221972
rect 600648 221960 600654 222012
rect 600792 222000 600820 222108
rect 600958 222096 600964 222148
rect 601016 222136 601022 222148
rect 607766 222136 607772 222148
rect 601016 222108 607772 222136
rect 601016 222096 601022 222108
rect 607766 222096 607772 222108
rect 607824 222096 607830 222148
rect 601142 222000 601148 222012
rect 600792 221972 601148 222000
rect 601142 221960 601148 221972
rect 601200 221960 601206 222012
rect 543240 221836 597692 221864
rect 543240 221824 543246 221836
rect 597830 221824 597836 221876
rect 597888 221864 597894 221876
rect 607306 221864 607312 221876
rect 597888 221836 607312 221864
rect 597888 221824 597894 221836
rect 607306 221824 607312 221836
rect 607364 221824 607370 221876
rect 68094 221688 68100 221740
rect 68152 221728 68158 221740
rect 147490 221728 147496 221740
rect 68152 221700 147496 221728
rect 68152 221688 68158 221700
rect 147490 221688 147496 221700
rect 147548 221688 147554 221740
rect 147766 221688 147772 221740
rect 147824 221728 147830 221740
rect 147824 221700 157334 221728
rect 147824 221688 147830 221700
rect 61470 221552 61476 221604
rect 61528 221592 61534 221604
rect 137278 221592 137284 221604
rect 61528 221564 137284 221592
rect 61528 221552 61534 221564
rect 137278 221552 137284 221564
rect 137336 221552 137342 221604
rect 137462 221552 137468 221604
rect 137520 221592 137526 221604
rect 137520 221564 142660 221592
rect 137520 221552 137526 221564
rect 64598 221416 64604 221468
rect 64656 221456 64662 221468
rect 138290 221456 138296 221468
rect 64656 221428 138296 221456
rect 64656 221416 64662 221428
rect 138290 221416 138296 221428
rect 138348 221416 138354 221468
rect 138474 221416 138480 221468
rect 138532 221456 138538 221468
rect 142430 221456 142436 221468
rect 138532 221428 142436 221456
rect 138532 221416 138538 221428
rect 142430 221416 142436 221428
rect 142488 221416 142494 221468
rect 142632 221456 142660 221564
rect 142798 221552 142804 221604
rect 142856 221592 142862 221604
rect 147306 221592 147312 221604
rect 142856 221564 147312 221592
rect 142856 221552 142862 221564
rect 147306 221552 147312 221564
rect 147364 221552 147370 221604
rect 157306 221592 157334 221700
rect 161658 221688 161664 221740
rect 161716 221728 161722 221740
rect 224402 221728 224408 221740
rect 161716 221700 224408 221728
rect 161716 221688 161722 221700
rect 224402 221688 224408 221700
rect 224460 221688 224466 221740
rect 227070 221688 227076 221740
rect 227128 221728 227134 221740
rect 272702 221728 272708 221740
rect 227128 221700 272708 221728
rect 227128 221688 227134 221700
rect 272702 221688 272708 221700
rect 272760 221688 272766 221740
rect 275278 221728 275284 221740
rect 272904 221700 275284 221728
rect 204898 221592 204904 221604
rect 157306 221564 204904 221592
rect 204898 221552 204904 221564
rect 204956 221552 204962 221604
rect 205082 221552 205088 221604
rect 205140 221592 205146 221604
rect 205140 221564 212304 221592
rect 205140 221552 205146 221564
rect 142982 221456 142988 221468
rect 142632 221428 142988 221456
rect 142982 221416 142988 221428
rect 143040 221416 143046 221468
rect 148410 221416 148416 221468
rect 148468 221456 148474 221468
rect 211982 221456 211988 221468
rect 148468 221428 211988 221456
rect 148468 221416 148474 221428
rect 211982 221416 211988 221428
rect 212040 221416 212046 221468
rect 212276 221456 212304 221564
rect 214650 221552 214656 221604
rect 214708 221592 214714 221604
rect 258534 221592 258540 221604
rect 214708 221564 258540 221592
rect 214708 221552 214714 221564
rect 258534 221552 258540 221564
rect 258592 221552 258598 221604
rect 258718 221552 258724 221604
rect 258776 221592 258782 221604
rect 272904 221592 272932 221700
rect 275278 221688 275284 221700
rect 275336 221688 275342 221740
rect 278314 221688 278320 221740
rect 278372 221728 278378 221740
rect 313458 221728 313464 221740
rect 278372 221700 313464 221728
rect 278372 221688 278378 221700
rect 313458 221688 313464 221700
rect 313516 221688 313522 221740
rect 331398 221688 331404 221740
rect 331456 221728 331462 221740
rect 353938 221728 353944 221740
rect 331456 221700 353944 221728
rect 331456 221688 331462 221700
rect 353938 221688 353944 221700
rect 353996 221688 354002 221740
rect 359550 221688 359556 221740
rect 359608 221728 359614 221740
rect 376846 221728 376852 221740
rect 359608 221700 376852 221728
rect 359608 221688 359614 221700
rect 376846 221688 376852 221700
rect 376904 221688 376910 221740
rect 484302 221688 484308 221740
rect 484360 221728 484366 221740
rect 496078 221728 496084 221740
rect 484360 221700 496084 221728
rect 484360 221688 484366 221700
rect 496078 221688 496084 221700
rect 496136 221688 496142 221740
rect 503438 221688 503444 221740
rect 503496 221728 503502 221740
rect 521746 221728 521752 221740
rect 503496 221700 521752 221728
rect 503496 221688 503502 221700
rect 521746 221688 521752 221700
rect 521804 221688 521810 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 546586 221728 546592 221740
rect 522908 221700 546592 221728
rect 522908 221688 522914 221700
rect 546586 221688 546592 221700
rect 546644 221688 546650 221740
rect 547138 221688 547144 221740
rect 547196 221728 547202 221740
rect 547196 221700 555924 221728
rect 547196 221688 547202 221700
rect 258776 221564 272932 221592
rect 258776 221552 258782 221564
rect 275094 221552 275100 221604
rect 275152 221592 275158 221604
rect 310882 221592 310888 221604
rect 275152 221564 310888 221592
rect 275152 221552 275158 221564
rect 310882 221552 310888 221564
rect 310940 221552 310946 221604
rect 314562 221552 314568 221604
rect 314620 221592 314626 221604
rect 340874 221592 340880 221604
rect 314620 221564 340880 221592
rect 314620 221552 314626 221564
rect 340874 221552 340880 221564
rect 340932 221552 340938 221604
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361942 221592 361948 221604
rect 341392 221564 361948 221592
rect 341392 221552 341398 221564
rect 361942 221552 361948 221564
rect 362000 221552 362006 221604
rect 377766 221552 377772 221604
rect 377824 221592 377830 221604
rect 390002 221592 390008 221604
rect 377824 221564 390008 221592
rect 377824 221552 377830 221564
rect 390002 221552 390008 221564
rect 390060 221552 390066 221604
rect 456702 221552 456708 221604
rect 456760 221592 456766 221604
rect 462130 221592 462136 221604
rect 456760 221564 462136 221592
rect 456760 221552 456766 221564
rect 462130 221552 462136 221564
rect 462188 221552 462194 221604
rect 496262 221552 496268 221604
rect 496320 221592 496326 221604
rect 513374 221592 513380 221604
rect 496320 221564 513380 221592
rect 496320 221552 496326 221564
rect 513374 221552 513380 221564
rect 513432 221552 513438 221604
rect 529750 221552 529756 221604
rect 529808 221592 529814 221604
rect 555418 221592 555424 221604
rect 529808 221564 555424 221592
rect 529808 221552 529814 221564
rect 555418 221552 555424 221564
rect 555476 221552 555482 221604
rect 555896 221592 555924 221700
rect 556062 221688 556068 221740
rect 556120 221728 556126 221740
rect 562962 221728 562968 221740
rect 556120 221700 562968 221728
rect 556120 221688 556126 221700
rect 562962 221688 562968 221700
rect 563020 221688 563026 221740
rect 563790 221688 563796 221740
rect 563848 221728 563854 221740
rect 567378 221728 567384 221740
rect 563848 221700 567384 221728
rect 563848 221688 563854 221700
rect 567378 221688 567384 221700
rect 567436 221688 567442 221740
rect 567562 221688 567568 221740
rect 567620 221728 567626 221740
rect 567620 221700 601004 221728
rect 567620 221688 567626 221700
rect 556338 221592 556344 221604
rect 555896 221564 556344 221592
rect 556338 221552 556344 221564
rect 556396 221552 556402 221604
rect 556798 221552 556804 221604
rect 556856 221592 556862 221604
rect 567470 221592 567476 221604
rect 556856 221564 567476 221592
rect 556856 221552 556862 221564
rect 567470 221552 567476 221564
rect 567528 221592 567534 221604
rect 567746 221592 567752 221604
rect 567528 221564 567752 221592
rect 567528 221552 567534 221564
rect 567746 221552 567752 221564
rect 567804 221552 567810 221604
rect 568114 221552 568120 221604
rect 568172 221592 568178 221604
rect 597830 221592 597836 221604
rect 568172 221564 597836 221592
rect 568172 221552 568178 221564
rect 597830 221552 597836 221564
rect 597888 221552 597894 221604
rect 600976 221592 601004 221700
rect 601326 221688 601332 221740
rect 601384 221728 601390 221740
rect 606570 221728 606576 221740
rect 601384 221700 606576 221728
rect 601384 221688 601390 221700
rect 606570 221688 606576 221700
rect 606628 221688 606634 221740
rect 610250 221592 610256 221604
rect 600976 221564 610256 221592
rect 610250 221552 610256 221564
rect 610308 221552 610314 221604
rect 655698 221552 655704 221604
rect 655756 221592 655762 221604
rect 659562 221592 659568 221604
rect 655756 221564 659568 221592
rect 655756 221552 655762 221564
rect 659562 221552 659568 221564
rect 659620 221552 659626 221604
rect 232130 221456 232136 221468
rect 212276 221428 232136 221456
rect 232130 221416 232136 221428
rect 232188 221416 232194 221468
rect 241146 221416 241152 221468
rect 241204 221456 241210 221468
rect 285674 221456 285680 221468
rect 241204 221428 285680 221456
rect 241204 221416 241210 221428
rect 285674 221416 285680 221428
rect 285732 221416 285738 221468
rect 285950 221416 285956 221468
rect 286008 221456 286014 221468
rect 289814 221456 289820 221468
rect 286008 221428 289820 221456
rect 286008 221416 286014 221428
rect 289814 221416 289820 221428
rect 289872 221416 289878 221468
rect 289998 221416 290004 221468
rect 290056 221456 290062 221468
rect 321738 221456 321744 221468
rect 290056 221428 321744 221456
rect 290056 221416 290062 221428
rect 321738 221416 321744 221428
rect 321796 221416 321802 221468
rect 338850 221416 338856 221468
rect 338908 221456 338914 221468
rect 338908 221428 354674 221456
rect 338908 221416 338914 221428
rect 117774 221280 117780 221332
rect 117832 221320 117838 221332
rect 117832 221292 118188 221320
rect 117832 221280 117838 221292
rect 107838 221144 107844 221196
rect 107896 221184 107902 221196
rect 117958 221184 117964 221196
rect 107896 221156 117964 221184
rect 107896 221144 107902 221156
rect 117958 221144 117964 221156
rect 118016 221144 118022 221196
rect 118160 221184 118188 221292
rect 118418 221280 118424 221332
rect 118476 221320 118482 221332
rect 177390 221320 177396 221332
rect 118476 221292 177396 221320
rect 118476 221280 118482 221292
rect 177390 221280 177396 221292
rect 177448 221280 177454 221332
rect 178218 221280 178224 221332
rect 178276 221320 178282 221332
rect 181254 221320 181260 221332
rect 178276 221292 181260 221320
rect 178276 221280 178282 221292
rect 181254 221280 181260 221292
rect 181312 221280 181318 221332
rect 181438 221280 181444 221332
rect 181496 221320 181502 221332
rect 195238 221320 195244 221332
rect 181496 221292 195244 221320
rect 181496 221280 181502 221292
rect 195238 221280 195244 221292
rect 195296 221280 195302 221332
rect 195422 221280 195428 221332
rect 195480 221320 195486 221332
rect 245102 221320 245108 221332
rect 195480 221292 245108 221320
rect 195480 221280 195486 221292
rect 245102 221280 245108 221292
rect 245160 221280 245166 221332
rect 258534 221280 258540 221332
rect 258592 221320 258598 221332
rect 265710 221320 265716 221332
rect 258592 221292 265716 221320
rect 258592 221280 258598 221292
rect 265710 221280 265716 221292
rect 265768 221280 265774 221332
rect 273438 221280 273444 221332
rect 273496 221320 273502 221332
rect 309226 221320 309232 221332
rect 273496 221292 309232 221320
rect 273496 221280 273502 221292
rect 309226 221280 309232 221292
rect 309284 221280 309290 221332
rect 354646 221320 354674 221428
rect 362034 221416 362040 221468
rect 362092 221456 362098 221468
rect 379882 221456 379888 221468
rect 362092 221428 379888 221456
rect 362092 221416 362098 221428
rect 379882 221416 379888 221428
rect 379940 221416 379946 221468
rect 391014 221416 391020 221468
rect 391072 221456 391078 221468
rect 400306 221456 400312 221468
rect 391072 221428 400312 221456
rect 391072 221416 391078 221428
rect 400306 221416 400312 221428
rect 400364 221416 400370 221468
rect 405090 221416 405096 221468
rect 405148 221456 405154 221468
rect 414198 221456 414204 221468
rect 405148 221428 414204 221456
rect 405148 221416 405154 221428
rect 414198 221416 414204 221428
rect 414256 221416 414262 221468
rect 452562 221416 452568 221468
rect 452620 221456 452626 221468
rect 456702 221456 456708 221468
rect 452620 221428 456708 221456
rect 452620 221416 452626 221428
rect 456702 221416 456708 221428
rect 456760 221416 456766 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538674 221456 538680 221468
rect 483808 221428 538680 221456
rect 483808 221416 483814 221428
rect 538674 221416 538680 221428
rect 538732 221416 538738 221468
rect 550634 221416 550640 221468
rect 550692 221456 550698 221468
rect 600958 221456 600964 221468
rect 550692 221428 600964 221456
rect 550692 221416 550698 221428
rect 600958 221416 600964 221428
rect 601016 221416 601022 221468
rect 601142 221416 601148 221468
rect 601200 221456 601206 221468
rect 610066 221456 610072 221468
rect 601200 221428 610072 221456
rect 601200 221416 601206 221428
rect 610066 221416 610072 221428
rect 610124 221416 610130 221468
rect 654134 221416 654140 221468
rect 654192 221456 654198 221468
rect 655882 221456 655888 221468
rect 654192 221428 655888 221456
rect 654192 221416 654198 221428
rect 655882 221416 655888 221428
rect 655940 221416 655946 221468
rect 362310 221320 362316 221332
rect 354646 221292 362316 221320
rect 362310 221280 362316 221292
rect 362368 221280 362374 221332
rect 548058 221212 548064 221264
rect 548116 221252 548122 221264
rect 567746 221252 567752 221264
rect 548116 221224 567752 221252
rect 548116 221212 548122 221224
rect 567746 221212 567752 221224
rect 567804 221212 567810 221264
rect 567930 221212 567936 221264
rect 567988 221252 567994 221264
rect 568942 221252 568948 221264
rect 567988 221224 568948 221252
rect 567988 221212 567994 221224
rect 568942 221212 568948 221224
rect 569000 221212 569006 221264
rect 569126 221212 569132 221264
rect 569184 221252 569190 221264
rect 608686 221252 608692 221264
rect 569184 221224 608692 221252
rect 569184 221212 569190 221224
rect 608686 221212 608692 221224
rect 608744 221212 608750 221264
rect 137094 221184 137100 221196
rect 118160 221156 137100 221184
rect 137094 221144 137100 221156
rect 137152 221144 137158 221196
rect 137278 221144 137284 221196
rect 137336 221184 137342 221196
rect 143994 221184 144000 221196
rect 137336 221156 144000 221184
rect 137336 221144 137342 221156
rect 143994 221144 144000 221156
rect 144052 221144 144058 221196
rect 144178 221144 144184 221196
rect 144236 221184 144242 221196
rect 203242 221184 203248 221196
rect 144236 221156 203248 221184
rect 144236 221144 144242 221156
rect 203242 221144 203248 221156
rect 203300 221144 203306 221196
rect 205082 221184 205088 221196
rect 204732 221156 205088 221184
rect 117774 221008 117780 221060
rect 117832 221048 117838 221060
rect 187878 221048 187884 221060
rect 117832 221020 187884 221048
rect 117832 221008 117838 221020
rect 187878 221008 187884 221020
rect 187936 221008 187942 221060
rect 188154 221008 188160 221060
rect 188212 221048 188218 221060
rect 195054 221048 195060 221060
rect 188212 221020 195060 221048
rect 188212 221008 188218 221020
rect 195054 221008 195060 221020
rect 195112 221008 195118 221060
rect 195238 221008 195244 221060
rect 195296 221048 195302 221060
rect 204732 221048 204760 221156
rect 205082 221144 205088 221156
rect 205140 221144 205146 221196
rect 206002 221144 206008 221196
rect 206060 221184 206066 221196
rect 258350 221184 258356 221196
rect 206060 221156 258356 221184
rect 206060 221144 206066 221156
rect 258350 221144 258356 221156
rect 258408 221144 258414 221196
rect 542078 221076 542084 221128
rect 542136 221116 542142 221128
rect 549254 221116 549260 221128
rect 542136 221088 549260 221116
rect 542136 221076 542142 221088
rect 549254 221076 549260 221088
rect 549312 221076 549318 221128
rect 550450 221076 550456 221128
rect 550508 221116 550514 221128
rect 554222 221116 554228 221128
rect 550508 221088 554228 221116
rect 550508 221076 550514 221088
rect 554222 221076 554228 221088
rect 554280 221076 554286 221128
rect 558178 221076 558184 221128
rect 558236 221116 558242 221128
rect 608870 221116 608876 221128
rect 558236 221088 608876 221116
rect 558236 221076 558242 221088
rect 608870 221076 608876 221088
rect 608928 221076 608934 221128
rect 195296 221020 204760 221048
rect 195296 221008 195302 221020
rect 204898 221008 204904 221060
rect 204956 221048 204962 221060
rect 211614 221048 211620 221060
rect 204956 221020 211620 221048
rect 204956 221008 204962 221020
rect 211614 221008 211620 221020
rect 211672 221008 211678 221060
rect 211982 221008 211988 221060
rect 212040 221048 212046 221060
rect 214190 221048 214196 221060
rect 212040 221020 214196 221048
rect 212040 221008 212046 221020
rect 214190 221008 214196 221020
rect 214248 221008 214254 221060
rect 237098 221008 237104 221060
rect 237156 221048 237162 221060
rect 280430 221048 280436 221060
rect 237156 221020 280436 221048
rect 237156 221008 237162 221020
rect 280430 221008 280436 221020
rect 280488 221008 280494 221060
rect 415026 221008 415032 221060
rect 415084 221048 415090 221060
rect 420178 221048 420184 221060
rect 415084 221020 420184 221048
rect 415084 221008 415090 221020
rect 420178 221008 420184 221020
rect 420236 221008 420242 221060
rect 545758 220940 545764 220992
rect 545816 220980 545822 220992
rect 601326 220980 601332 220992
rect 545816 220952 601332 220980
rect 545816 220940 545822 220952
rect 601326 220940 601332 220952
rect 601384 220940 601390 220992
rect 606018 220980 606024 220992
rect 601528 220952 606024 220980
rect 108022 220872 108028 220924
rect 108080 220912 108086 220924
rect 108080 220884 108528 220912
rect 108080 220872 108086 220884
rect 97718 220736 97724 220788
rect 97776 220776 97782 220788
rect 108500 220776 108528 220884
rect 114462 220872 114468 220924
rect 114520 220912 114526 220924
rect 118418 220912 118424 220924
rect 114520 220884 118424 220912
rect 114520 220872 114526 220884
rect 118418 220872 118424 220884
rect 118476 220872 118482 220924
rect 128538 220872 128544 220924
rect 128596 220912 128602 220924
rect 198918 220912 198924 220924
rect 128596 220884 198924 220912
rect 128596 220872 128602 220884
rect 198918 220872 198924 220884
rect 198976 220872 198982 220924
rect 203242 220872 203248 220924
rect 203300 220912 203306 220924
rect 206462 220912 206468 220924
rect 203300 220884 206468 220912
rect 203300 220872 203306 220884
rect 206462 220872 206468 220884
rect 206520 220872 206526 220924
rect 256050 220872 256056 220924
rect 256108 220912 256114 220924
rect 261386 220912 261392 220924
rect 256108 220884 261392 220912
rect 256108 220872 256114 220884
rect 261386 220872 261392 220884
rect 261444 220872 261450 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423766 220844 423772 220856
rect 420696 220816 423772 220844
rect 420696 220804 420702 220816
rect 423766 220804 423772 220816
rect 423824 220804 423830 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471698 220844 471704 220856
rect 466144 220816 471704 220844
rect 466144 220804 466150 220816
rect 471698 220804 471704 220816
rect 471756 220804 471762 220856
rect 518434 220804 518440 220856
rect 518492 220844 518498 220856
rect 600406 220844 600412 220856
rect 518492 220816 600412 220844
rect 518492 220804 518498 220816
rect 600406 220804 600412 220816
rect 600464 220804 600470 220856
rect 600590 220804 600596 220856
rect 600648 220844 600654 220856
rect 601528 220844 601556 220952
rect 606018 220940 606024 220952
rect 606076 220940 606082 220992
rect 600648 220816 601556 220844
rect 600648 220804 600654 220816
rect 137278 220776 137284 220788
rect 97776 220748 108252 220776
rect 108500 220748 137284 220776
rect 97776 220736 97782 220748
rect 108224 220708 108252 220748
rect 137278 220736 137284 220748
rect 137336 220736 137342 220788
rect 137462 220736 137468 220788
rect 137520 220776 137526 220788
rect 197722 220776 197728 220788
rect 137520 220748 197728 220776
rect 137520 220736 137526 220748
rect 197722 220736 197728 220748
rect 197780 220736 197786 220788
rect 198090 220736 198096 220788
rect 198148 220776 198154 220788
rect 252738 220776 252744 220788
rect 198148 220748 252744 220776
rect 198148 220736 198154 220748
rect 252738 220736 252744 220748
rect 252796 220736 252802 220788
rect 253566 220736 253572 220788
rect 253624 220776 253630 220788
rect 293310 220776 293316 220788
rect 253624 220748 293316 220776
rect 253624 220736 253630 220748
rect 293310 220736 293316 220748
rect 293368 220736 293374 220788
rect 296990 220736 296996 220788
rect 297048 220776 297054 220788
rect 310698 220776 310704 220788
rect 297048 220748 310704 220776
rect 297048 220736 297054 220748
rect 310698 220736 310704 220748
rect 310756 220736 310762 220788
rect 311802 220736 311808 220788
rect 311860 220776 311866 220788
rect 327074 220776 327080 220788
rect 311860 220748 327080 220776
rect 311860 220736 311866 220748
rect 327074 220736 327080 220748
rect 327132 220736 327138 220788
rect 329282 220736 329288 220788
rect 329340 220776 329346 220788
rect 331950 220776 331956 220788
rect 329340 220748 331956 220776
rect 329340 220736 329346 220748
rect 331950 220736 331956 220748
rect 332008 220736 332014 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418246 220776 418252 220788
rect 414256 220748 418252 220776
rect 414256 220736 414262 220748
rect 418246 220736 418252 220748
rect 418304 220736 418310 220788
rect 455230 220736 455236 220788
rect 455288 220776 455294 220788
rect 458818 220776 458824 220788
rect 455288 220748 458824 220776
rect 455288 220736 455294 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 475378 220736 475384 220788
rect 475436 220776 475442 220788
rect 476206 220776 476212 220788
rect 475436 220748 476212 220776
rect 475436 220736 475442 220748
rect 476206 220736 476212 220748
rect 476264 220736 476270 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 601970 220736 601976 220788
rect 602028 220776 602034 220788
rect 617242 220776 617248 220788
rect 602028 220748 617248 220776
rect 602028 220736 602034 220748
rect 617242 220736 617248 220748
rect 617300 220736 617306 220788
rect 108224 220680 108436 220708
rect 91278 220600 91284 220652
rect 91336 220640 91342 220652
rect 108022 220640 108028 220652
rect 91336 220612 108028 220640
rect 91336 220600 91342 220612
rect 108022 220600 108028 220612
rect 108080 220600 108086 220652
rect 108408 220640 108436 220680
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 172698 220640 172704 220652
rect 108408 220612 172704 220640
rect 172698 220600 172704 220612
rect 172756 220600 172762 220652
rect 177206 220600 177212 220652
rect 177264 220640 177270 220652
rect 182634 220640 182640 220652
rect 177264 220612 182640 220640
rect 177264 220600 177270 220612
rect 182634 220600 182640 220612
rect 182692 220600 182698 220652
rect 183094 220600 183100 220652
rect 183152 220640 183158 220652
rect 184198 220640 184204 220652
rect 183152 220612 184204 220640
rect 183152 220600 183158 220612
rect 184198 220600 184204 220612
rect 184256 220600 184262 220652
rect 184382 220600 184388 220652
rect 184440 220640 184446 220652
rect 234062 220640 234068 220652
rect 184440 220612 234068 220640
rect 184440 220600 184446 220612
rect 234062 220600 234068 220612
rect 234120 220600 234126 220652
rect 240318 220600 240324 220652
rect 240376 220640 240382 220652
rect 283006 220640 283012 220652
rect 240376 220612 283012 220640
rect 240376 220600 240382 220612
rect 283006 220600 283012 220612
rect 283064 220600 283070 220652
rect 296622 220600 296628 220652
rect 296680 220640 296686 220652
rect 327442 220640 327448 220652
rect 296680 220612 327448 220640
rect 296680 220600 296686 220612
rect 327442 220600 327448 220612
rect 327500 220600 327506 220652
rect 328086 220600 328092 220652
rect 328144 220640 328150 220652
rect 351362 220640 351368 220652
rect 328144 220612 351368 220640
rect 328144 220600 328150 220612
rect 351362 220600 351368 220612
rect 351420 220600 351426 220652
rect 473998 220600 474004 220652
rect 474056 220640 474062 220652
rect 475378 220640 475384 220652
rect 474056 220612 475384 220640
rect 474056 220600 474062 220612
rect 475378 220600 475384 220612
rect 475436 220600 475442 220652
rect 493962 220600 493968 220652
rect 494020 220640 494026 220652
rect 508498 220640 508504 220652
rect 494020 220612 508504 220640
rect 494020 220600 494026 220612
rect 508498 220600 508504 220612
rect 508556 220600 508562 220652
rect 511258 220600 511264 220652
rect 511316 220640 511322 220652
rect 527542 220640 527548 220652
rect 511316 220612 527548 220640
rect 511316 220600 511322 220612
rect 527542 220600 527548 220612
rect 527600 220600 527606 220652
rect 541710 220600 541716 220652
rect 541768 220640 541774 220652
rect 545942 220640 545948 220652
rect 541768 220612 545948 220640
rect 541768 220600 541774 220612
rect 545942 220600 545948 220612
rect 546000 220600 546006 220652
rect 552382 220640 552388 220652
rect 546144 220612 552388 220640
rect 82998 220464 83004 220516
rect 83056 220504 83062 220516
rect 83056 220476 152504 220504
rect 83056 220464 83062 220476
rect 76374 220328 76380 220380
rect 76432 220368 76438 220380
rect 150020 220368 150026 220380
rect 76432 220340 150026 220368
rect 76432 220328 76438 220340
rect 150020 220328 150026 220340
rect 150078 220328 150084 220380
rect 150894 220328 150900 220380
rect 150952 220368 150958 220380
rect 152274 220368 152280 220380
rect 150952 220340 152280 220368
rect 150952 220328 150958 220340
rect 152274 220328 152280 220340
rect 152332 220328 152338 220380
rect 152476 220368 152504 220476
rect 152642 220464 152648 220516
rect 152700 220504 152706 220516
rect 167178 220504 167184 220516
rect 152700 220476 167184 220504
rect 152700 220464 152706 220476
rect 167178 220464 167184 220476
rect 167236 220464 167242 220516
rect 170766 220464 170772 220516
rect 170824 220504 170830 220516
rect 229278 220504 229284 220516
rect 170824 220476 229284 220504
rect 170824 220464 170830 220476
rect 229278 220464 229284 220476
rect 229336 220464 229342 220516
rect 254394 220464 254400 220516
rect 254452 220504 254458 220516
rect 296806 220504 296812 220516
rect 254452 220476 296812 220504
rect 254452 220464 254458 220476
rect 296806 220464 296812 220476
rect 296864 220464 296870 220516
rect 299934 220464 299940 220516
rect 299992 220504 299998 220516
rect 330018 220504 330024 220516
rect 299992 220476 330024 220504
rect 299992 220464 299998 220476
rect 330018 220464 330024 220476
rect 330076 220464 330082 220516
rect 371142 220464 371148 220516
rect 371200 220504 371206 220516
rect 385218 220504 385224 220516
rect 371200 220476 385224 220504
rect 371200 220464 371206 220476
rect 385218 220464 385224 220476
rect 385276 220464 385282 220516
rect 482278 220464 482284 220516
rect 482336 220504 482342 220516
rect 491938 220504 491944 220516
rect 482336 220476 491944 220504
rect 482336 220464 482342 220476
rect 491938 220464 491944 220476
rect 491996 220464 492002 220516
rect 507026 220464 507032 220516
rect 507084 220504 507090 220516
rect 522022 220504 522028 220516
rect 507084 220476 522028 220504
rect 507084 220464 507090 220476
rect 522022 220464 522028 220476
rect 522080 220464 522086 220516
rect 522298 220464 522304 220516
rect 522356 220504 522362 220516
rect 539962 220504 539968 220516
rect 522356 220476 539968 220504
rect 522356 220464 522362 220476
rect 539962 220464 539968 220476
rect 540020 220504 540026 220516
rect 540020 220476 543734 220504
rect 540020 220464 540026 220476
rect 157334 220368 157340 220380
rect 152476 220340 157340 220368
rect 157334 220328 157340 220340
rect 157392 220328 157398 220380
rect 157518 220328 157524 220380
rect 157576 220368 157582 220380
rect 210234 220368 210240 220380
rect 157576 220340 210240 220368
rect 157576 220328 157582 220340
rect 210234 220328 210240 220340
rect 210292 220328 210298 220380
rect 214006 220368 214012 220380
rect 210436 220340 214012 220368
rect 66438 220192 66444 220244
rect 66496 220232 66502 220244
rect 147490 220232 147496 220244
rect 66496 220204 147496 220232
rect 66496 220192 66502 220204
rect 147490 220192 147496 220204
rect 147548 220192 147554 220244
rect 147628 220192 147634 220244
rect 147686 220232 147692 220244
rect 152642 220232 152648 220244
rect 147686 220204 152648 220232
rect 147686 220192 147692 220204
rect 152642 220192 152648 220204
rect 152700 220192 152706 220244
rect 152826 220192 152832 220244
rect 152884 220232 152890 220244
rect 210436 220232 210464 220340
rect 214006 220328 214012 220340
rect 214064 220328 214070 220380
rect 229186 220328 229192 220380
rect 229244 220368 229250 220380
rect 276106 220368 276112 220380
rect 229244 220340 276112 220368
rect 229244 220328 229250 220340
rect 276106 220328 276112 220340
rect 276164 220328 276170 220380
rect 280062 220328 280068 220380
rect 280120 220368 280126 220380
rect 314102 220368 314108 220380
rect 280120 220340 314108 220368
rect 280120 220328 280126 220340
rect 314102 220328 314108 220340
rect 314160 220328 314166 220380
rect 323118 220328 323124 220380
rect 323176 220368 323182 220380
rect 348142 220368 348148 220380
rect 323176 220340 348148 220368
rect 323176 220328 323182 220340
rect 348142 220328 348148 220340
rect 348200 220328 348206 220380
rect 352926 220328 352932 220380
rect 352984 220368 352990 220380
rect 371418 220368 371424 220380
rect 352984 220340 371424 220368
rect 352984 220328 352990 220340
rect 371418 220328 371424 220340
rect 371476 220328 371482 220380
rect 436278 220328 436284 220380
rect 436336 220368 436342 220380
rect 437014 220368 437020 220380
rect 436336 220340 437020 220368
rect 436336 220328 436342 220340
rect 437014 220328 437020 220340
rect 437072 220328 437078 220380
rect 469122 220328 469128 220380
rect 469180 220368 469186 220380
rect 474550 220368 474556 220380
rect 469180 220340 474556 220368
rect 469180 220328 469186 220340
rect 474550 220328 474556 220340
rect 474608 220328 474614 220380
rect 481542 220328 481548 220380
rect 481600 220368 481606 220380
rect 492766 220368 492772 220380
rect 481600 220340 492772 220368
rect 481600 220328 481606 220340
rect 492766 220328 492772 220340
rect 492824 220328 492830 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 510982 220368 510988 220380
rect 496504 220340 510988 220368
rect 496504 220328 496510 220340
rect 510982 220328 510988 220340
rect 511040 220328 511046 220380
rect 517146 220328 517152 220380
rect 517204 220368 517210 220380
rect 539134 220368 539140 220380
rect 517204 220340 539140 220368
rect 517204 220328 517210 220340
rect 539134 220328 539140 220340
rect 539192 220328 539198 220380
rect 543706 220368 543734 220476
rect 543826 220464 543832 220516
rect 543884 220504 543890 220516
rect 546144 220504 546172 220612
rect 552382 220600 552388 220612
rect 552440 220640 552446 220652
rect 557534 220640 557540 220652
rect 552440 220612 557540 220640
rect 552440 220600 552446 220612
rect 557534 220600 557540 220612
rect 557592 220600 557598 220652
rect 558546 220600 558552 220652
rect 558604 220640 558610 220652
rect 559926 220640 559932 220652
rect 558604 220612 559932 220640
rect 558604 220600 558610 220612
rect 559926 220600 559932 220612
rect 559984 220640 559990 220652
rect 626626 220640 626632 220652
rect 559984 220612 626632 220640
rect 559984 220600 559990 220612
rect 626626 220600 626632 220612
rect 626684 220600 626690 220652
rect 543884 220476 546172 220504
rect 543884 220464 543890 220476
rect 546310 220464 546316 220516
rect 546368 220504 546374 220516
rect 553486 220504 553492 220516
rect 546368 220476 553492 220504
rect 546368 220464 546374 220476
rect 553486 220464 553492 220476
rect 553544 220464 553550 220516
rect 554222 220464 554228 220516
rect 554280 220504 554286 220516
rect 625246 220504 625252 220516
rect 554280 220476 625252 220504
rect 554280 220464 554286 220476
rect 625246 220464 625252 220476
rect 625304 220464 625310 220516
rect 622670 220368 622676 220380
rect 543706 220340 622676 220368
rect 622670 220328 622676 220340
rect 622728 220328 622734 220380
rect 211338 220232 211344 220244
rect 152884 220204 210464 220232
rect 210528 220204 211344 220232
rect 152884 220192 152890 220204
rect 63126 220056 63132 220108
rect 63184 220096 63190 220108
rect 140774 220096 140780 220108
rect 63184 220068 140780 220096
rect 63184 220056 63190 220068
rect 140774 220056 140780 220068
rect 140832 220056 140838 220108
rect 140958 220056 140964 220108
rect 141016 220096 141022 220108
rect 147030 220096 147036 220108
rect 141016 220068 147036 220096
rect 141016 220056 141022 220068
rect 147030 220056 147036 220068
rect 147088 220056 147094 220108
rect 150710 220056 150716 220108
rect 150768 220096 150774 220108
rect 210528 220096 210556 220204
rect 211338 220192 211344 220204
rect 211396 220192 211402 220244
rect 217134 220192 217140 220244
rect 217192 220232 217198 220244
rect 265158 220232 265164 220244
rect 217192 220204 265164 220232
rect 217192 220192 217198 220204
rect 265158 220192 265164 220204
rect 265216 220192 265222 220244
rect 280890 220192 280896 220244
rect 280948 220232 280954 220244
rect 317506 220232 317512 220244
rect 280948 220204 317512 220232
rect 280948 220192 280954 220204
rect 317506 220192 317512 220204
rect 317564 220192 317570 220244
rect 332226 220192 332232 220244
rect 332284 220232 332290 220244
rect 357526 220232 357532 220244
rect 332284 220204 357532 220232
rect 332284 220192 332290 220204
rect 357526 220192 357532 220204
rect 357584 220192 357590 220244
rect 360378 220192 360384 220244
rect 360436 220232 360442 220244
rect 377398 220232 377404 220244
rect 360436 220204 377404 220232
rect 360436 220192 360442 220204
rect 377398 220192 377404 220204
rect 377456 220192 377462 220244
rect 390094 220192 390100 220244
rect 390152 220232 390158 220244
rect 401686 220232 401692 220244
rect 390152 220204 401692 220232
rect 390152 220192 390158 220204
rect 401686 220192 401692 220204
rect 401744 220192 401750 220244
rect 430114 220192 430120 220244
rect 430172 220232 430178 220244
rect 432046 220232 432052 220244
rect 430172 220204 432052 220232
rect 430172 220192 430178 220204
rect 432046 220192 432052 220204
rect 432104 220192 432110 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 472986 220192 472992 220244
rect 473044 220232 473050 220244
rect 482002 220232 482008 220244
rect 473044 220204 482008 220232
rect 473044 220192 473050 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 488442 220192 488448 220244
rect 488500 220232 488506 220244
rect 502702 220232 502708 220244
rect 488500 220204 502708 220232
rect 488500 220192 488506 220204
rect 502702 220192 502708 220204
rect 502760 220192 502766 220244
rect 504174 220192 504180 220244
rect 504232 220232 504238 220244
rect 515214 220232 515220 220244
rect 504232 220204 515220 220232
rect 504232 220192 504238 220204
rect 515214 220192 515220 220204
rect 515272 220232 515278 220244
rect 515950 220232 515956 220244
rect 515272 220204 515956 220232
rect 515272 220192 515278 220204
rect 515950 220192 515956 220204
rect 516008 220192 516014 220244
rect 521562 220192 521568 220244
rect 521620 220232 521626 220244
rect 543826 220232 543832 220244
rect 521620 220204 543832 220232
rect 521620 220192 521626 220204
rect 543826 220192 543832 220204
rect 543884 220192 543890 220244
rect 544010 220192 544016 220244
rect 544068 220232 544074 220244
rect 559374 220232 559380 220244
rect 544068 220204 559380 220232
rect 544068 220192 544074 220204
rect 559374 220192 559380 220204
rect 559432 220192 559438 220244
rect 559558 220192 559564 220244
rect 559616 220232 559622 220244
rect 563238 220232 563244 220244
rect 559616 220204 563244 220232
rect 559616 220192 559622 220204
rect 563238 220192 563244 220204
rect 563296 220192 563302 220244
rect 566918 220192 566924 220244
rect 566976 220232 566982 220244
rect 571242 220232 571248 220244
rect 566976 220204 571248 220232
rect 566976 220192 566982 220204
rect 571242 220192 571248 220204
rect 571300 220192 571306 220244
rect 571886 220192 571892 220244
rect 571944 220232 571950 220244
rect 628006 220232 628012 220244
rect 571944 220204 628012 220232
rect 571944 220192 571950 220204
rect 628006 220192 628012 220204
rect 628064 220192 628070 220244
rect 563422 220124 563428 220176
rect 563480 220164 563486 220176
rect 566734 220164 566740 220176
rect 563480 220136 566740 220164
rect 563480 220124 563486 220136
rect 566734 220124 566740 220136
rect 566792 220124 566798 220176
rect 150768 220068 210556 220096
rect 150768 220056 150774 220068
rect 211338 220056 211344 220108
rect 211396 220096 211402 220108
rect 263042 220096 263048 220108
rect 211396 220068 263048 220096
rect 211396 220056 211402 220068
rect 263042 220056 263048 220068
rect 263100 220056 263106 220108
rect 263318 220056 263324 220108
rect 263376 220096 263382 220108
rect 301038 220096 301044 220108
rect 263376 220068 301044 220096
rect 263376 220056 263382 220068
rect 301038 220056 301044 220068
rect 301096 220056 301102 220108
rect 318150 220056 318156 220108
rect 318208 220096 318214 220108
rect 343726 220096 343732 220108
rect 318208 220068 343732 220096
rect 318208 220056 318214 220068
rect 343726 220056 343732 220068
rect 343784 220056 343790 220108
rect 345474 220056 345480 220108
rect 345532 220096 345538 220108
rect 367370 220096 367376 220108
rect 345532 220068 367376 220096
rect 345532 220056 345538 220068
rect 367370 220056 367376 220068
rect 367428 220056 367434 220108
rect 367830 220056 367836 220108
rect 367888 220096 367894 220108
rect 382458 220096 382464 220108
rect 367888 220068 382464 220096
rect 367888 220056 367894 220068
rect 382458 220056 382464 220068
rect 382516 220056 382522 220108
rect 382734 220056 382740 220108
rect 382792 220096 382798 220108
rect 394786 220096 394792 220108
rect 382792 220068 394792 220096
rect 382792 220056 382798 220068
rect 394786 220056 394792 220068
rect 394844 220056 394850 220108
rect 397638 220056 397644 220108
rect 397696 220096 397702 220108
rect 405826 220096 405832 220108
rect 397696 220068 405832 220096
rect 397696 220056 397702 220068
rect 405826 220056 405832 220068
rect 405884 220056 405890 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 431954 220056 431960 220108
rect 432012 220096 432018 220108
rect 434806 220096 434812 220108
rect 432012 220068 434812 220096
rect 432012 220056 432018 220068
rect 434806 220056 434812 220068
rect 434864 220056 434870 220108
rect 478506 220056 478512 220108
rect 478564 220096 478570 220108
rect 489454 220096 489460 220108
rect 478564 220068 489460 220096
rect 478564 220056 478570 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 492306 220056 492312 220108
rect 492364 220096 492370 220108
rect 507670 220096 507676 220108
rect 492364 220068 507676 220096
rect 492364 220056 492370 220068
rect 507670 220056 507676 220068
rect 507728 220056 507734 220108
rect 527818 220056 527824 220108
rect 527876 220096 527882 220108
rect 543688 220096 543694 220108
rect 527876 220068 543694 220096
rect 527876 220056 527882 220068
rect 543688 220056 543694 220068
rect 543746 220056 543752 220108
rect 549990 220056 549996 220108
rect 550048 220096 550054 220108
rect 550450 220096 550456 220108
rect 550048 220068 550456 220096
rect 550048 220056 550054 220068
rect 550450 220056 550456 220068
rect 550508 220056 550514 220108
rect 553486 220056 553492 220108
rect 553544 220096 553550 220108
rect 553544 220068 553900 220096
rect 553544 220056 553550 220068
rect 549438 220028 549444 220040
rect 543936 220000 549444 220028
rect 111242 219920 111248 219972
rect 111300 219960 111306 219972
rect 177206 219960 177212 219972
rect 111300 219932 177212 219960
rect 111300 219920 111306 219932
rect 177206 219920 177212 219932
rect 177264 219920 177270 219972
rect 177390 219920 177396 219972
rect 177448 219960 177454 219972
rect 184382 219960 184388 219972
rect 177448 219932 184388 219960
rect 177448 219920 177454 219932
rect 184382 219920 184388 219932
rect 184440 219920 184446 219972
rect 190638 219920 190644 219972
rect 190696 219960 190702 219972
rect 244458 219960 244464 219972
rect 190696 219932 244464 219960
rect 190696 219920 190702 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 256878 219920 256884 219972
rect 256936 219960 256942 219972
rect 295886 219960 295892 219972
rect 256936 219932 295892 219960
rect 256936 219920 256942 219932
rect 295886 219920 295892 219932
rect 295944 219920 295950 219972
rect 306742 219920 306748 219972
rect 306800 219960 306806 219972
rect 320358 219960 320364 219972
rect 306800 219932 320364 219960
rect 306800 219920 306806 219932
rect 320358 219920 320364 219932
rect 320416 219920 320422 219972
rect 543936 219960 543964 220000
rect 549438 219988 549444 220000
rect 549496 219988 549502 220040
rect 543706 219932 543964 219960
rect 553872 219960 553900 220068
rect 554958 220056 554964 220108
rect 555016 220096 555022 220108
rect 556062 220096 556068 220108
rect 555016 220068 556068 220096
rect 555016 220056 555022 220068
rect 556062 220056 556068 220068
rect 556120 220056 556126 220108
rect 556338 220056 556344 220108
rect 556396 220096 556402 220108
rect 557350 220096 557356 220108
rect 556396 220068 557356 220096
rect 556396 220056 556402 220068
rect 557350 220056 557356 220068
rect 557408 220056 557414 220108
rect 557534 220056 557540 220108
rect 557592 220096 557598 220108
rect 625430 220096 625436 220108
rect 557592 220068 563054 220096
rect 557592 220056 557598 220068
rect 563026 220028 563054 220068
rect 569926 220068 625436 220096
rect 569926 220028 569954 220068
rect 625430 220056 625436 220068
rect 625488 220056 625494 220108
rect 647234 220056 647240 220108
rect 647292 220096 647298 220108
rect 652754 220096 652760 220108
rect 647292 220068 652760 220096
rect 647292 220056 647298 220068
rect 652754 220056 652760 220068
rect 652812 220056 652818 220108
rect 563026 220000 569954 220028
rect 676030 219988 676036 220040
rect 676088 220028 676094 220040
rect 677042 220028 677048 220040
rect 676088 220000 677048 220028
rect 676088 219988 676094 220000
rect 677042 219988 677048 220000
rect 677100 219988 677106 220040
rect 562686 219960 562692 219972
rect 553872 219932 562692 219960
rect 542262 219852 542268 219904
rect 542320 219892 542326 219904
rect 543706 219892 543734 219932
rect 562686 219920 562692 219932
rect 562744 219920 562750 219972
rect 582374 219920 582380 219972
rect 582432 219960 582438 219972
rect 582432 219932 589274 219960
rect 582432 219920 582438 219932
rect 542320 219864 543734 219892
rect 542320 219852 542326 219864
rect 547598 219852 547604 219904
rect 547656 219892 547662 219904
rect 553670 219892 553676 219904
rect 547656 219864 553676 219892
rect 547656 219852 547662 219864
rect 553670 219852 553676 219864
rect 553728 219852 553734 219904
rect 562870 219852 562876 219904
rect 562928 219892 562934 219904
rect 572070 219892 572076 219904
rect 562928 219864 572076 219892
rect 562928 219852 562934 219864
rect 572070 219852 572076 219864
rect 572128 219852 572134 219904
rect 573174 219852 573180 219904
rect 573232 219892 573238 219904
rect 582190 219892 582196 219904
rect 573232 219864 582196 219892
rect 573232 219852 573238 219864
rect 582190 219852 582196 219864
rect 582248 219852 582254 219904
rect 589246 219892 589274 219932
rect 626810 219892 626816 219904
rect 589246 219864 626816 219892
rect 626810 219852 626816 219864
rect 626868 219852 626874 219904
rect 124398 219784 124404 219836
rect 124456 219824 124462 219836
rect 193490 219824 193496 219836
rect 124456 219796 193496 219824
rect 124456 219784 124462 219796
rect 193490 219784 193496 219796
rect 193548 219784 193554 219836
rect 197262 219784 197268 219836
rect 197320 219824 197326 219836
rect 249886 219824 249892 219836
rect 197320 219796 249892 219824
rect 197320 219784 197326 219796
rect 249886 219784 249892 219796
rect 249944 219784 249950 219836
rect 293586 219784 293592 219836
rect 293644 219824 293650 219836
rect 299750 219824 299756 219836
rect 293644 219796 299756 219824
rect 293644 219784 293650 219796
rect 299750 219784 299756 219796
rect 299808 219784 299814 219836
rect 522022 219716 522028 219768
rect 522080 219756 522086 219768
rect 522574 219756 522580 219768
rect 522080 219728 522580 219756
rect 522080 219716 522086 219728
rect 522574 219716 522580 219728
rect 522632 219716 522638 219768
rect 531314 219716 531320 219768
rect 531372 219756 531378 219768
rect 532510 219756 532516 219768
rect 531372 219728 532516 219756
rect 531372 219716 531378 219728
rect 532510 219716 532516 219728
rect 532568 219756 532574 219768
rect 621014 219756 621020 219768
rect 532568 219728 621020 219756
rect 532568 219716 532574 219728
rect 621014 219716 621020 219728
rect 621072 219716 621078 219768
rect 676030 219716 676036 219768
rect 676088 219756 676094 219768
rect 677410 219756 677416 219768
rect 676088 219728 677416 219756
rect 676088 219716 676094 219728
rect 677410 219716 677416 219728
rect 677468 219716 677474 219768
rect 131022 219648 131028 219700
rect 131080 219688 131086 219700
rect 131080 219660 137140 219688
rect 131080 219648 131086 219660
rect 137112 219552 137140 219660
rect 137278 219648 137284 219700
rect 137336 219688 137342 219700
rect 147490 219688 147496 219700
rect 137336 219660 147496 219688
rect 137336 219648 137342 219660
rect 147490 219648 147496 219660
rect 147548 219648 147554 219700
rect 148042 219648 148048 219700
rect 148100 219688 148106 219700
rect 205818 219688 205824 219700
rect 148100 219660 205824 219688
rect 148100 219648 148106 219660
rect 205818 219648 205824 219660
rect 205876 219648 205882 219700
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 668394 219648 668400 219700
rect 668452 219688 668458 219700
rect 669314 219688 669320 219700
rect 668452 219660 669320 219688
rect 668452 219648 668458 219660
rect 669314 219648 669320 219660
rect 669372 219648 669378 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 520182 219580 520188 219632
rect 520240 219620 520246 219632
rect 618254 219620 618260 219632
rect 520240 219592 572392 219620
rect 520240 219580 520246 219592
rect 137462 219552 137468 219564
rect 132512 219524 134012 219552
rect 137112 219524 137468 219552
rect 105814 219444 105820 219496
rect 105872 219484 105878 219496
rect 105872 219456 107148 219484
rect 105872 219444 105878 219456
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 72234 219376 72240 219428
rect 72292 219416 72298 219428
rect 73154 219416 73160 219428
rect 72292 219388 73160 219416
rect 72292 219376 72298 219388
rect 73154 219376 73160 219388
rect 73212 219376 73218 219428
rect 80514 219376 80520 219428
rect 80572 219416 80578 219428
rect 90266 219416 90272 219428
rect 80572 219388 90272 219416
rect 80572 219376 80578 219388
rect 90266 219376 90272 219388
rect 90324 219376 90330 219428
rect 90450 219376 90456 219428
rect 90508 219416 90514 219428
rect 90508 219388 103514 219416
rect 90508 219376 90514 219388
rect 103486 219280 103514 219388
rect 106918 219280 106924 219292
rect 103486 219252 106924 219280
rect 106918 219240 106924 219252
rect 106976 219240 106982 219292
rect 107120 219280 107148 219456
rect 117958 219376 117964 219428
rect 118016 219416 118022 219428
rect 119246 219416 119252 219428
rect 118016 219388 119252 219416
rect 118016 219376 118022 219388
rect 119246 219376 119252 219388
rect 119304 219376 119310 219428
rect 119430 219376 119436 219428
rect 119488 219416 119494 219428
rect 119982 219416 119988 219428
rect 119488 219388 119988 219416
rect 119488 219376 119494 219388
rect 119982 219376 119988 219388
rect 120040 219376 120046 219428
rect 126054 219376 126060 219428
rect 126112 219416 126118 219428
rect 126882 219416 126888 219428
rect 126112 219388 126888 219416
rect 126112 219376 126118 219388
rect 126882 219376 126888 219388
rect 126940 219376 126946 219428
rect 127710 219376 127716 219428
rect 127768 219416 127774 219428
rect 128262 219416 128268 219428
rect 127768 219388 128268 219416
rect 127768 219376 127774 219388
rect 128262 219376 128268 219388
rect 128320 219376 128326 219428
rect 130194 219376 130200 219428
rect 130252 219416 130258 219428
rect 132512 219416 132540 219524
rect 130252 219388 132540 219416
rect 130252 219376 130258 219388
rect 132678 219376 132684 219428
rect 132736 219416 132742 219428
rect 133782 219416 133788 219428
rect 132736 219388 133788 219416
rect 132736 219376 132742 219388
rect 133782 219376 133788 219388
rect 133840 219376 133846 219428
rect 133984 219416 134012 219524
rect 137462 219512 137468 219524
rect 137520 219512 137526 219564
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 203426 219552 203432 219564
rect 137704 219524 203432 219552
rect 137704 219512 137710 219524
rect 203426 219512 203432 219524
rect 203484 219512 203490 219564
rect 210234 219512 210240 219564
rect 210292 219552 210298 219564
rect 218606 219552 218612 219564
rect 210292 219524 218612 219552
rect 210292 219512 210298 219524
rect 218606 219512 218612 219524
rect 218664 219512 218670 219564
rect 270770 219512 270776 219564
rect 270828 219552 270834 219564
rect 279234 219552 279240 219564
rect 270828 219524 279240 219552
rect 270828 219512 270834 219524
rect 279234 219512 279240 219524
rect 279292 219512 279298 219564
rect 515950 219512 515956 219564
rect 516008 219552 516014 219564
rect 572364 219552 572392 219592
rect 572732 219592 618260 219620
rect 572732 219552 572760 219592
rect 618254 219580 618260 219592
rect 618312 219580 618318 219632
rect 516008 219524 520044 219552
rect 572364 219524 572760 219552
rect 516008 219512 516014 219524
rect 221642 219444 221648 219496
rect 221700 219484 221706 219496
rect 221700 219456 222056 219484
rect 221700 219444 221706 219456
rect 142430 219416 142436 219428
rect 133984 219388 142436 219416
rect 142430 219376 142436 219388
rect 142488 219376 142494 219428
rect 142614 219376 142620 219428
rect 142672 219416 142678 219428
rect 143166 219416 143172 219428
rect 142672 219388 143172 219416
rect 142672 219376 142678 219388
rect 143166 219376 143172 219388
rect 143224 219376 143230 219428
rect 143626 219376 143632 219428
rect 143684 219416 143690 219428
rect 197906 219416 197912 219428
rect 143684 219388 197912 219416
rect 143684 219376 143690 219388
rect 197906 219376 197912 219388
rect 197964 219376 197970 219428
rect 199746 219376 199752 219428
rect 199804 219416 199810 219428
rect 204714 219416 204720 219428
rect 199804 219388 204720 219416
rect 199804 219376 199810 219388
rect 204714 219376 204720 219388
rect 204772 219376 204778 219428
rect 208854 219376 208860 219428
rect 208912 219416 208918 219428
rect 209774 219416 209780 219428
rect 208912 219388 209780 219416
rect 208912 219376 208918 219388
rect 209774 219376 209780 219388
rect 209832 219376 209838 219428
rect 222028 219416 222056 219456
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 232498 219416 232504 219428
rect 222028 219388 232504 219416
rect 232498 219376 232504 219388
rect 232556 219376 232562 219428
rect 233694 219376 233700 219428
rect 233752 219416 233758 219428
rect 234614 219416 234620 219428
rect 233752 219388 234620 219416
rect 233752 219376 233758 219388
rect 234614 219376 234620 219388
rect 234672 219376 234678 219428
rect 234816 219388 243584 219416
rect 152366 219280 152372 219292
rect 107120 219252 152372 219280
rect 152366 219240 152372 219252
rect 152424 219240 152430 219292
rect 152550 219240 152556 219292
rect 152608 219280 152614 219292
rect 153102 219280 153108 219292
rect 152608 219252 153108 219280
rect 152608 219240 152614 219252
rect 153102 219240 153108 219252
rect 153160 219240 153166 219292
rect 153378 219240 153384 219292
rect 153436 219280 153442 219292
rect 158990 219280 158996 219292
rect 153436 219252 158996 219280
rect 153436 219240 153442 219252
rect 158990 219240 158996 219252
rect 159048 219240 159054 219292
rect 159174 219240 159180 219292
rect 159232 219280 159238 219292
rect 160002 219280 160008 219292
rect 159232 219252 160008 219280
rect 159232 219240 159238 219252
rect 160002 219240 160008 219252
rect 160060 219240 160066 219292
rect 160186 219240 160192 219292
rect 160244 219280 160250 219292
rect 163958 219280 163964 219292
rect 160244 219252 163964 219280
rect 160244 219240 160250 219252
rect 163958 219240 163964 219252
rect 164016 219240 164022 219292
rect 164970 219240 164976 219292
rect 165028 219280 165034 219292
rect 165430 219280 165436 219292
rect 165028 219252 165436 219280
rect 165028 219240 165034 219252
rect 165430 219240 165436 219252
rect 165488 219240 165494 219292
rect 165798 219240 165804 219292
rect 165856 219280 165862 219292
rect 166534 219280 166540 219292
rect 165856 219252 166540 219280
rect 165856 219240 165862 219252
rect 166534 219240 166540 219252
rect 166592 219240 166598 219292
rect 168926 219280 168932 219292
rect 166736 219252 168932 219280
rect 85298 219104 85304 219156
rect 85356 219144 85362 219156
rect 117958 219144 117964 219156
rect 85356 219116 117964 219144
rect 85356 219104 85362 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 119246 219104 119252 219156
rect 119304 219144 119310 219156
rect 123386 219144 123392 219156
rect 119304 219116 123392 219144
rect 119304 219104 119310 219116
rect 123386 219104 123392 219116
rect 123444 219104 123450 219156
rect 123570 219104 123576 219156
rect 123628 219144 123634 219156
rect 128722 219144 128728 219156
rect 123628 219116 128728 219144
rect 123628 219104 123634 219116
rect 128722 219104 128728 219116
rect 128780 219104 128786 219156
rect 131850 219104 131856 219156
rect 131908 219144 131914 219156
rect 132402 219144 132408 219156
rect 131908 219116 132408 219144
rect 131908 219104 131914 219116
rect 132402 219104 132408 219116
rect 132460 219104 132466 219156
rect 132604 219116 138014 219144
rect 70578 218968 70584 219020
rect 70636 219008 70642 219020
rect 132604 219008 132632 219116
rect 70636 218980 132632 219008
rect 70636 218968 70642 218980
rect 134426 218968 134432 219020
rect 134484 219008 134490 219020
rect 135070 219008 135076 219020
rect 134484 218980 135076 219008
rect 134484 218968 134490 218980
rect 135070 218968 135076 218980
rect 135128 218968 135134 219020
rect 135990 218968 135996 219020
rect 136048 219008 136054 219020
rect 136542 219008 136548 219020
rect 136048 218980 136548 219008
rect 136048 218968 136054 218980
rect 136542 218968 136548 218980
rect 136600 218968 136606 219020
rect 136818 218968 136824 219020
rect 136876 219008 136882 219020
rect 137830 219008 137836 219020
rect 136876 218980 137836 219008
rect 136876 218968 136882 218980
rect 137830 218968 137836 218980
rect 137888 218968 137894 219020
rect 137986 219008 138014 219116
rect 138106 219104 138112 219156
rect 138164 219144 138170 219156
rect 143626 219144 143632 219156
rect 138164 219116 143632 219144
rect 138164 219104 138170 219116
rect 143626 219104 143632 219116
rect 143684 219104 143690 219156
rect 143810 219104 143816 219156
rect 143868 219144 143874 219156
rect 152274 219144 152280 219156
rect 143868 219116 152280 219144
rect 143868 219104 143874 219116
rect 152274 219104 152280 219116
rect 152332 219104 152338 219156
rect 166736 219144 166764 219252
rect 168926 219240 168932 219252
rect 168984 219240 168990 219292
rect 169294 219240 169300 219292
rect 169352 219280 169358 219292
rect 169352 219252 190454 219280
rect 169352 219240 169358 219252
rect 152476 219116 166764 219144
rect 139946 219008 139952 219020
rect 137986 218980 139952 219008
rect 139946 218968 139952 218980
rect 140004 218968 140010 219020
rect 140130 218968 140136 219020
rect 140188 219008 140194 219020
rect 142246 219008 142252 219020
rect 140188 218980 142252 219008
rect 140188 218968 140194 218980
rect 142246 218968 142252 218980
rect 142304 218968 142310 219020
rect 142430 218968 142436 219020
rect 142488 219008 142494 219020
rect 152476 219008 152504 219116
rect 166994 219104 167000 219156
rect 167052 219144 167058 219156
rect 190086 219144 190092 219156
rect 167052 219116 190092 219144
rect 167052 219104 167058 219116
rect 190086 219104 190092 219116
rect 190144 219104 190150 219156
rect 190426 219144 190454 219252
rect 193122 219240 193128 219292
rect 193180 219280 193186 219292
rect 195422 219280 195428 219292
rect 193180 219252 195428 219280
rect 193180 219240 193186 219252
rect 195422 219240 195428 219252
rect 195480 219240 195486 219292
rect 196066 219240 196072 219292
rect 196124 219280 196130 219292
rect 199378 219280 199384 219292
rect 196124 219252 199384 219280
rect 196124 219240 196130 219252
rect 199378 219240 199384 219252
rect 199436 219240 199442 219292
rect 226886 219280 226892 219292
rect 200086 219252 226892 219280
rect 195054 219144 195060 219156
rect 190426 219116 195060 219144
rect 195054 219104 195060 219116
rect 195112 219104 195118 219156
rect 195238 219104 195244 219156
rect 195296 219144 195302 219156
rect 200086 219144 200114 219252
rect 226886 219240 226892 219252
rect 226944 219240 226950 219292
rect 232866 219240 232872 219292
rect 232924 219280 232930 219292
rect 234816 219280 234844 219388
rect 232924 219252 234844 219280
rect 232924 219240 232930 219252
rect 237834 219240 237840 219292
rect 237892 219280 237898 219292
rect 239398 219280 239404 219292
rect 237892 219252 239404 219280
rect 237892 219240 237898 219252
rect 239398 219240 239404 219252
rect 239456 219240 239462 219292
rect 243556 219280 243584 219388
rect 246114 219376 246120 219428
rect 246172 219416 246178 219428
rect 285950 219416 285956 219428
rect 246172 219388 285956 219416
rect 246172 219376 246178 219388
rect 285950 219376 285956 219388
rect 286008 219376 286014 219428
rect 287514 219376 287520 219428
rect 287572 219416 287578 219428
rect 288434 219416 288440 219428
rect 287572 219388 288440 219416
rect 287572 219376 287578 219388
rect 288434 219376 288440 219388
rect 288492 219376 288498 219428
rect 291654 219376 291660 219428
rect 291712 219416 291718 219428
rect 324682 219416 324688 219428
rect 291712 219388 324688 219416
rect 291712 219376 291718 219388
rect 324682 219376 324688 219388
rect 324740 219376 324746 219428
rect 325602 219376 325608 219428
rect 325660 219416 325666 219428
rect 326338 219416 326344 219428
rect 325660 219388 326344 219416
rect 325660 219376 325666 219388
rect 326338 219376 326344 219388
rect 326396 219376 326402 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 366358 219416 366364 219428
rect 352156 219388 366364 219416
rect 352156 219376 352162 219388
rect 366358 219376 366364 219388
rect 366416 219376 366422 219428
rect 374454 219376 374460 219428
rect 374512 219416 374518 219428
rect 375374 219416 375380 219428
rect 374512 219388 375380 219416
rect 374512 219376 374518 219388
rect 375374 219376 375380 219388
rect 375432 219376 375438 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384298 219416 384304 219428
rect 380308 219388 384304 219416
rect 380308 219376 380314 219388
rect 384298 219376 384304 219388
rect 384356 219376 384362 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 403434 219376 403440 219428
rect 403492 219416 403498 219428
rect 404354 219416 404360 219428
rect 403492 219388 404360 219416
rect 403492 219376 403498 219388
rect 404354 219376 404360 219388
rect 404412 219376 404418 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 520016 219484 520044 219524
rect 557718 219484 557724 219496
rect 520016 219456 557724 219484
rect 557718 219444 557724 219456
rect 557776 219444 557782 219496
rect 558730 219444 558736 219496
rect 558788 219484 558794 219496
rect 558788 219456 572300 219484
rect 558788 219444 558794 219456
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 438210 219376 438216 219428
rect 438268 219416 438274 219428
rect 438854 219416 438860 219428
rect 438268 219388 438860 219416
rect 438268 219376 438274 219388
rect 438854 219376 438860 219388
rect 438912 219376 438918 219428
rect 439866 219376 439872 219428
rect 439924 219416 439930 219428
rect 440326 219416 440332 219428
rect 439924 219388 440332 219416
rect 439924 219376 439930 219388
rect 440326 219376 440332 219388
rect 440384 219376 440390 219428
rect 488718 219376 488724 219428
rect 488776 219416 488782 219428
rect 489178 219416 489184 219428
rect 488776 219388 489184 219416
rect 488776 219376 488782 219388
rect 489178 219376 489184 219388
rect 489236 219376 489242 219428
rect 518802 219376 518808 219428
rect 518860 219416 518866 219428
rect 519814 219416 519820 219428
rect 518860 219388 519820 219416
rect 518860 219376 518866 219388
rect 519814 219376 519820 219388
rect 519872 219376 519878 219428
rect 572272 219416 572300 219456
rect 572824 219456 601694 219484
rect 572824 219416 572852 219456
rect 558012 219388 558316 219416
rect 572272 219388 572852 219416
rect 504634 219308 504640 219360
rect 504692 219348 504698 219360
rect 505278 219348 505284 219360
rect 504692 219320 505284 219348
rect 504692 219308 504698 219320
rect 505278 219308 505284 219320
rect 505336 219308 505342 219360
rect 540238 219308 540244 219360
rect 540296 219348 540302 219360
rect 540790 219348 540796 219360
rect 540296 219320 540796 219348
rect 540296 219308 540302 219320
rect 540790 219308 540796 219320
rect 540848 219348 540854 219360
rect 542262 219348 542268 219360
rect 540848 219320 542268 219348
rect 540848 219308 540854 219320
rect 542262 219308 542268 219320
rect 542320 219308 542326 219360
rect 542446 219308 542452 219360
rect 542504 219348 542510 219360
rect 555602 219348 555608 219360
rect 542504 219320 555608 219348
rect 542504 219308 542510 219320
rect 555602 219308 555608 219320
rect 555660 219308 555666 219360
rect 555786 219308 555792 219360
rect 555844 219348 555850 219360
rect 558012 219348 558040 219388
rect 555844 219320 558040 219348
rect 558288 219348 558316 219388
rect 571978 219348 571984 219360
rect 558288 219320 571984 219348
rect 555844 219308 555850 219320
rect 571978 219308 571984 219320
rect 572036 219308 572042 219360
rect 573818 219308 573824 219360
rect 573876 219348 573882 219360
rect 575290 219348 575296 219360
rect 573876 219320 575296 219348
rect 573876 219308 573882 219320
rect 575290 219308 575296 219320
rect 575348 219308 575354 219360
rect 582190 219308 582196 219360
rect 582248 219348 582254 219360
rect 599026 219348 599032 219360
rect 582248 219320 599032 219348
rect 582248 219308 582254 219320
rect 599026 219308 599032 219320
rect 599084 219308 599090 219360
rect 601666 219348 601694 219456
rect 601786 219444 601792 219496
rect 601844 219484 601850 219496
rect 628190 219484 628196 219496
rect 601844 219456 628196 219484
rect 601844 219444 601850 219456
rect 628190 219444 628196 219456
rect 628248 219444 628254 219496
rect 676214 219376 676220 219428
rect 676272 219416 676278 219428
rect 677594 219416 677600 219428
rect 676272 219388 677600 219416
rect 676272 219376 676278 219388
rect 677594 219376 677600 219388
rect 677652 219376 677658 219428
rect 601970 219348 601976 219360
rect 601666 219320 601976 219348
rect 601970 219308 601976 219320
rect 602028 219308 602034 219360
rect 270770 219280 270776 219292
rect 243556 219252 270776 219280
rect 270770 219240 270776 219252
rect 270828 219240 270834 219292
rect 327258 219240 327264 219292
rect 327316 219280 327322 219292
rect 327316 219252 345014 219280
rect 327316 219240 327322 219252
rect 195296 219116 200114 219144
rect 200408 219116 201724 219144
rect 195296 219104 195302 219116
rect 142488 218980 152504 219008
rect 142488 218968 142494 218980
rect 152734 218968 152740 219020
rect 152792 219008 152798 219020
rect 166258 219008 166264 219020
rect 152792 218980 166264 219008
rect 152792 218968 152798 218980
rect 166258 218968 166264 218980
rect 166316 218968 166322 219020
rect 167178 218968 167184 219020
rect 167236 219008 167242 219020
rect 200408 219008 200436 219116
rect 167236 218980 200436 219008
rect 167236 218968 167242 218980
rect 200574 218968 200580 219020
rect 200632 219008 200638 219020
rect 201494 219008 201500 219020
rect 200632 218980 201500 219008
rect 200632 218968 200638 218980
rect 201494 218968 201500 218980
rect 201552 218968 201558 219020
rect 201696 219008 201724 219116
rect 204714 219104 204720 219156
rect 204772 219144 204778 219156
rect 246298 219144 246304 219156
rect 204772 219116 246304 219144
rect 204772 219104 204778 219116
rect 246298 219104 246304 219116
rect 246356 219104 246362 219156
rect 258534 219104 258540 219156
rect 258592 219144 258598 219156
rect 259270 219144 259276 219156
rect 258592 219116 259276 219144
rect 258592 219104 258598 219116
rect 259270 219104 259276 219116
rect 259328 219104 259334 219156
rect 259454 219104 259460 219156
rect 259512 219144 259518 219156
rect 291838 219144 291844 219156
rect 259512 219116 291844 219144
rect 259512 219104 259518 219116
rect 291838 219104 291844 219116
rect 291896 219104 291902 219156
rect 294138 219104 294144 219156
rect 294196 219144 294202 219156
rect 311802 219144 311808 219156
rect 294196 219116 311808 219144
rect 294196 219104 294202 219116
rect 311802 219104 311808 219116
rect 311860 219104 311866 219156
rect 315666 219104 315672 219156
rect 315724 219144 315730 219156
rect 317966 219144 317972 219156
rect 315724 219116 317972 219144
rect 315724 219104 315730 219116
rect 317966 219104 317972 219116
rect 318024 219104 318030 219156
rect 320634 219104 320640 219156
rect 320692 219144 320698 219156
rect 340138 219144 340144 219156
rect 320692 219116 340144 219144
rect 320692 219104 320698 219116
rect 340138 219104 340144 219116
rect 340196 219104 340202 219156
rect 344986 219144 345014 219252
rect 383562 219240 383568 219292
rect 383620 219280 383626 219292
rect 387058 219280 387064 219292
rect 383620 219252 387064 219280
rect 383620 219240 383626 219252
rect 387058 219240 387064 219252
rect 387116 219240 387122 219292
rect 450722 219240 450728 219292
rect 450780 219280 450786 219292
rect 453850 219280 453856 219292
rect 450780 219252 453856 219280
rect 450780 219240 450786 219252
rect 453850 219240 453856 219252
rect 453908 219240 453914 219292
rect 479702 219240 479708 219292
rect 479760 219280 479766 219292
rect 480346 219280 480352 219292
rect 479760 219252 480352 219280
rect 479760 219240 479766 219252
rect 480346 219240 480352 219252
rect 480404 219240 480410 219292
rect 534166 219240 534172 219292
rect 534224 219280 534230 219292
rect 534626 219280 534632 219292
rect 534224 219252 534632 219280
rect 534224 219240 534230 219252
rect 534626 219240 534632 219252
rect 534684 219240 534690 219292
rect 544930 219172 544936 219224
rect 544988 219212 544994 219224
rect 553486 219212 553492 219224
rect 544988 219184 553492 219212
rect 544988 219172 544994 219184
rect 553486 219172 553492 219184
rect 553544 219172 553550 219224
rect 566550 219212 566556 219224
rect 558886 219184 566556 219212
rect 345658 219144 345664 219156
rect 344986 219116 345664 219144
rect 345658 219104 345664 219116
rect 345716 219104 345722 219156
rect 352558 219144 352564 219156
rect 348758 219116 352564 219144
rect 204898 219008 204904 219020
rect 201696 218980 204904 219008
rect 204898 218968 204904 218980
rect 204956 218968 204962 219020
rect 206370 218968 206376 219020
rect 206428 219008 206434 219020
rect 255866 219008 255872 219020
rect 206428 218980 255872 219008
rect 206428 218968 206434 218980
rect 255866 218968 255872 218980
rect 255924 218968 255930 219020
rect 259270 218968 259276 219020
rect 259328 219008 259334 219020
rect 293586 219008 293592 219020
rect 259328 218980 293592 219008
rect 259328 218968 259334 218980
rect 293586 218968 293592 218980
rect 293644 218968 293650 219020
rect 300762 218968 300768 219020
rect 300820 219008 300826 219020
rect 329282 219008 329288 219020
rect 300820 218980 329288 219008
rect 300820 218968 300826 218980
rect 329282 218968 329288 218980
rect 329340 218968 329346 219020
rect 333698 218968 333704 219020
rect 333756 219008 333762 219020
rect 348758 219008 348786 219116
rect 352558 219104 352564 219116
rect 352616 219104 352622 219156
rect 354398 219104 354404 219156
rect 354456 219144 354462 219156
rect 355502 219144 355508 219156
rect 354456 219116 355508 219144
rect 354456 219104 354462 219116
rect 355502 219104 355508 219116
rect 355560 219104 355566 219156
rect 358722 219104 358728 219156
rect 358780 219144 358786 219156
rect 364978 219144 364984 219156
rect 358780 219116 364984 219144
rect 358780 219104 358786 219116
rect 364978 219104 364984 219116
rect 365036 219104 365042 219156
rect 419166 219104 419172 219156
rect 419224 219144 419230 219156
rect 422662 219144 422668 219156
rect 419224 219116 422668 219144
rect 419224 219104 419230 219116
rect 422662 219104 422668 219116
rect 422720 219104 422726 219156
rect 483566 219104 483572 219156
rect 483624 219144 483630 219156
rect 490282 219144 490288 219156
rect 483624 219116 490288 219144
rect 483624 219104 483630 219116
rect 490282 219104 490288 219116
rect 490340 219104 490346 219156
rect 503070 219104 503076 219156
rect 503128 219144 503134 219156
rect 503530 219144 503536 219156
rect 503128 219116 503536 219144
rect 503128 219104 503134 219116
rect 503530 219104 503536 219116
rect 503588 219104 503594 219156
rect 507118 219104 507124 219156
rect 507176 219144 507182 219156
rect 514938 219144 514944 219156
rect 507176 219116 514944 219144
rect 507176 219104 507182 219116
rect 514938 219104 514944 219116
rect 514996 219104 515002 219156
rect 535178 219104 535184 219156
rect 535236 219144 535242 219156
rect 544010 219144 544016 219156
rect 535236 219116 544016 219144
rect 535236 219104 535242 219116
rect 544010 219104 544016 219116
rect 544068 219104 544074 219156
rect 558270 219144 558276 219156
rect 553688 219116 558276 219144
rect 544470 219036 544476 219088
rect 544528 219076 544534 219088
rect 544528 219048 549254 219076
rect 544528 219036 544534 219048
rect 333756 218980 348786 219008
rect 333756 218968 333762 218980
rect 351362 218968 351368 219020
rect 351420 219008 351426 219020
rect 355226 219008 355232 219020
rect 351420 218980 355232 219008
rect 351420 218968 351426 218980
rect 355226 218968 355232 218980
rect 355284 218968 355290 219020
rect 355410 218968 355416 219020
rect 355468 219008 355474 219020
rect 369118 219008 369124 219020
rect 355468 218980 369124 219008
rect 355468 218968 355474 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 373626 218968 373632 219020
rect 373684 219008 373690 219020
rect 380066 219008 380072 219020
rect 373684 218980 380072 219008
rect 373684 218968 373690 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 384390 218968 384396 219020
rect 384448 219008 384454 219020
rect 393958 219008 393964 219020
rect 384448 218980 393964 219008
rect 384448 218968 384454 218980
rect 393958 218968 393964 218980
rect 394016 218968 394022 219020
rect 401778 218968 401784 219020
rect 401836 219008 401842 219020
rect 407758 219008 407764 219020
rect 401836 218980 407764 219008
rect 401836 218968 401842 218980
rect 407758 218968 407764 218980
rect 407816 218968 407822 219020
rect 514754 218968 514760 219020
rect 514812 219008 514818 219020
rect 519814 219008 519820 219020
rect 514812 218980 519820 219008
rect 514812 218968 514818 218980
rect 519814 218968 519820 218980
rect 519872 218968 519878 219020
rect 524414 218968 524420 219020
rect 524472 219008 524478 219020
rect 544194 219008 544200 219020
rect 524472 218980 544200 219008
rect 524472 218968 524478 218980
rect 544194 218968 544200 218980
rect 544252 218968 544258 219020
rect 549226 219008 549254 219048
rect 553688 219008 553716 219116
rect 558270 219104 558276 219116
rect 558328 219104 558334 219156
rect 558730 219104 558736 219156
rect 558788 219144 558794 219156
rect 558886 219144 558914 219184
rect 566550 219172 566556 219184
rect 566608 219172 566614 219224
rect 567838 219172 567844 219224
rect 567896 219212 567902 219224
rect 573266 219212 573272 219224
rect 567896 219184 573272 219212
rect 567896 219172 567902 219184
rect 573266 219172 573272 219184
rect 573324 219172 573330 219224
rect 573450 219172 573456 219224
rect 573508 219212 573514 219224
rect 582282 219212 582288 219224
rect 573508 219184 582288 219212
rect 573508 219172 573514 219184
rect 582282 219172 582288 219184
rect 582340 219172 582346 219224
rect 558788 219116 558914 219144
rect 558788 219104 558794 219116
rect 567010 219104 567016 219156
rect 567068 219144 567074 219156
rect 567068 219116 567700 219144
rect 567068 219104 567074 219116
rect 549226 218980 553716 219008
rect 553854 218968 553860 219020
rect 553912 219008 553918 219020
rect 555234 219008 555240 219020
rect 553912 218980 555240 219008
rect 553912 218968 553918 218980
rect 555234 218968 555240 218980
rect 555292 218968 555298 219020
rect 555602 218968 555608 219020
rect 555660 219008 555666 219020
rect 567194 219008 567200 219020
rect 555660 218980 557856 219008
rect 555660 218968 555666 218980
rect 62298 218832 62304 218884
rect 62356 218872 62362 218884
rect 76558 218872 76564 218884
rect 62356 218844 76564 218872
rect 62356 218832 62362 218844
rect 76558 218832 76564 218844
rect 76616 218832 76622 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 152090 218872 152096 218884
rect 83884 218844 152096 218872
rect 83884 218832 83890 218844
rect 152090 218832 152096 218844
rect 152148 218832 152154 218884
rect 152274 218832 152280 218884
rect 152332 218872 152338 218884
rect 166442 218872 166448 218884
rect 152332 218844 166448 218872
rect 152332 218832 152338 218844
rect 166442 218832 166448 218844
rect 166500 218832 166506 218884
rect 167178 218832 167184 218884
rect 167236 218872 167242 218884
rect 215938 218872 215944 218884
rect 167236 218844 215944 218872
rect 167236 218832 167242 218844
rect 215938 218832 215944 218844
rect 215996 218832 216002 218884
rect 217962 218832 217968 218884
rect 218020 218872 218026 218884
rect 220078 218872 220084 218884
rect 218020 218844 220084 218872
rect 218020 218832 218026 218844
rect 220078 218832 220084 218844
rect 220136 218832 220142 218884
rect 220280 218844 224448 218872
rect 77202 218696 77208 218748
rect 77260 218736 77266 218748
rect 147490 218736 147496 218748
rect 77260 218708 147496 218736
rect 77260 218696 77266 218708
rect 147490 218696 147496 218708
rect 147548 218696 147554 218748
rect 152734 218736 152740 218748
rect 147646 218708 152740 218736
rect 59814 218560 59820 218612
rect 59872 218600 59878 218612
rect 69566 218600 69572 218612
rect 59872 218572 69572 218600
rect 59872 218560 59878 218572
rect 69566 218560 69572 218572
rect 69624 218560 69630 218612
rect 92934 218560 92940 218612
rect 92992 218600 92998 218612
rect 93762 218600 93768 218612
rect 92992 218572 93768 218600
rect 92992 218560 92998 218572
rect 93762 218560 93768 218572
rect 93820 218560 93826 218612
rect 139946 218600 139952 218612
rect 103486 218572 139952 218600
rect 93762 218424 93768 218476
rect 93820 218464 93826 218476
rect 103486 218464 103514 218572
rect 139946 218560 139952 218572
rect 140004 218560 140010 218612
rect 140130 218560 140136 218612
rect 140188 218600 140194 218612
rect 143810 218600 143816 218612
rect 140188 218572 143816 218600
rect 140188 218560 140194 218572
rect 143810 218560 143816 218572
rect 143868 218560 143874 218612
rect 144270 218560 144276 218612
rect 144328 218600 144334 218612
rect 144822 218600 144828 218612
rect 144328 218572 144828 218600
rect 144328 218560 144334 218572
rect 144822 218560 144828 218572
rect 144880 218560 144886 218612
rect 146754 218560 146760 218612
rect 146812 218600 146818 218612
rect 147646 218600 147674 218708
rect 152734 218696 152740 218708
rect 152792 218696 152798 218748
rect 152918 218696 152924 218748
rect 152976 218736 152982 218748
rect 156322 218736 156328 218748
rect 152976 218708 156328 218736
rect 152976 218696 152982 218708
rect 156322 218696 156328 218708
rect 156380 218696 156386 218748
rect 156690 218696 156696 218748
rect 156748 218736 156754 218748
rect 162118 218736 162124 218748
rect 156748 218708 162124 218736
rect 156748 218696 156754 218708
rect 162118 218696 162124 218708
rect 162176 218696 162182 218748
rect 166258 218736 166264 218748
rect 162320 218708 166264 218736
rect 146812 218572 147674 218600
rect 146812 218560 146818 218572
rect 149054 218560 149060 218612
rect 149112 218600 149118 218612
rect 157978 218600 157984 218612
rect 149112 218572 157984 218600
rect 149112 218560 149118 218572
rect 157978 218560 157984 218572
rect 158036 218560 158042 218612
rect 158990 218560 158996 218612
rect 159048 218600 159054 218612
rect 162320 218600 162348 218708
rect 166258 218696 166264 218708
rect 166316 218696 166322 218748
rect 167362 218696 167368 218748
rect 167420 218736 167426 218748
rect 213178 218736 213184 218748
rect 167420 218708 213184 218736
rect 167420 218696 167426 218708
rect 213178 218696 213184 218708
rect 213236 218696 213242 218748
rect 213546 218696 213552 218748
rect 213604 218736 213610 218748
rect 217318 218736 217324 218748
rect 213604 218708 217324 218736
rect 213604 218696 213610 218708
rect 217318 218696 217324 218708
rect 217376 218696 217382 218748
rect 218790 218696 218796 218748
rect 218848 218736 218854 218748
rect 219342 218736 219348 218748
rect 218848 218708 219348 218736
rect 218848 218696 218854 218708
rect 219342 218696 219348 218708
rect 219400 218696 219406 218748
rect 219618 218696 219624 218748
rect 219676 218736 219682 218748
rect 220280 218736 220308 218844
rect 219676 218708 220308 218736
rect 219676 218696 219682 218708
rect 221090 218696 221096 218748
rect 221148 218736 221154 218748
rect 224218 218736 224224 218748
rect 221148 218708 224224 218736
rect 221148 218696 221154 218708
rect 224218 218696 224224 218708
rect 224276 218696 224282 218748
rect 224420 218736 224448 218844
rect 225966 218832 225972 218884
rect 226024 218872 226030 218884
rect 226024 218844 264330 218872
rect 226024 218832 226030 218844
rect 264146 218736 264152 218748
rect 224420 218708 264152 218736
rect 264146 218696 264152 218708
rect 264204 218696 264210 218748
rect 159048 218572 162348 218600
rect 159048 218560 159054 218572
rect 162670 218560 162676 218612
rect 162728 218600 162734 218612
rect 166534 218600 166540 218612
rect 162728 218572 166540 218600
rect 162728 218560 162734 218572
rect 166534 218560 166540 218572
rect 166592 218560 166598 218612
rect 169938 218560 169944 218612
rect 169996 218600 170002 218612
rect 181070 218600 181076 218612
rect 169996 218572 181076 218600
rect 169996 218560 170002 218572
rect 181070 218560 181076 218572
rect 181128 218560 181134 218612
rect 182358 218560 182364 218612
rect 182416 218600 182422 218612
rect 183278 218600 183284 218612
rect 182416 218572 183284 218600
rect 182416 218560 182422 218572
rect 183278 218560 183284 218572
rect 183336 218560 183342 218612
rect 195238 218600 195244 218612
rect 186286 218572 195244 218600
rect 93820 218436 103514 218464
rect 93820 218424 93826 218436
rect 113634 218424 113640 218476
rect 113692 218464 113698 218476
rect 119982 218464 119988 218476
rect 113692 218436 119988 218464
rect 113692 218424 113698 218436
rect 119982 218424 119988 218436
rect 120040 218424 120046 218476
rect 128722 218424 128728 218476
rect 128780 218464 128786 218476
rect 174538 218464 174544 218476
rect 128780 218436 174544 218464
rect 128780 218424 128786 218436
rect 174538 218424 174544 218436
rect 174596 218424 174602 218476
rect 174722 218424 174728 218476
rect 174780 218464 174786 218476
rect 186286 218464 186314 218572
rect 195238 218560 195244 218572
rect 195296 218560 195302 218612
rect 195422 218560 195428 218612
rect 195480 218600 195486 218612
rect 243446 218600 243452 218612
rect 195480 218572 243452 218600
rect 195480 218560 195486 218572
rect 243446 218560 243452 218572
rect 243504 218560 243510 218612
rect 252738 218560 252744 218612
rect 252796 218600 252802 218612
rect 259454 218600 259460 218612
rect 252796 218572 259460 218600
rect 252796 218560 252802 218572
rect 259454 218560 259460 218572
rect 259512 218560 259518 218612
rect 264302 218600 264330 218844
rect 274266 218832 274272 218884
rect 274324 218872 274330 218884
rect 280706 218872 280712 218884
rect 274324 218844 280712 218872
rect 274324 218832 274330 218844
rect 280706 218832 280712 218844
rect 280764 218832 280770 218884
rect 281074 218832 281080 218884
rect 281132 218872 281138 218884
rect 312538 218872 312544 218884
rect 281132 218844 312544 218872
rect 281132 218832 281138 218844
rect 312538 218832 312544 218844
rect 312596 218832 312602 218884
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 329098 218872 329104 218884
rect 314068 218844 329104 218872
rect 314068 218832 314074 218844
rect 329098 218832 329104 218844
rect 329156 218832 329162 218884
rect 337194 218832 337200 218884
rect 337252 218872 337258 218884
rect 357710 218872 357716 218884
rect 337252 218844 357716 218872
rect 337252 218832 337258 218844
rect 357710 218832 357716 218844
rect 357768 218832 357774 218884
rect 366726 218832 366732 218884
rect 366784 218872 366790 218884
rect 378778 218872 378784 218884
rect 366784 218844 378784 218872
rect 366784 218832 366790 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 386046 218832 386052 218884
rect 386104 218872 386110 218884
rect 396626 218872 396632 218884
rect 386104 218844 396632 218872
rect 386104 218832 386110 218844
rect 396626 218832 396632 218844
rect 396684 218832 396690 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412450 218872 412456 218884
rect 411772 218844 412456 218872
rect 411772 218832 411778 218844
rect 412450 218832 412456 218844
rect 412508 218832 412514 218884
rect 505830 218832 505836 218884
rect 505888 218872 505894 218884
rect 505888 218844 519124 218872
rect 505888 218832 505894 218844
rect 265986 218696 265992 218748
rect 266044 218736 266050 218748
rect 302878 218736 302884 218748
rect 266044 218708 302884 218736
rect 266044 218696 266050 218708
rect 302878 218696 302884 218708
rect 302936 218696 302942 218748
rect 307386 218696 307392 218748
rect 307444 218736 307450 218748
rect 337010 218736 337016 218748
rect 307444 218708 337016 218736
rect 307444 218696 307450 218708
rect 337010 218696 337016 218708
rect 337068 218696 337074 218748
rect 340506 218696 340512 218748
rect 340564 218736 340570 218748
rect 360838 218736 360844 218748
rect 340564 218708 360844 218736
rect 340564 218696 340570 218708
rect 360838 218696 360844 218708
rect 360896 218696 360902 218748
rect 379146 218696 379152 218748
rect 379204 218736 379210 218748
rect 392118 218736 392124 218748
rect 379204 218708 392124 218736
rect 379204 218696 379210 218708
rect 392118 218696 392124 218708
rect 392176 218696 392182 218748
rect 395798 218696 395804 218748
rect 395856 218736 395862 218748
rect 404538 218736 404544 218748
rect 395856 218708 404544 218736
rect 395856 218696 395862 218708
rect 404538 218696 404544 218708
rect 404596 218696 404602 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 460198 218696 460204 218748
rect 460256 218736 460262 218748
rect 461302 218736 461308 218748
rect 460256 218708 461308 218736
rect 460256 218696 460262 218708
rect 461302 218696 461308 218708
rect 461360 218696 461366 218748
rect 518802 218736 518808 218748
rect 514726 218708 518808 218736
rect 502518 218628 502524 218680
rect 502576 218668 502582 218680
rect 505002 218668 505008 218680
rect 502576 218640 505008 218668
rect 502576 218628 502582 218640
rect 505002 218628 505008 218640
rect 505060 218628 505066 218680
rect 267826 218600 267832 218612
rect 264302 218572 267832 218600
rect 267826 218560 267832 218572
rect 267884 218560 267890 218612
rect 272610 218560 272616 218612
rect 272668 218600 272674 218612
rect 296990 218600 296996 218612
rect 272668 218572 296996 218600
rect 272668 218560 272674 218572
rect 296990 218560 296996 218572
rect 297048 218560 297054 218612
rect 429930 218560 429936 218612
rect 429988 218600 429994 218612
rect 432690 218600 432696 218612
rect 429988 218572 432696 218600
rect 429988 218560 429994 218572
rect 432690 218560 432696 218572
rect 432748 218560 432754 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 514726 218600 514754 218708
rect 518802 218696 518808 218708
rect 518860 218696 518866 218748
rect 519096 218736 519124 218844
rect 519538 218832 519544 218884
rect 519596 218872 519602 218884
rect 526438 218872 526444 218884
rect 519596 218844 526444 218872
rect 519596 218832 519602 218844
rect 526438 218832 526444 218844
rect 526496 218832 526502 218884
rect 533430 218832 533436 218884
rect 533488 218872 533494 218884
rect 533890 218872 533896 218884
rect 533488 218844 533896 218872
rect 533488 218832 533494 218844
rect 533890 218832 533896 218844
rect 533948 218832 533954 218884
rect 537570 218832 537576 218884
rect 537628 218872 537634 218884
rect 537628 218844 548472 218872
rect 537628 218832 537634 218844
rect 524598 218736 524604 218748
rect 519096 218708 524604 218736
rect 524598 218696 524604 218708
rect 524656 218696 524662 218748
rect 525058 218696 525064 218748
rect 525116 218736 525122 218748
rect 529382 218736 529388 218748
rect 525116 218708 529388 218736
rect 525116 218696 525122 218708
rect 529382 218696 529388 218708
rect 529440 218696 529446 218748
rect 533614 218696 533620 218748
rect 533672 218736 533678 218748
rect 534350 218736 534356 218748
rect 533672 218708 534356 218736
rect 533672 218696 533678 218708
rect 534350 218696 534356 218708
rect 534408 218696 534414 218748
rect 534994 218696 535000 218748
rect 535052 218736 535058 218748
rect 547966 218736 547972 218748
rect 535052 218708 547972 218736
rect 535052 218696 535058 218708
rect 547966 218696 547972 218708
rect 548024 218696 548030 218748
rect 548444 218736 548472 218844
rect 549070 218832 549076 218884
rect 549128 218872 549134 218884
rect 556154 218872 556160 218884
rect 549128 218844 556160 218872
rect 549128 218832 549134 218844
rect 556154 218832 556160 218844
rect 556212 218832 556218 218884
rect 557828 218872 557856 218980
rect 558380 218980 567200 219008
rect 558380 218940 558408 218980
rect 567194 218968 567200 218980
rect 567252 218968 567258 219020
rect 567672 219008 567700 219116
rect 572254 219036 572260 219088
rect 572312 219076 572318 219088
rect 574554 219076 574560 219088
rect 572312 219048 574560 219076
rect 572312 219036 572318 219048
rect 574554 219036 574560 219048
rect 574612 219036 574618 219088
rect 571794 219008 571800 219020
rect 567672 218980 571800 219008
rect 571794 218968 571800 218980
rect 571852 218968 571858 219020
rect 574738 218968 574744 219020
rect 574796 219008 574802 219020
rect 586514 219008 586520 219020
rect 574796 218980 586520 219008
rect 574796 218968 574802 218980
rect 586514 218968 586520 218980
rect 586572 218968 586578 219020
rect 572898 218940 572904 218952
rect 558196 218912 558408 218940
rect 571996 218912 572904 218940
rect 558196 218872 558224 218912
rect 557828 218844 558224 218872
rect 559742 218832 559748 218884
rect 559800 218872 559806 218884
rect 567838 218872 567844 218884
rect 559800 218844 567844 218872
rect 559800 218832 559806 218844
rect 567838 218832 567844 218844
rect 567896 218832 567902 218884
rect 568022 218832 568028 218884
rect 568080 218872 568086 218884
rect 571996 218872 572024 218912
rect 572898 218900 572904 218912
rect 572956 218900 572962 218952
rect 568080 218844 572024 218872
rect 568080 218832 568086 218844
rect 573082 218832 573088 218884
rect 573140 218872 573146 218884
rect 591666 218872 591672 218884
rect 573140 218844 591672 218872
rect 573140 218832 573146 218844
rect 591666 218832 591672 218844
rect 591724 218832 591730 218884
rect 548444 218708 548564 218736
rect 544470 218600 544476 218612
rect 509896 218572 514754 218600
rect 524386 218572 544476 218600
rect 174780 218436 186314 218464
rect 174780 218424 174786 218436
rect 186498 218424 186504 218476
rect 186556 218464 186562 218476
rect 235166 218464 235172 218476
rect 186556 218436 235172 218464
rect 186556 218424 186562 218436
rect 235166 218424 235172 218436
rect 235224 218424 235230 218476
rect 239490 218424 239496 218476
rect 239548 218464 239554 218476
rect 272426 218464 272432 218476
rect 239548 218436 272432 218464
rect 239548 218424 239554 218436
rect 272426 218424 272432 218436
rect 272484 218424 272490 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 281074 218464 281080 218476
rect 279292 218436 281080 218464
rect 279292 218424 279298 218436
rect 281074 218424 281080 218436
rect 281132 218424 281138 218476
rect 285858 218424 285864 218476
rect 285916 218464 285922 218476
rect 306742 218464 306748 218476
rect 285916 218436 306748 218464
rect 285916 218424 285922 218436
rect 306742 218424 306748 218436
rect 306800 218424 306806 218476
rect 482922 218424 482928 218476
rect 482980 218464 482986 218476
rect 485314 218464 485320 218476
rect 482980 218436 485320 218464
rect 482980 218424 482986 218436
rect 485314 218424 485320 218436
rect 485372 218424 485378 218476
rect 501046 218424 501052 218476
rect 501104 218464 501110 218476
rect 509896 218464 509924 218572
rect 501104 218436 509924 218464
rect 501104 218424 501110 218436
rect 510338 218424 510344 218476
rect 510396 218464 510402 218476
rect 524386 218464 524414 218572
rect 544470 218560 544476 218572
rect 544528 218560 544534 218612
rect 548536 218600 548564 218708
rect 548702 218696 548708 218748
rect 548760 218736 548766 218748
rect 555786 218736 555792 218748
rect 548760 218708 555792 218736
rect 548760 218696 548766 218708
rect 555786 218696 555792 218708
rect 555844 218696 555850 218748
rect 555988 218708 558868 218736
rect 555988 218600 556016 218708
rect 548536 218572 556016 218600
rect 556154 218560 556160 218612
rect 556212 218600 556218 218612
rect 558546 218600 558552 218612
rect 556212 218572 558552 218600
rect 556212 218560 556218 218572
rect 558546 218560 558552 218572
rect 558604 218560 558610 218612
rect 558840 218600 558868 218708
rect 559098 218696 559104 218748
rect 559156 218736 559162 218748
rect 562870 218736 562876 218748
rect 559156 218708 562876 218736
rect 559156 218696 559162 218708
rect 562870 218696 562876 218708
rect 562928 218696 562934 218748
rect 563054 218696 563060 218748
rect 563112 218736 563118 218748
rect 572070 218736 572076 218748
rect 563112 218708 572076 218736
rect 563112 218696 563118 218708
rect 572070 218696 572076 218708
rect 572128 218696 572134 218748
rect 572438 218696 572444 218748
rect 572496 218736 572502 218748
rect 575106 218736 575112 218748
rect 572496 218708 575112 218736
rect 572496 218696 572502 218708
rect 575106 218696 575112 218708
rect 575164 218696 575170 218748
rect 582190 218696 582196 218748
rect 582248 218736 582254 218748
rect 586330 218736 586336 218748
rect 582248 218708 586336 218736
rect 582248 218696 582254 218708
rect 586330 218696 586336 218708
rect 586388 218696 586394 218748
rect 562870 218600 562876 218612
rect 558840 218572 562876 218600
rect 562870 218560 562876 218572
rect 562928 218560 562934 218612
rect 567010 218600 567016 218612
rect 563348 218572 567016 218600
rect 510396 218436 524414 218464
rect 510396 218424 510402 218436
rect 527542 218424 527548 218476
rect 527600 218464 527606 218476
rect 563348 218464 563376 218572
rect 567010 218560 567016 218572
rect 567068 218560 567074 218612
rect 567194 218560 567200 218612
rect 567252 218600 567258 218612
rect 597462 218600 597468 218612
rect 567252 218572 572208 218600
rect 567252 218560 567258 218572
rect 527600 218436 563376 218464
rect 527600 218424 527606 218436
rect 563514 218424 563520 218476
rect 563572 218464 563578 218476
rect 572180 218464 572208 218572
rect 572640 218572 597468 218600
rect 572640 218464 572668 218572
rect 597462 218560 597468 218572
rect 597520 218560 597526 218612
rect 573450 218464 573456 218476
rect 563572 218436 572116 218464
rect 572180 218436 572668 218464
rect 572732 218436 573456 218464
rect 563572 218424 563578 218436
rect 75546 218288 75552 218340
rect 75604 218328 75610 218340
rect 83458 218328 83464 218340
rect 75604 218300 83464 218328
rect 75604 218288 75610 218300
rect 83458 218288 83464 218300
rect 83516 218288 83522 218340
rect 100386 218288 100392 218340
rect 100444 218328 100450 218340
rect 105814 218328 105820 218340
rect 100444 218300 105820 218328
rect 100444 218288 100450 218300
rect 105814 218288 105820 218300
rect 105872 218288 105878 218340
rect 107010 218288 107016 218340
rect 107068 218328 107074 218340
rect 149054 218328 149060 218340
rect 107068 218300 149060 218328
rect 107068 218288 107074 218300
rect 149054 218288 149060 218300
rect 149112 218288 149118 218340
rect 149238 218288 149244 218340
rect 149296 218328 149302 218340
rect 150342 218328 150348 218340
rect 149296 218300 150348 218328
rect 149296 218288 149302 218300
rect 150342 218288 150348 218300
rect 150400 218288 150406 218340
rect 150526 218288 150532 218340
rect 150584 218328 150590 218340
rect 157242 218328 157248 218340
rect 150584 218300 157248 218328
rect 150584 218288 150590 218300
rect 157242 218288 157248 218300
rect 157300 218288 157306 218340
rect 159818 218328 159824 218340
rect 157536 218300 159824 218328
rect 56318 218152 56324 218204
rect 56376 218192 56382 218204
rect 62758 218192 62764 218204
rect 56376 218164 62764 218192
rect 56376 218152 56382 218164
rect 62758 218152 62764 218164
rect 62816 218152 62822 218204
rect 79686 218152 79692 218204
rect 79744 218192 79750 218204
rect 82078 218192 82084 218204
rect 79744 218164 82084 218192
rect 79744 218152 79750 218164
rect 82078 218152 82084 218164
rect 82136 218152 82142 218204
rect 119982 218152 119988 218204
rect 120040 218192 120046 218204
rect 157536 218192 157564 218300
rect 159818 218288 159824 218300
rect 159876 218288 159882 218340
rect 160002 218288 160008 218340
rect 160060 218328 160066 218340
rect 162670 218328 162676 218340
rect 160060 218300 162676 218328
rect 160060 218288 160066 218300
rect 162670 218288 162676 218300
rect 162728 218288 162734 218340
rect 162854 218288 162860 218340
rect 162912 218328 162918 218340
rect 166442 218328 166448 218340
rect 162912 218300 166448 218328
rect 162912 218288 162918 218300
rect 166442 218288 166448 218300
rect 166500 218288 166506 218340
rect 166626 218288 166632 218340
rect 166684 218328 166690 218340
rect 213546 218328 213552 218340
rect 166684 218300 213552 218328
rect 166684 218288 166690 218300
rect 213546 218288 213552 218300
rect 213604 218288 213610 218340
rect 216306 218288 216312 218340
rect 216364 218328 216370 218340
rect 221642 218328 221648 218340
rect 216364 218300 221648 218328
rect 216364 218288 216370 218300
rect 221642 218288 221648 218300
rect 221700 218288 221706 218340
rect 224586 218288 224592 218340
rect 224644 218328 224650 218340
rect 225598 218328 225604 218340
rect 224644 218300 225604 218328
rect 224644 218288 224650 218300
rect 225598 218288 225604 218300
rect 225656 218288 225662 218340
rect 227898 218288 227904 218340
rect 227956 218328 227962 218340
rect 229186 218328 229192 218340
rect 227956 218300 229192 218328
rect 227956 218288 227962 218300
rect 229186 218288 229192 218300
rect 229244 218288 229250 218340
rect 244458 218288 244464 218340
rect 244516 218328 244522 218340
rect 247678 218328 247684 218340
rect 244516 218300 247684 218328
rect 244516 218288 244522 218300
rect 247678 218288 247684 218300
rect 247736 218288 247742 218340
rect 365346 218288 365352 218340
rect 365404 218328 365410 218340
rect 373258 218328 373264 218340
rect 365404 218300 373264 218328
rect 365404 218288 365410 218300
rect 373258 218288 373264 218300
rect 373316 218288 373322 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429562 218328 429568 218340
rect 426676 218300 429568 218328
rect 426676 218288 426682 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 475562 218288 475568 218340
rect 475620 218328 475626 218340
rect 482830 218328 482836 218340
rect 475620 218300 482836 218328
rect 475620 218288 475626 218300
rect 482830 218288 482836 218300
rect 482888 218288 482894 218340
rect 500034 218288 500040 218340
rect 500092 218328 500098 218340
rect 507118 218328 507124 218340
rect 500092 218300 507124 218328
rect 500092 218288 500098 218300
rect 507118 218288 507124 218300
rect 507176 218288 507182 218340
rect 507670 218288 507676 218340
rect 507728 218328 507734 218340
rect 507728 218300 529244 218328
rect 507728 218288 507734 218300
rect 120040 218164 157564 218192
rect 120040 218152 120046 218164
rect 157702 218152 157708 218204
rect 157760 218192 157766 218204
rect 161290 218192 161296 218204
rect 157760 218164 161296 218192
rect 157760 218152 157766 218164
rect 161290 218152 161296 218164
rect 161348 218152 161354 218204
rect 162118 218152 162124 218204
rect 162176 218192 162182 218204
rect 167638 218192 167644 218204
rect 162176 218164 167644 218192
rect 162176 218152 162182 218164
rect 167638 218152 167644 218164
rect 167696 218152 167702 218204
rect 168098 218152 168104 218204
rect 168156 218192 168162 218204
rect 171042 218192 171048 218204
rect 168156 218164 171048 218192
rect 168156 218152 168162 218164
rect 171042 218152 171048 218164
rect 171100 218152 171106 218204
rect 171594 218152 171600 218204
rect 171652 218192 171658 218204
rect 171652 218164 175412 218192
rect 171652 218152 171658 218164
rect 55674 218016 55680 218068
rect 55732 218056 55738 218068
rect 56502 218056 56508 218068
rect 55732 218028 56508 218056
rect 55732 218016 55738 218028
rect 56502 218016 56508 218028
rect 56560 218016 56566 218068
rect 57330 218016 57336 218068
rect 57388 218056 57394 218068
rect 57882 218056 57888 218068
rect 57388 218028 57888 218056
rect 57388 218016 57394 218028
rect 57882 218016 57888 218028
rect 57940 218016 57946 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 61286 218056 61292 218068
rect 58216 218028 61292 218056
rect 58216 218016 58222 218028
rect 61286 218016 61292 218028
rect 61344 218016 61350 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 73890 218016 73896 218068
rect 73948 218056 73954 218068
rect 74442 218056 74448 218068
rect 73948 218028 74448 218056
rect 73948 218016 73954 218028
rect 74442 218016 74448 218028
rect 74500 218016 74506 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 82722 218056 82728 218068
rect 82228 218028 82728 218056
rect 82228 218016 82234 218028
rect 82722 218016 82728 218028
rect 82780 218016 82786 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85482 218056 85488 218068
rect 84712 218028 85488 218056
rect 84712 218016 84718 218028
rect 85482 218016 85488 218028
rect 85540 218016 85546 218068
rect 86310 218016 86316 218068
rect 86368 218056 86374 218068
rect 86862 218056 86868 218068
rect 86368 218028 86868 218056
rect 86368 218016 86374 218028
rect 86862 218016 86868 218028
rect 86920 218016 86926 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 94590 218016 94596 218068
rect 94648 218056 94654 218068
rect 95142 218056 95148 218068
rect 94648 218028 95148 218056
rect 94648 218016 94654 218028
rect 95142 218016 95148 218028
rect 95200 218016 95206 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 101214 218016 101220 218068
rect 101272 218056 101278 218068
rect 102134 218056 102140 218068
rect 101272 218028 102140 218056
rect 101272 218016 101278 218028
rect 102134 218016 102140 218028
rect 102192 218016 102198 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 103698 218016 103704 218068
rect 103756 218056 103762 218068
rect 104802 218056 104808 218068
rect 103756 218028 104808 218056
rect 103756 218016 103762 218028
rect 104802 218016 104808 218028
rect 104860 218016 104866 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 110322 218016 110328 218068
rect 110380 218056 110386 218068
rect 110966 218056 110972 218068
rect 110380 218028 110972 218056
rect 110380 218016 110386 218028
rect 110966 218016 110972 218028
rect 111024 218016 111030 218068
rect 111978 218016 111984 218068
rect 112036 218056 112042 218068
rect 112806 218056 112812 218068
rect 112036 218028 112812 218056
rect 112036 218016 112042 218028
rect 112806 218016 112812 218028
rect 112864 218016 112870 218068
rect 115290 218016 115296 218068
rect 115348 218056 115354 218068
rect 115750 218056 115756 218068
rect 115348 218028 115756 218056
rect 115348 218016 115354 218028
rect 115750 218016 115756 218028
rect 115808 218016 115814 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 120258 218016 120264 218068
rect 120316 218056 120322 218068
rect 162854 218056 162860 218068
rect 120316 218028 162860 218056
rect 120316 218016 120322 218028
rect 162854 218016 162860 218028
rect 162912 218016 162918 218068
rect 163314 218016 163320 218068
rect 163372 218056 163378 218068
rect 163372 218028 164234 218056
rect 163372 218016 163378 218028
rect 164206 217920 164234 218028
rect 167454 218016 167460 218068
rect 167512 218056 167518 218068
rect 168282 218056 168288 218068
rect 167512 218028 168288 218056
rect 167512 218016 167518 218028
rect 168282 218016 168288 218028
rect 168340 218016 168346 218068
rect 169110 218016 169116 218068
rect 169168 218056 169174 218068
rect 169570 218056 169576 218068
rect 169168 218028 169576 218056
rect 169168 218016 169174 218028
rect 169570 218016 169576 218028
rect 169628 218016 169634 218068
rect 173250 218016 173256 218068
rect 173308 218056 173314 218068
rect 173308 218028 173940 218056
rect 173308 218016 173314 218028
rect 169294 217920 169300 217932
rect 164206 217892 169300 217920
rect 169294 217880 169300 217892
rect 169352 217880 169358 217932
rect 173912 217920 173940 218028
rect 174078 218016 174084 218068
rect 174136 218056 174142 218068
rect 175182 218056 175188 218068
rect 174136 218028 175188 218056
rect 174136 218016 174142 218028
rect 175182 218016 175188 218028
rect 175240 218016 175246 218068
rect 175384 218056 175412 218164
rect 175734 218152 175740 218204
rect 175792 218192 175798 218204
rect 176470 218192 176476 218204
rect 175792 218164 176476 218192
rect 175792 218152 175798 218164
rect 176470 218152 176476 218164
rect 176528 218152 176534 218204
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 221090 218192 221096 218204
rect 179932 218164 221096 218192
rect 179932 218152 179938 218164
rect 221090 218152 221096 218164
rect 221148 218152 221154 218204
rect 221274 218152 221280 218204
rect 221332 218192 221338 218204
rect 221826 218192 221832 218204
rect 221332 218164 221832 218192
rect 221332 218152 221338 218164
rect 221826 218152 221832 218164
rect 221884 218152 221890 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 223390 218192 223396 218204
rect 222988 218164 223396 218192
rect 222988 218152 222994 218164
rect 223390 218152 223396 218164
rect 223448 218152 223454 218204
rect 223758 218152 223764 218204
rect 223816 218192 223822 218204
rect 224862 218192 224868 218204
rect 223816 218164 224868 218192
rect 223816 218152 223822 218164
rect 224862 218152 224868 218164
rect 224920 218152 224926 218204
rect 225414 218152 225420 218204
rect 225472 218192 225478 218204
rect 226150 218192 226156 218204
rect 225472 218164 226156 218192
rect 225472 218152 225478 218164
rect 226150 218152 226156 218164
rect 226208 218152 226214 218204
rect 229554 218152 229560 218204
rect 229612 218192 229618 218204
rect 231026 218192 231032 218204
rect 229612 218164 231032 218192
rect 229612 218152 229618 218164
rect 231026 218152 231032 218164
rect 231084 218152 231090 218204
rect 231210 218152 231216 218204
rect 231268 218192 231274 218204
rect 231670 218192 231676 218204
rect 231268 218164 231676 218192
rect 231268 218152 231274 218164
rect 231670 218152 231676 218164
rect 231728 218152 231734 218204
rect 232038 218152 232044 218204
rect 232096 218192 232102 218204
rect 233142 218192 233148 218204
rect 232096 218164 233148 218192
rect 232096 218152 232102 218164
rect 233142 218152 233148 218164
rect 233200 218152 233206 218204
rect 235350 218152 235356 218204
rect 235408 218192 235414 218204
rect 235902 218192 235908 218204
rect 235408 218164 235908 218192
rect 235408 218152 235414 218164
rect 235902 218152 235908 218164
rect 235960 218152 235966 218204
rect 236178 218152 236184 218204
rect 236236 218192 236242 218204
rect 236914 218192 236920 218204
rect 236236 218164 236920 218192
rect 236236 218152 236242 218164
rect 236914 218152 236920 218164
rect 236972 218152 236978 218204
rect 249058 218192 249064 218204
rect 238726 218164 249064 218192
rect 176286 218056 176292 218068
rect 175384 218028 176292 218056
rect 176286 218016 176292 218028
rect 176344 218016 176350 218068
rect 176562 218016 176568 218068
rect 176620 218056 176626 218068
rect 177574 218056 177580 218068
rect 176620 218028 177580 218056
rect 176620 218016 176626 218028
rect 177574 218016 177580 218028
rect 177632 218016 177638 218068
rect 189810 218016 189816 218068
rect 189868 218056 189874 218068
rect 190270 218056 190276 218068
rect 189868 218028 190276 218056
rect 189868 218016 189874 218028
rect 190270 218016 190276 218028
rect 190328 218016 190334 218068
rect 192110 218056 192116 218068
rect 190426 218028 192116 218056
rect 174722 217920 174728 217932
rect 173912 217892 174728 217920
rect 174722 217880 174728 217892
rect 174780 217880 174786 217932
rect 190086 217880 190092 217932
rect 190144 217920 190150 217932
rect 190426 217920 190454 218028
rect 192110 218016 192116 218028
rect 192168 218016 192174 218068
rect 192294 218016 192300 218068
rect 192352 218056 192358 218068
rect 192938 218056 192944 218068
rect 192352 218028 192944 218056
rect 192352 218016 192358 218028
rect 192938 218016 192944 218028
rect 192996 218016 193002 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 196434 218016 196440 218068
rect 196492 218056 196498 218068
rect 197078 218056 197084 218068
rect 196492 218028 197084 218056
rect 196492 218016 196498 218028
rect 197078 218016 197084 218028
rect 197136 218016 197142 218068
rect 198918 218016 198924 218068
rect 198976 218056 198982 218068
rect 200022 218056 200028 218068
rect 198976 218028 200028 218056
rect 198976 218016 198982 218028
rect 200022 218016 200028 218028
rect 200080 218016 200086 218068
rect 202230 218016 202236 218068
rect 202288 218056 202294 218068
rect 202690 218056 202696 218068
rect 202288 218028 202696 218056
rect 202288 218016 202294 218028
rect 202690 218016 202696 218028
rect 202748 218016 202754 218068
rect 203058 218016 203064 218068
rect 203116 218056 203122 218068
rect 203702 218056 203708 218068
rect 203116 218028 203708 218056
rect 203116 218016 203122 218028
rect 203702 218016 203708 218028
rect 203760 218016 203766 218068
rect 204714 218016 204720 218068
rect 204772 218056 204778 218068
rect 206002 218056 206008 218068
rect 204772 218028 206008 218056
rect 204772 218016 204778 218028
rect 206002 218016 206008 218028
rect 206060 218016 206066 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 212994 218016 213000 218068
rect 213052 218056 213058 218068
rect 213052 218028 215340 218056
rect 213052 218016 213058 218028
rect 190144 217892 190454 217920
rect 215312 217920 215340 218028
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216490 218056 216496 218068
rect 215536 218028 216496 218056
rect 215536 218016 215542 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 238726 218056 238754 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251726 218192 251732 218204
rect 249484 218164 251732 218192
rect 249484 218152 249490 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 269298 218152 269304 218204
rect 269356 218192 269362 218204
rect 273898 218192 273904 218204
rect 269356 218164 273904 218192
rect 269356 218152 269362 218164
rect 273898 218152 273904 218164
rect 273956 218152 273962 218204
rect 299106 218152 299112 218204
rect 299164 218192 299170 218204
rect 300302 218192 300308 218204
rect 299164 218164 300308 218192
rect 299164 218152 299170 218164
rect 300302 218152 300308 218164
rect 300360 218152 300366 218204
rect 302418 218152 302424 218204
rect 302476 218192 302482 218204
rect 304626 218192 304632 218204
rect 302476 218164 304632 218192
rect 302476 218152 302482 218164
rect 304626 218152 304632 218164
rect 304684 218152 304690 218204
rect 310698 218152 310704 218204
rect 310756 218192 310762 218204
rect 315298 218192 315304 218204
rect 310756 218164 315304 218192
rect 310756 218152 310762 218164
rect 315298 218152 315304 218164
rect 315356 218152 315362 218204
rect 330662 218152 330668 218204
rect 330720 218192 330726 218204
rect 333238 218192 333244 218204
rect 330720 218164 333244 218192
rect 330720 218152 330726 218164
rect 333238 218152 333244 218164
rect 333296 218152 333302 218204
rect 348786 218152 348792 218204
rect 348844 218192 348850 218204
rect 351178 218192 351184 218204
rect 348844 218164 351184 218192
rect 348844 218152 348850 218164
rect 351178 218152 351184 218164
rect 351236 218152 351242 218204
rect 364518 218152 364524 218204
rect 364576 218192 364582 218204
rect 367646 218192 367652 218204
rect 364576 218164 367652 218192
rect 364576 218152 364582 218164
rect 367646 218152 367652 218164
rect 367704 218152 367710 218204
rect 369486 218152 369492 218204
rect 369544 218192 369550 218204
rect 370498 218192 370504 218204
rect 369544 218164 370504 218192
rect 369544 218152 369550 218164
rect 370498 218152 370504 218164
rect 370556 218152 370562 218204
rect 376938 218152 376944 218204
rect 376996 218192 377002 218204
rect 382918 218192 382924 218204
rect 376996 218164 382924 218192
rect 376996 218152 377002 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 386874 218152 386880 218204
rect 386932 218192 386938 218204
rect 388438 218192 388444 218204
rect 386932 218164 388444 218192
rect 386932 218152 386938 218164
rect 388438 218152 388444 218164
rect 388496 218152 388502 218204
rect 394326 218152 394332 218204
rect 394384 218192 394390 218204
rect 402238 218192 402244 218204
rect 394384 218164 402244 218192
rect 394384 218152 394390 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 427906 218192 427912 218204
rect 425848 218164 427912 218192
rect 425848 218152 425854 218164
rect 427906 218152 427912 218164
rect 427964 218152 427970 218204
rect 428458 218152 428464 218204
rect 428516 218192 428522 218204
rect 430114 218192 430120 218204
rect 428516 218164 430120 218192
rect 428516 218152 428522 218164
rect 430114 218152 430120 218164
rect 430172 218152 430178 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 435726 218152 435732 218204
rect 435784 218192 435790 218204
rect 436646 218192 436652 218204
rect 435784 218164 436652 218192
rect 435784 218152 435790 218164
rect 436646 218152 436652 218164
rect 436704 218152 436710 218204
rect 455046 218152 455052 218204
rect 455104 218192 455110 218204
rect 460474 218192 460480 218204
rect 455104 218164 460480 218192
rect 455104 218152 455110 218164
rect 460474 218152 460480 218164
rect 460532 218152 460538 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 494606 218152 494612 218204
rect 494664 218192 494670 218204
rect 495250 218192 495256 218204
rect 494664 218164 495256 218192
rect 494664 218152 494670 218164
rect 495250 218152 495256 218164
rect 495308 218192 495314 218204
rect 519538 218192 519544 218204
rect 495308 218164 519544 218192
rect 495308 218152 495314 218164
rect 519538 218152 519544 218164
rect 519596 218152 519602 218204
rect 519814 218152 519820 218204
rect 519872 218192 519878 218204
rect 524414 218192 524420 218204
rect 519872 218164 524420 218192
rect 519872 218152 519878 218164
rect 524414 218152 524420 218164
rect 524472 218152 524478 218204
rect 529216 218192 529244 218300
rect 529382 218288 529388 218340
rect 529440 218328 529446 218340
rect 571886 218328 571892 218340
rect 529440 218300 571892 218328
rect 529440 218288 529446 218300
rect 571886 218288 571892 218300
rect 571944 218288 571950 218340
rect 572088 218328 572116 218436
rect 572732 218328 572760 218436
rect 573450 218424 573456 218436
rect 573508 218424 573514 218476
rect 573634 218424 573640 218476
rect 573692 218464 573698 218476
rect 606478 218464 606484 218476
rect 573692 218436 606484 218464
rect 573692 218424 573698 218436
rect 606478 218424 606484 218436
rect 606536 218424 606542 218476
rect 572088 218300 572760 218328
rect 573266 218288 573272 218340
rect 573324 218328 573330 218340
rect 574370 218328 574376 218340
rect 573324 218300 574376 218328
rect 573324 218288 573330 218300
rect 574370 218288 574376 218300
rect 574428 218288 574434 218340
rect 574554 218288 574560 218340
rect 574612 218328 574618 218340
rect 605282 218328 605288 218340
rect 574612 218300 605288 218328
rect 574612 218288 574618 218300
rect 605282 218288 605288 218300
rect 605340 218288 605346 218340
rect 548702 218192 548708 218204
rect 529216 218164 548708 218192
rect 548702 218152 548708 218164
rect 548760 218152 548766 218204
rect 548886 218152 548892 218204
rect 548944 218192 548950 218204
rect 553486 218192 553492 218204
rect 548944 218164 553492 218192
rect 548944 218152 548950 218164
rect 553486 218152 553492 218164
rect 553544 218152 553550 218204
rect 553670 218152 553676 218204
rect 553728 218192 553734 218204
rect 553728 218164 560432 218192
rect 553728 218152 553734 218164
rect 560404 218124 560432 218164
rect 563330 218152 563336 218204
rect 563388 218192 563394 218204
rect 571978 218192 571984 218204
rect 563388 218164 571984 218192
rect 563388 218152 563394 218164
rect 571978 218152 571984 218164
rect 572036 218152 572042 218204
rect 572162 218152 572168 218204
rect 572220 218192 572226 218204
rect 574922 218192 574928 218204
rect 572220 218164 574928 218192
rect 572220 218152 572226 218164
rect 574922 218152 574928 218164
rect 574980 218152 574986 218204
rect 586330 218152 586336 218204
rect 586388 218192 586394 218204
rect 594978 218192 594984 218204
rect 586388 218164 594984 218192
rect 586388 218152 586394 218164
rect 594978 218152 594984 218164
rect 595036 218152 595042 218204
rect 596910 218152 596916 218204
rect 596968 218192 596974 218204
rect 601326 218192 601332 218204
rect 596968 218164 601332 218192
rect 596968 218152 596974 218164
rect 601326 218152 601332 218164
rect 601384 218152 601390 218204
rect 563008 218124 563014 218136
rect 560404 218096 563014 218124
rect 563008 218084 563014 218096
rect 563066 218084 563072 218136
rect 216692 218028 238754 218056
rect 216692 217920 216720 218028
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249702 218056 249708 218068
rect 248656 218028 249708 218056
rect 248656 218016 248662 218028
rect 249702 218016 249708 218028
rect 249760 218016 249766 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 251174 218056 251180 218068
rect 250312 218028 251180 218056
rect 250312 218016 250318 218028
rect 251174 218016 251180 218028
rect 251232 218016 251238 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 262674 218016 262680 218068
rect 262732 218056 262738 218068
rect 263594 218056 263600 218068
rect 262732 218028 263600 218056
rect 262732 218016 262738 218028
rect 263594 218016 263600 218028
rect 263652 218016 263658 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 266814 218016 266820 218068
rect 266872 218056 266878 218068
rect 267688 218056 267694 218068
rect 266872 218028 267694 218056
rect 266872 218016 266878 218028
rect 267688 218016 267694 218028
rect 267746 218016 267752 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 269022 218056 269028 218068
rect 268528 218028 269028 218056
rect 268528 218016 268534 218028
rect 269022 218016 269028 218028
rect 269080 218016 269086 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 271598 218056 271604 218068
rect 271012 218028 271604 218056
rect 271012 218016 271018 218028
rect 271598 218016 271604 218028
rect 271656 218016 271662 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278498 218056 278504 218068
rect 277636 218028 278504 218056
rect 277636 218016 277642 218028
rect 278498 218016 278504 218028
rect 278556 218016 278562 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282546 218056 282552 218068
rect 281776 218028 282552 218056
rect 281776 218016 281782 218028
rect 282546 218016 282552 218028
rect 282604 218016 282610 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289630 218056 289636 218068
rect 289228 218028 289636 218056
rect 289228 218016 289234 218028
rect 289630 218016 289636 218028
rect 289688 218016 289694 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 295794 218016 295800 218068
rect 295852 218056 295858 218068
rect 296438 218056 296444 218068
rect 295852 218028 296444 218056
rect 295852 218016 295858 218028
rect 296438 218016 296444 218028
rect 296496 218016 296502 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 298002 218056 298008 218068
rect 297508 218028 298008 218056
rect 297508 218016 297514 218028
rect 298002 218016 298008 218028
rect 298060 218016 298066 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299290 218056 299296 218068
rect 298336 218028 299296 218056
rect 298336 218016 298342 218028
rect 299290 218016 299296 218028
rect 299348 218016 299354 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 305546 218056 305552 218068
rect 304132 218028 305552 218056
rect 304132 218016 304138 218028
rect 305546 218016 305552 218028
rect 305604 218016 305610 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306282 218056 306288 218068
rect 305788 218028 306288 218056
rect 305788 218016 305794 218028
rect 306282 218016 306288 218028
rect 306340 218016 306346 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308766 218056 308772 218068
rect 308272 218028 308772 218056
rect 308272 218016 308278 218028
rect 308766 218016 308772 218028
rect 308824 218016 308830 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 314562 218056 314568 218068
rect 312412 218028 314568 218056
rect 312412 218016 312418 218028
rect 314562 218016 314568 218028
rect 314620 218016 314626 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315850 218056 315856 218068
rect 314896 218028 315856 218056
rect 314896 218016 314902 218028
rect 315850 218016 315856 218028
rect 315908 218016 315914 218068
rect 316494 218016 316500 218068
rect 316552 218056 316558 218068
rect 317138 218056 317144 218068
rect 316552 218028 317144 218056
rect 316552 218016 316558 218028
rect 317138 218016 317144 218028
rect 317196 218016 317202 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319990 218056 319996 218068
rect 319036 218028 319996 218056
rect 319036 218016 319042 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 328914 218016 328920 218068
rect 328972 218056 328978 218068
rect 330478 218056 330484 218068
rect 328972 218028 330484 218056
rect 328972 218016 328978 218028
rect 330478 218016 330484 218028
rect 330536 218016 330542 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335262 218056 335268 218068
rect 334768 218028 335268 218056
rect 334768 218016 334774 218028
rect 335262 218016 335268 218028
rect 335320 218016 335326 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 336366 218056 336372 218068
rect 335596 218028 336372 218056
rect 335596 218016 335602 218028
rect 336366 218016 336372 218028
rect 336424 218016 336430 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 342990 218016 342996 218068
rect 343048 218056 343054 218068
rect 343542 218056 343548 218068
rect 343048 218028 343548 218056
rect 343048 218016 343054 218028
rect 343542 218016 343548 218028
rect 343600 218016 343606 218068
rect 347130 218016 347136 218068
rect 347188 218056 347194 218068
rect 347590 218056 347596 218068
rect 347188 218028 347596 218056
rect 347188 218016 347194 218028
rect 347590 218016 347596 218028
rect 347648 218016 347654 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 353754 218016 353760 218068
rect 353812 218056 353818 218068
rect 354582 218056 354588 218068
rect 353812 218028 354588 218056
rect 353812 218016 353818 218028
rect 354582 218016 354588 218028
rect 354640 218016 354646 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357342 218056 357348 218068
rect 356296 218028 357348 218056
rect 356296 218016 356302 218028
rect 357342 218016 357348 218028
rect 357400 218016 357406 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 359366 218056 359372 218068
rect 357952 218028 359372 218056
rect 357952 218016 357958 218028
rect 359366 218016 359372 218028
rect 359424 218016 359430 218068
rect 363690 218016 363696 218068
rect 363748 218056 363754 218068
rect 364150 218056 364156 218068
rect 363748 218028 364156 218056
rect 363748 218016 363754 218028
rect 364150 218016 364156 218028
rect 364208 218016 364214 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366910 218056 366916 218068
rect 366232 218028 366916 218056
rect 366232 218016 366238 218028
rect 366910 218016 366916 218028
rect 366968 218016 366974 218068
rect 368658 218016 368664 218068
rect 368716 218056 368722 218068
rect 369762 218056 369768 218068
rect 368716 218028 369768 218056
rect 368716 218016 368722 218028
rect 369762 218016 369768 218028
rect 369820 218016 369826 218068
rect 370314 218016 370320 218068
rect 370372 218056 370378 218068
rect 370958 218056 370964 218068
rect 370372 218028 370964 218056
rect 370372 218016 370378 218028
rect 370958 218016 370964 218028
rect 371016 218016 371022 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373810 218056 373816 218068
rect 372856 218028 373816 218056
rect 372856 218016 372862 218028
rect 373810 218016 373816 218028
rect 373868 218016 373874 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376570 218056 376576 218068
rect 376168 218028 376576 218056
rect 376168 218016 376174 218028
rect 376570 218016 376576 218028
rect 376628 218016 376634 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379330 218056 379336 218068
rect 378652 218028 379336 218056
rect 378652 218016 378658 218028
rect 379330 218016 379336 218028
rect 379388 218016 379394 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 381722 218056 381728 218068
rect 381136 218028 381728 218056
rect 381136 218016 381142 218028
rect 381722 218016 381728 218028
rect 381780 218016 381786 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386322 218056 386328 218068
rect 385276 218028 386328 218056
rect 385276 218016 385282 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 388530 218016 388536 218068
rect 388588 218056 388594 218068
rect 389082 218056 389088 218068
rect 388588 218028 389088 218056
rect 388588 218016 388594 218028
rect 389082 218016 389088 218028
rect 389140 218016 389146 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390278 218056 390284 218068
rect 389416 218028 390284 218056
rect 389416 218016 389422 218028
rect 390278 218016 390284 218028
rect 390336 218016 390342 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393222 218056 393228 218068
rect 392728 218028 393228 218056
rect 392728 218016 392734 218028
rect 393222 218016 393228 218028
rect 393280 218016 393286 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394602 218056 394608 218068
rect 393556 218028 394608 218056
rect 393556 218016 393562 218028
rect 394602 218016 394608 218028
rect 394660 218016 394666 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395982 218056 395988 218068
rect 395212 218028 395988 218056
rect 395212 218016 395218 218028
rect 395982 218016 395988 218028
rect 396040 218016 396046 218068
rect 396810 218016 396816 218068
rect 396868 218056 396874 218068
rect 397362 218056 397368 218068
rect 396868 218028 397368 218056
rect 396868 218016 396874 218028
rect 397362 218016 397368 218028
rect 397420 218016 397426 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 401410 218056 401416 218068
rect 401008 218028 401416 218056
rect 401008 218016 401014 218028
rect 401410 218016 401416 218028
rect 401468 218016 401474 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 418338 218016 418344 218068
rect 418396 218056 418402 218068
rect 419442 218056 419448 218068
rect 418396 218028 419448 218056
rect 418396 218016 418402 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 428274 218056 428280 218068
rect 427504 218028 428280 218056
rect 427504 218016 427510 218028
rect 428274 218016 428280 218028
rect 428332 218016 428338 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434898 218016 434904 218068
rect 434956 218056 434962 218068
rect 436278 218056 436284 218068
rect 434956 218028 436284 218056
rect 434956 218016 434962 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437750 218056 437756 218068
rect 436612 218028 437756 218056
rect 436612 218016 436618 218028
rect 437750 218016 437756 218028
rect 437808 218016 437814 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455506 218056 455512 218068
rect 453356 218028 455512 218056
rect 453356 218016 453362 218028
rect 455506 218016 455512 218028
rect 455564 218016 455570 218068
rect 456702 218016 456708 218068
rect 456760 218056 456766 218068
rect 457162 218056 457168 218068
rect 456760 218028 457168 218056
rect 456760 218016 456766 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 471698 218016 471704 218068
rect 471756 218056 471762 218068
rect 472894 218056 472900 218068
rect 471756 218028 472900 218056
rect 471756 218016 471762 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 488718 218016 488724 218068
rect 488776 218056 488782 218068
rect 497550 218056 497556 218068
rect 488776 218028 497556 218056
rect 488776 218016 488782 218028
rect 497550 218016 497556 218028
rect 497608 218016 497614 218068
rect 505278 218016 505284 218068
rect 505336 218056 505342 218068
rect 505646 218056 505652 218068
rect 505336 218028 505652 218056
rect 505336 218016 505342 218028
rect 505646 218016 505652 218028
rect 505704 218056 505710 218068
rect 613838 218056 613844 218068
rect 505704 218028 553302 218056
rect 505704 218016 505710 218028
rect 553274 217988 553302 218028
rect 553596 218028 560294 218056
rect 553596 217988 553624 218028
rect 553274 217960 553624 217988
rect 560266 217988 560294 218028
rect 569926 218028 613844 218056
rect 569926 217988 569954 218028
rect 613838 218016 613844 218028
rect 613896 218016 613902 218068
rect 560266 217960 569954 217988
rect 215312 217892 216720 217920
rect 540946 217892 550634 217920
rect 190144 217880 190150 217892
rect 528370 217812 528376 217864
rect 528428 217852 528434 217864
rect 540946 217852 540974 217892
rect 528428 217824 540974 217852
rect 550606 217852 550634 217892
rect 602890 217852 602896 217864
rect 550606 217824 602896 217852
rect 528428 217812 528434 217824
rect 602890 217812 602896 217824
rect 602948 217812 602954 217864
rect 604086 217812 604092 217864
rect 604144 217852 604150 217864
rect 612274 217852 612280 217864
rect 604144 217824 612280 217852
rect 604144 217812 604150 217824
rect 612274 217812 612280 217824
rect 612332 217812 612338 217864
rect 524598 217676 524604 217728
rect 524656 217716 524662 217728
rect 524656 217688 534212 217716
rect 524656 217676 524662 217688
rect 533614 217580 533620 217592
rect 524386 217552 533620 217580
rect 523402 217472 523408 217524
rect 523460 217512 523466 217524
rect 524386 217512 524414 217552
rect 533614 217540 533620 217552
rect 533672 217540 533678 217592
rect 534184 217580 534212 217688
rect 534350 217676 534356 217728
rect 534408 217716 534414 217728
rect 542078 217716 542084 217728
rect 534408 217688 542084 217716
rect 534408 217676 534414 217688
rect 542078 217676 542084 217688
rect 542136 217676 542142 217728
rect 542262 217676 542268 217728
rect 542320 217716 542326 217728
rect 548426 217716 548432 217728
rect 542320 217688 548432 217716
rect 542320 217676 542326 217688
rect 548426 217676 548432 217688
rect 548484 217676 548490 217728
rect 596910 217716 596916 217728
rect 548628 217688 596916 217716
rect 535178 217580 535184 217592
rect 534184 217552 535184 217580
rect 535178 217540 535184 217552
rect 535236 217540 535242 217592
rect 535914 217540 535920 217592
rect 535972 217580 535978 217592
rect 535972 217552 538720 217580
rect 535972 217540 535978 217552
rect 523460 217484 524414 217512
rect 523460 217472 523466 217484
rect 538692 217444 538720 217552
rect 538858 217540 538864 217592
rect 538916 217580 538922 217592
rect 542998 217580 543004 217592
rect 538916 217552 543004 217580
rect 538916 217540 538922 217552
rect 542998 217540 543004 217552
rect 543056 217540 543062 217592
rect 548628 217512 548656 217688
rect 596910 217676 596916 217688
rect 596968 217676 596974 217728
rect 597094 217676 597100 217728
rect 597152 217716 597158 217728
rect 604454 217716 604460 217728
rect 597152 217688 604460 217716
rect 597152 217676 597158 217688
rect 604454 217676 604460 217688
rect 604512 217676 604518 217728
rect 605282 217676 605288 217728
rect 605340 217716 605346 217728
rect 615678 217716 615684 217728
rect 605340 217688 615684 217716
rect 605340 217676 605346 217688
rect 615678 217676 615684 217688
rect 615736 217676 615742 217728
rect 549438 217540 549444 217592
rect 549496 217580 549502 217592
rect 562042 217580 562048 217592
rect 549496 217552 562048 217580
rect 549496 217540 549502 217552
rect 562042 217540 562048 217552
rect 562100 217540 562106 217592
rect 562502 217540 562508 217592
rect 562560 217580 562566 217592
rect 609054 217580 609060 217592
rect 562560 217552 609060 217580
rect 562560 217540 562566 217552
rect 609054 217540 609060 217552
rect 609112 217540 609118 217592
rect 543844 217484 548656 217512
rect 542262 217444 542268 217456
rect 538692 217416 542268 217444
rect 542262 217404 542268 217416
rect 542320 217404 542326 217456
rect 543274 217404 543280 217456
rect 543332 217444 543338 217456
rect 543844 217444 543872 217484
rect 543332 217416 543872 217444
rect 543332 217404 543338 217416
rect 548794 217404 548800 217456
rect 548852 217444 548858 217456
rect 566182 217444 566188 217456
rect 548852 217416 566188 217444
rect 548852 217404 548858 217416
rect 566182 217404 566188 217416
rect 566240 217404 566246 217456
rect 567010 217404 567016 217456
rect 567068 217444 567074 217456
rect 597094 217444 597100 217456
rect 567068 217416 597100 217444
rect 567068 217404 567074 217416
rect 597094 217404 597100 217416
rect 597152 217404 597158 217456
rect 603442 217444 603448 217456
rect 597296 217416 603448 217444
rect 544010 217336 544016 217388
rect 544068 217376 544074 217388
rect 544068 217348 545068 217376
rect 544068 217336 544074 217348
rect 533430 217268 533436 217320
rect 533488 217308 533494 217320
rect 543182 217308 543188 217320
rect 533488 217280 543188 217308
rect 533488 217268 533494 217280
rect 543182 217268 543188 217280
rect 543240 217268 543246 217320
rect 545040 217308 545068 217348
rect 565262 217308 565268 217320
rect 545040 217280 565268 217308
rect 565262 217268 565268 217280
rect 565320 217268 565326 217320
rect 565814 217268 565820 217320
rect 565872 217308 565878 217320
rect 597094 217308 597100 217320
rect 565872 217280 597100 217308
rect 565872 217268 565878 217280
rect 597094 217268 597100 217280
rect 597152 217268 597158 217320
rect 145052 217200 145058 217252
rect 145110 217240 145116 217252
rect 147766 217240 147772 217252
rect 145110 217212 147772 217240
rect 145110 217200 145116 217212
rect 147766 217200 147772 217212
rect 147824 217200 147830 217252
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 543826 217200 543832 217252
rect 543884 217240 543890 217252
rect 543884 217212 544424 217240
rect 543884 217200 543890 217212
rect 530900 217132 530906 217184
rect 530958 217172 530964 217184
rect 541894 217172 541900 217184
rect 530958 217144 541900 217172
rect 530958 217132 530964 217144
rect 541894 217132 541900 217144
rect 541952 217132 541958 217184
rect 543458 217172 543464 217184
rect 543200 217144 543464 217172
rect 147536 217064 147542 217116
rect 147594 217104 147600 217116
rect 150710 217104 150716 217116
rect 147594 217076 150716 217104
rect 147594 217064 147600 217076
rect 150710 217064 150716 217076
rect 150768 217064 150774 217116
rect 520964 217064 520970 217116
rect 521022 217104 521028 217116
rect 521022 217076 524414 217104
rect 521022 217064 521028 217076
rect 524386 217036 524414 217076
rect 543200 217036 543228 217144
rect 543458 217132 543464 217144
rect 543516 217132 543522 217184
rect 524386 217008 543228 217036
rect 544396 217036 544424 217212
rect 544654 217132 544660 217184
rect 544712 217172 544718 217184
rect 564618 217172 564624 217184
rect 544712 217144 564624 217172
rect 544712 217132 544718 217144
rect 564618 217132 564624 217144
rect 564676 217132 564682 217184
rect 565998 217172 566004 217184
rect 564912 217144 566004 217172
rect 564912 217036 564940 217144
rect 565998 217132 566004 217144
rect 566056 217132 566062 217184
rect 567194 217132 567200 217184
rect 567252 217132 567258 217184
rect 569310 217132 569316 217184
rect 569368 217172 569374 217184
rect 597296 217172 597324 217416
rect 603442 217404 603448 217416
rect 603500 217404 603506 217456
rect 597462 217268 597468 217320
rect 597520 217308 597526 217320
rect 601142 217308 601148 217320
rect 597520 217280 601148 217308
rect 597520 217268 597526 217280
rect 601142 217268 601148 217280
rect 601200 217268 601206 217320
rect 601326 217268 601332 217320
rect 601384 217308 601390 217320
rect 605098 217308 605104 217320
rect 601384 217280 605104 217308
rect 601384 217268 601390 217280
rect 605098 217268 605104 217280
rect 605156 217268 605162 217320
rect 606478 217268 606484 217320
rect 606536 217308 606542 217320
rect 616138 217308 616144 217320
rect 606536 217280 616144 217308
rect 606536 217268 606542 217280
rect 616138 217268 616144 217280
rect 616196 217268 616202 217320
rect 569368 217144 597324 217172
rect 569368 217132 569374 217144
rect 598842 217132 598848 217184
rect 598900 217172 598906 217184
rect 614114 217172 614120 217184
rect 598900 217144 614120 217172
rect 598900 217132 598906 217144
rect 614114 217132 614120 217144
rect 614172 217132 614178 217184
rect 566182 217064 566188 217116
rect 566240 217104 566246 217116
rect 567010 217104 567016 217116
rect 566240 217076 567016 217104
rect 566240 217064 566246 217076
rect 567010 217064 567016 217076
rect 567068 217064 567074 217116
rect 544396 217008 564940 217036
rect 567212 217036 567240 217132
rect 567212 217008 601004 217036
rect 574278 216860 574284 216912
rect 574336 216900 574342 216912
rect 574922 216900 574928 216912
rect 574336 216872 574928 216900
rect 574336 216860 574342 216872
rect 574922 216860 574928 216872
rect 574980 216860 574986 216912
rect 590838 216860 590844 216912
rect 590896 216900 590902 216912
rect 594794 216900 594800 216912
rect 590896 216872 594800 216900
rect 590896 216860 590902 216872
rect 594794 216860 594800 216872
rect 594852 216860 594858 216912
rect 594978 216860 594984 216912
rect 595036 216900 595042 216912
rect 598842 216900 598848 216912
rect 595036 216872 598848 216900
rect 595036 216860 595042 216872
rect 598842 216860 598848 216872
rect 598900 216860 598906 216912
rect 600976 216900 601004 217008
rect 601142 216996 601148 217048
rect 601200 217036 601206 217048
rect 623314 217036 623320 217048
rect 601200 217008 623320 217036
rect 601200 216996 601206 217008
rect 623314 216996 623320 217008
rect 623372 216996 623378 217048
rect 605834 216900 605840 216912
rect 600976 216872 605840 216900
rect 605834 216860 605840 216872
rect 605892 216860 605898 216912
rect 574554 216724 574560 216776
rect 574612 216764 574618 216776
rect 575658 216764 575664 216776
rect 574612 216736 575664 216764
rect 574612 216724 574618 216736
rect 575658 216724 575664 216736
rect 575716 216724 575722 216776
rect 590838 216724 590844 216776
rect 590896 216764 590902 216776
rect 592034 216764 592040 216776
rect 590896 216736 592040 216764
rect 590896 216724 590902 216736
rect 592034 216724 592040 216736
rect 592092 216724 592098 216776
rect 595622 216724 595628 216776
rect 595680 216764 595686 216776
rect 596266 216764 596272 216776
rect 595680 216736 596272 216764
rect 595680 216724 595686 216736
rect 596266 216724 596272 216736
rect 596324 216724 596330 216776
rect 597094 216724 597100 216776
rect 597152 216764 597158 216776
rect 603994 216764 604000 216776
rect 597152 216736 604000 216764
rect 597152 216724 597158 216736
rect 603994 216724 604000 216736
rect 604052 216724 604058 216776
rect 574186 216588 574192 216640
rect 574244 216628 574250 216640
rect 576118 216628 576124 216640
rect 574244 216600 576124 216628
rect 574244 216588 574250 216600
rect 576118 216588 576124 216600
rect 576176 216588 576182 216640
rect 576854 216452 576860 216504
rect 576912 216492 576918 216504
rect 586698 216492 586704 216504
rect 576912 216464 586704 216492
rect 576912 216452 576918 216464
rect 586698 216452 586704 216464
rect 586756 216452 586762 216504
rect 595990 216384 595996 216436
rect 596048 216424 596054 216436
rect 596818 216424 596824 216436
rect 596048 216396 596824 216424
rect 596048 216384 596054 216396
rect 596818 216384 596824 216396
rect 596876 216384 596882 216436
rect 599762 215908 599768 215960
rect 599820 215948 599826 215960
rect 613378 215948 613384 215960
rect 599820 215920 613384 215948
rect 599820 215908 599826 215920
rect 613378 215908 613384 215920
rect 613436 215908 613442 215960
rect 582098 215840 582104 215892
rect 582156 215880 582162 215892
rect 595990 215880 595996 215892
rect 582156 215852 595996 215880
rect 582156 215840 582162 215852
rect 595990 215840 595996 215852
rect 596048 215840 596054 215892
rect 613838 215364 613844 215416
rect 613896 215404 613902 215416
rect 615034 215404 615040 215416
rect 613896 215376 615040 215404
rect 613896 215364 613902 215376
rect 615034 215364 615040 215376
rect 615092 215364 615098 215416
rect 636654 215296 636660 215348
rect 636712 215336 636718 215348
rect 639598 215336 639604 215348
rect 636712 215308 639604 215336
rect 636712 215296 636718 215308
rect 639598 215296 639604 215308
rect 639656 215296 639662 215348
rect 574738 215228 574744 215280
rect 574796 215268 574802 215280
rect 621658 215268 621664 215280
rect 574796 215240 621664 215268
rect 574796 215228 574802 215240
rect 621658 215228 621664 215240
rect 621716 215228 621722 215280
rect 574278 215092 574284 215144
rect 574336 215132 574342 215144
rect 619634 215132 619640 215144
rect 574336 215104 619640 215132
rect 574336 215092 574342 215104
rect 619634 215092 619640 215104
rect 619692 215092 619698 215144
rect 675846 215092 675852 215144
rect 675904 215132 675910 215144
rect 677226 215132 677232 215144
rect 675904 215104 677232 215132
rect 675904 215092 675910 215104
rect 677226 215092 677232 215104
rect 677284 215092 677290 215144
rect 577682 214956 577688 215008
rect 577740 214996 577746 215008
rect 626074 214996 626080 215008
rect 577740 214968 626080 214996
rect 577740 214956 577746 214968
rect 626074 214956 626080 214968
rect 626132 214956 626138 215008
rect 663518 214888 663524 214940
rect 663576 214928 663582 214940
rect 664438 214928 664444 214940
rect 663576 214900 664444 214928
rect 663576 214888 663582 214900
rect 664438 214888 664444 214900
rect 664496 214888 664502 214940
rect 575106 214820 575112 214872
rect 575164 214860 575170 214872
rect 622394 214860 622400 214872
rect 575164 214832 622400 214860
rect 575164 214820 575170 214832
rect 622394 214820 622400 214832
rect 622452 214820 622458 214872
rect 575658 214684 575664 214736
rect 575716 214724 575722 214736
rect 616690 214724 616696 214736
rect 575716 214696 616696 214724
rect 575716 214684 575722 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 616874 214684 616880 214736
rect 616932 214724 616938 214736
rect 617794 214724 617800 214736
rect 616932 214696 617800 214724
rect 616932 214684 616938 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 624418 214684 624424 214736
rect 624476 214724 624482 214736
rect 633802 214724 633808 214736
rect 624476 214696 633808 214724
rect 624476 214684 624482 214696
rect 633802 214684 633808 214696
rect 633860 214684 633866 214736
rect 575934 214548 575940 214600
rect 575992 214588 575998 214600
rect 575992 214560 625154 214588
rect 575992 214548 575998 214560
rect 576118 214412 576124 214464
rect 576176 214452 576182 214464
rect 620002 214452 620008 214464
rect 576176 214424 620008 214452
rect 576176 214412 576182 214424
rect 620002 214412 620008 214424
rect 620060 214412 620066 214464
rect 625126 214452 625154 214560
rect 626626 214548 626632 214600
rect 626684 214588 626690 214600
rect 627178 214588 627184 214600
rect 626684 214560 627184 214588
rect 626684 214548 626690 214560
rect 627178 214548 627184 214560
rect 627236 214548 627242 214600
rect 630766 214548 630772 214600
rect 630824 214588 630830 214600
rect 631594 214588 631600 214600
rect 630824 214560 631600 214588
rect 630824 214548 630830 214560
rect 631594 214548 631600 214560
rect 631652 214548 631658 214600
rect 662046 214548 662052 214600
rect 662104 214588 662110 214600
rect 663242 214588 663248 214600
rect 662104 214560 663248 214588
rect 662104 214548 662110 214560
rect 663242 214548 663248 214560
rect 663300 214548 663306 214600
rect 628282 214452 628288 214464
rect 625126 214424 628288 214452
rect 628282 214412 628288 214424
rect 628340 214412 628346 214464
rect 658734 214344 658740 214396
rect 658792 214384 658798 214396
rect 661678 214384 661684 214396
rect 658792 214356 661684 214384
rect 658792 214344 658798 214356
rect 661678 214344 661684 214356
rect 661736 214344 661742 214396
rect 600406 214276 600412 214328
rect 600464 214316 600470 214328
rect 600774 214316 600780 214328
rect 600464 214288 600780 214316
rect 600464 214276 600470 214288
rect 600774 214276 600780 214288
rect 600832 214276 600838 214328
rect 608686 214276 608692 214328
rect 608744 214316 608750 214328
rect 609514 214316 609520 214328
rect 608744 214288 609520 214316
rect 608744 214276 608750 214288
rect 609514 214276 609520 214288
rect 609572 214276 609578 214328
rect 616690 214276 616696 214328
rect 616748 214316 616754 214328
rect 624418 214316 624424 214328
rect 616748 214288 624424 214316
rect 616748 214276 616754 214288
rect 624418 214276 624424 214288
rect 624476 214276 624482 214328
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 40678 213976 40684 213988
rect 35860 213948 40684 213976
rect 35860 213936 35866 213948
rect 40678 213936 40684 213948
rect 40736 213936 40742 213988
rect 626442 213868 626448 213920
rect 626500 213908 626506 213920
rect 629386 213908 629392 213920
rect 626500 213880 629392 213908
rect 626500 213868 626506 213880
rect 629386 213868 629392 213880
rect 629444 213868 629450 213920
rect 638310 213868 638316 213920
rect 638368 213908 638374 213920
rect 640058 213908 640064 213920
rect 638368 213880 640064 213908
rect 638368 213868 638374 213880
rect 640058 213868 640064 213880
rect 640116 213868 640122 213920
rect 648522 213868 648528 213920
rect 648580 213908 648586 213920
rect 650638 213908 650644 213920
rect 648580 213880 650644 213908
rect 648580 213868 648586 213880
rect 650638 213868 650644 213880
rect 650696 213868 650702 213920
rect 655698 213868 655704 213920
rect 655756 213908 655762 213920
rect 656802 213908 656808 213920
rect 655756 213880 656808 213908
rect 655756 213868 655762 213880
rect 656802 213868 656808 213880
rect 656860 213868 656866 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 645486 213732 645492 213784
rect 645544 213772 645550 213784
rect 651190 213772 651196 213784
rect 645544 213744 651196 213772
rect 645544 213732 645550 213744
rect 651190 213732 651196 213744
rect 651248 213732 651254 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 662966 213772 662972 213784
rect 661000 213744 662972 213772
rect 661000 213732 661006 213744
rect 662966 213732 662972 213744
rect 663024 213732 663030 213784
rect 575290 213596 575296 213648
rect 575348 213636 575354 213648
rect 601786 213636 601792 213648
rect 575348 213608 601792 213636
rect 575348 213596 575354 213608
rect 601786 213596 601792 213608
rect 601844 213596 601850 213648
rect 652018 213596 652024 213648
rect 652076 213636 652082 213648
rect 657998 213636 658004 213648
rect 652076 213608 658004 213636
rect 652076 213596 652082 213608
rect 657998 213596 658004 213608
rect 658056 213596 658062 213648
rect 659562 213596 659568 213648
rect 659620 213636 659626 213648
rect 664622 213636 664628 213648
rect 659620 213608 664628 213636
rect 659620 213596 659626 213608
rect 664622 213596 664628 213608
rect 664680 213596 664686 213648
rect 575474 213460 575480 213512
rect 575532 213500 575538 213512
rect 601234 213500 601240 213512
rect 575532 213472 601240 213500
rect 575532 213460 575538 213472
rect 601234 213460 601240 213472
rect 601292 213460 601298 213512
rect 639966 213460 639972 213512
rect 640024 213500 640030 213512
rect 642082 213500 642088 213512
rect 640024 213472 642088 213500
rect 640024 213460 640030 213472
rect 642082 213460 642088 213472
rect 642140 213460 642146 213512
rect 650454 213460 650460 213512
rect 650512 213500 650518 213512
rect 658918 213500 658924 213512
rect 650512 213472 658924 213500
rect 650512 213460 650518 213472
rect 658918 213460 658924 213472
rect 658976 213460 658982 213512
rect 576302 213324 576308 213376
rect 576360 213364 576366 213376
rect 612826 213364 612832 213376
rect 576360 213336 612832 213364
rect 576360 213324 576366 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 641622 213324 641628 213376
rect 641680 213364 641686 213376
rect 654778 213364 654784 213376
rect 641680 213336 654784 213364
rect 641680 213324 641686 213336
rect 654778 213324 654784 213336
rect 654836 213324 654842 213376
rect 574922 213188 574928 213240
rect 574980 213228 574986 213240
rect 623866 213228 623872 213240
rect 574980 213200 623872 213228
rect 574980 213188 574986 213200
rect 623866 213188 623872 213200
rect 623924 213188 623930 213240
rect 635550 213188 635556 213240
rect 635608 213228 635614 213240
rect 651834 213228 651840 213240
rect 635608 213200 651840 213228
rect 635608 213188 635614 213200
rect 651834 213188 651840 213200
rect 651892 213188 651898 213240
rect 652846 213188 652852 213240
rect 652904 213228 652910 213240
rect 660206 213228 660212 213240
rect 652904 213200 660212 213228
rect 652904 213188 652910 213200
rect 660206 213188 660212 213200
rect 660264 213188 660270 213240
rect 675846 213188 675852 213240
rect 675904 213228 675910 213240
rect 676674 213228 676680 213240
rect 675904 213200 676680 213228
rect 675904 213188 675910 213200
rect 676674 213188 676680 213200
rect 676732 213188 676738 213240
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 632698 212848 632704 212900
rect 632756 212888 632762 212900
rect 634354 212888 634360 212900
rect 632756 212860 634360 212888
rect 632756 212848 632762 212860
rect 634354 212848 634360 212860
rect 634412 212848 634418 212900
rect 628650 212712 628656 212764
rect 628708 212752 628714 212764
rect 632698 212752 632704 212764
rect 628708 212724 632704 212752
rect 628708 212712 628714 212724
rect 632698 212712 632704 212724
rect 632756 212712 632762 212764
rect 637206 212712 637212 212764
rect 637264 212752 637270 212764
rect 641438 212752 641444 212764
rect 637264 212724 641444 212752
rect 637264 212712 637270 212724
rect 641438 212712 641444 212724
rect 641496 212712 641502 212764
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 41690 211188 41696 211200
rect 35860 211160 41696 211188
rect 35860 211148 35866 211160
rect 41690 211148 41696 211160
rect 41748 211148 41754 211200
rect 610066 210264 610072 210316
rect 610124 210304 610130 210316
rect 610618 210304 610624 210316
rect 610124 210276 610624 210304
rect 610124 210264 610130 210276
rect 610618 210264 610624 210276
rect 610676 210264 610682 210316
rect 578786 209856 578792 209908
rect 578844 209896 578850 209908
rect 580994 209896 581000 209908
rect 578844 209868 581000 209896
rect 578844 209856 578850 209868
rect 580994 209856 581000 209868
rect 581052 209856 581058 209908
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 591298 208632 591304 208684
rect 591356 208672 591362 208684
rect 625126 208672 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 652260 209528 654134 209556
rect 652260 209516 652266 209528
rect 654106 209080 654134 209528
rect 667014 209080 667020 209092
rect 654106 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 591356 208644 625154 208672
rect 591356 208632 591362 208644
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 40034 208400 40040 208412
rect 35860 208372 40040 208400
rect 35860 208360 35866 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578602 208292 578608 208344
rect 578660 208332 578666 208344
rect 589458 208332 589464 208344
rect 578660 208304 589464 208332
rect 578660 208292 578666 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 579614 207612 579620 207664
rect 579672 207652 579678 207664
rect 589458 207652 589464 207664
rect 579672 207624 589464 207652
rect 579672 207612 579678 207624
rect 589458 207612 589464 207624
rect 589516 207612 589522 207664
rect 580994 206252 581000 206304
rect 581052 206292 581058 206304
rect 589642 206292 589648 206304
rect 581052 206264 589648 206292
rect 581052 206252 581058 206264
rect 589642 206252 589648 206264
rect 589700 206252 589706 206304
rect 578234 205776 578240 205828
rect 578292 205816 578298 205828
rect 580994 205816 581000 205828
rect 578292 205788 581000 205816
rect 578292 205776 578298 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 669314 199044 669320 199096
rect 669372 199084 669378 199096
rect 670786 199084 670792 199096
rect 669372 199056 670792 199084
rect 669372 199044 669378 199056
rect 670786 199044 670792 199056
rect 670844 199044 670850 199096
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 45462 196596 45468 196648
rect 45520 196636 45526 196648
rect 48774 196636 48780 196648
rect 45520 196608 48780 196636
rect 45520 196596 45526 196608
rect 48774 196596 48780 196608
rect 48832 196596 48838 196648
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 669406 194148 669412 194200
rect 669464 194188 669470 194200
rect 670786 194188 670792 194200
rect 669464 194160 670792 194188
rect 669464 194148 669470 194160
rect 670786 194148 670792 194160
rect 670844 194148 670850 194200
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 667934 189252 667940 189304
rect 667992 189292 667998 189304
rect 670786 189292 670792 189304
rect 667992 189264 670792 189292
rect 667992 189252 667998 189264
rect 670786 189252 670792 189264
rect 670844 189252 670850 189304
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 583018 175244 583024 175296
rect 583076 175284 583082 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 583076 175256 586514 175284
rect 583076 175244 583082 175256
rect 667934 174564 667940 174616
rect 667992 174604 667998 174616
rect 669774 174604 669780 174616
rect 667992 174576 669780 174604
rect 667992 174564 667998 174576
rect 669774 174564 669780 174576
rect 669832 174564 669838 174616
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 581638 171096 581644 171148
rect 581696 171136 581702 171148
rect 589458 171136 589464 171148
rect 581696 171108 589464 171136
rect 581696 171096 581702 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 579522 170960 579528 171012
rect 579580 171000 579586 171012
rect 583018 171000 583024 171012
rect 579580 170972 583024 171000
rect 579580 170960 579586 170972
rect 583018 170960 583024 170972
rect 583076 170960 583082 171012
rect 582374 169736 582380 169788
rect 582432 169776 582438 169788
rect 589458 169776 589464 169788
rect 582432 169748 589464 169776
rect 582432 169736 582438 169748
rect 589458 169736 589464 169748
rect 589516 169736 589522 169788
rect 578326 169668 578332 169720
rect 578384 169708 578390 169720
rect 580902 169708 580908 169720
rect 578384 169680 580908 169708
rect 578384 169668 578390 169680
rect 580902 169668 580908 169680
rect 580960 169668 580966 169720
rect 668026 169668 668032 169720
rect 668084 169708 668090 169720
rect 670326 169708 670332 169720
rect 668084 169680 670332 169708
rect 668084 169668 668090 169680
rect 670326 169668 670332 169680
rect 670384 169668 670390 169720
rect 579614 168376 579620 168428
rect 579672 168416 579678 168428
rect 589458 168416 589464 168428
rect 579672 168388 589464 168416
rect 579672 168376 579678 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578970 167152 578976 167204
rect 579028 167192 579034 167204
rect 581638 167192 581644 167204
rect 579028 167164 581644 167192
rect 579028 167152 579034 167164
rect 581638 167152 581644 167164
rect 581696 167152 581702 167204
rect 581638 167016 581644 167068
rect 581696 167056 581702 167068
rect 589458 167056 589464 167068
rect 581696 167028 589464 167056
rect 581696 167016 581702 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 578878 165520 578884 165572
rect 578936 165560 578942 165572
rect 582374 165560 582380 165572
rect 578936 165532 582380 165560
rect 578936 165520 578942 165532
rect 582374 165520 582380 165532
rect 582432 165520 582438 165572
rect 667934 164772 667940 164824
rect 667992 164812 667998 164824
rect 670142 164812 670148 164824
rect 667992 164784 670148 164812
rect 667992 164772 667998 164784
rect 670142 164772 670148 164784
rect 670200 164772 670206 164824
rect 585962 164228 585968 164280
rect 586020 164268 586026 164280
rect 589458 164268 589464 164280
rect 586020 164240 589464 164268
rect 586020 164228 586026 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 584398 162868 584404 162920
rect 584456 162908 584462 162920
rect 589458 162908 589464 162920
rect 584456 162880 589464 162908
rect 584456 162868 584462 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 676122 162800 676128 162852
rect 676180 162840 676186 162852
rect 678238 162840 678244 162852
rect 676180 162812 678244 162840
rect 676180 162800 676186 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 675938 162596 675944 162648
rect 675996 162636 676002 162648
rect 679618 162636 679624 162648
rect 675996 162608 679624 162636
rect 675996 162596 676002 162608
rect 679618 162596 679624 162608
rect 679676 162596 679682 162648
rect 675846 161712 675852 161764
rect 675904 161752 675910 161764
rect 680998 161752 681004 161764
rect 675904 161724 681004 161752
rect 675904 161712 675910 161724
rect 680998 161712 681004 161724
rect 681056 161712 681062 161764
rect 580258 161440 580264 161492
rect 580316 161480 580322 161492
rect 589458 161480 589464 161492
rect 580316 161452 589464 161480
rect 580316 161440 580322 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 582374 160080 582380 160132
rect 582432 160120 582438 160132
rect 589458 160120 589464 160132
rect 582432 160092 589464 160120
rect 582432 160080 582438 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 579246 160012 579252 160064
rect 579304 160052 579310 160064
rect 581638 160052 581644 160064
rect 579304 160024 581644 160052
rect 579304 160012 579310 160024
rect 581638 160012 581644 160024
rect 581696 160012 581702 160064
rect 581822 158788 581828 158840
rect 581880 158828 581886 158840
rect 589458 158828 589464 158840
rect 581880 158800 589464 158828
rect 581880 158788 581886 158800
rect 589458 158788 589464 158800
rect 589516 158788 589522 158840
rect 579154 158652 579160 158704
rect 579212 158692 579218 158704
rect 585962 158692 585968 158704
rect 579212 158664 585968 158692
rect 579212 158652 579218 158664
rect 585962 158652 585968 158664
rect 586020 158652 586026 158704
rect 585778 157360 585784 157412
rect 585836 157400 585842 157412
rect 589458 157400 589464 157412
rect 585836 157372 589464 157400
rect 585836 157360 585842 157372
rect 589458 157360 589464 157372
rect 589516 157360 589522 157412
rect 579522 155864 579528 155916
rect 579580 155904 579586 155916
rect 584398 155904 584404 155916
rect 579580 155876 584404 155904
rect 579580 155864 579586 155876
rect 584398 155864 584404 155876
rect 584456 155864 584462 155916
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 578234 154504 578240 154556
rect 578292 154544 578298 154556
rect 580258 154544 580264 154556
rect 578292 154516 580264 154544
rect 578292 154504 578298 154516
rect 580258 154504 580264 154516
rect 580316 154504 580322 154556
rect 580442 153212 580448 153264
rect 580500 153252 580506 153264
rect 589458 153252 589464 153264
rect 580500 153224 589464 153252
rect 580500 153212 580506 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 582374 152776 582380 152788
rect 578292 152748 582380 152776
rect 578292 152736 578298 152748
rect 582374 152736 582380 152748
rect 582432 152736 582438 152788
rect 583018 151784 583024 151836
rect 583076 151824 583082 151836
rect 589458 151824 589464 151836
rect 583076 151796 589464 151824
rect 583076 151784 583082 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 581822 150600 581828 150612
rect 578936 150572 581828 150600
rect 578936 150560 578942 150572
rect 581822 150560 581828 150572
rect 581880 150560 581886 150612
rect 581638 150424 581644 150476
rect 581696 150464 581702 150476
rect 589458 150464 589464 150476
rect 581696 150436 589464 150464
rect 581696 150424 581702 150436
rect 589458 150424 589464 150436
rect 589516 150424 589522 150476
rect 579522 147364 579528 147416
rect 579580 147404 579586 147416
rect 585778 147404 585784 147416
rect 579580 147376 585784 147404
rect 579580 147364 579586 147376
rect 585778 147364 585784 147376
rect 585836 147364 585842 147416
rect 587342 146276 587348 146328
rect 587400 146316 587406 146328
rect 589366 146316 589372 146328
rect 587400 146288 589372 146316
rect 587400 146276 587406 146288
rect 589366 146276 589372 146288
rect 589424 146276 589430 146328
rect 668486 146004 668492 146056
rect 668544 146044 668550 146056
rect 670786 146044 670792 146056
rect 668544 146016 670792 146044
rect 668544 146004 668550 146016
rect 670786 146004 670792 146016
rect 670844 146004 670850 146056
rect 578878 145528 578884 145580
rect 578936 145568 578942 145580
rect 589182 145568 589188 145580
rect 578936 145540 589188 145568
rect 578936 145528 578942 145540
rect 589182 145528 589188 145540
rect 589240 145528 589246 145580
rect 585778 144916 585784 144968
rect 585836 144956 585842 144968
rect 589458 144956 589464 144968
rect 585836 144928 589464 144956
rect 585836 144916 585842 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 578602 143148 578608 143200
rect 578660 143188 578666 143200
rect 580442 143188 580448 143200
rect 578660 143160 580448 143188
rect 578660 143148 578666 143160
rect 580442 143148 580448 143160
rect 580500 143148 580506 143200
rect 580258 142128 580264 142180
rect 580316 142168 580322 142180
rect 589458 142168 589464 142180
rect 580316 142140 589464 142168
rect 580316 142128 580322 142140
rect 589458 142128 589464 142140
rect 589516 142128 589522 142180
rect 579522 140564 579528 140616
rect 579580 140604 579586 140616
rect 583018 140604 583024 140616
rect 579580 140576 583024 140604
rect 579580 140564 579586 140576
rect 583018 140564 583024 140576
rect 583076 140564 583082 140616
rect 584398 139408 584404 139460
rect 584456 139448 584462 139460
rect 589458 139448 589464 139460
rect 584456 139420 589464 139448
rect 584456 139408 584462 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578694 139340 578700 139392
rect 578752 139380 578758 139392
rect 581638 139380 581644 139392
rect 578752 139352 581644 139380
rect 578752 139340 578758 139352
rect 581638 139340 581644 139352
rect 581696 139340 581702 139392
rect 581638 136620 581644 136672
rect 581696 136660 581702 136672
rect 589458 136660 589464 136672
rect 581696 136632 589464 136660
rect 581696 136620 581702 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 668026 136280 668032 136332
rect 668084 136320 668090 136332
rect 669958 136320 669964 136332
rect 668084 136292 669964 136320
rect 668084 136280 668090 136292
rect 669958 136280 669964 136292
rect 670016 136280 670022 136332
rect 578326 135872 578332 135924
rect 578384 135912 578390 135924
rect 587342 135912 587348 135924
rect 578384 135884 587348 135912
rect 578384 135872 578390 135884
rect 587342 135872 587348 135884
rect 587400 135872 587406 135924
rect 587158 135260 587164 135312
rect 587216 135300 587222 135312
rect 589274 135300 589280 135312
rect 587216 135272 589280 135300
rect 587216 135260 587222 135272
rect 589274 135260 589280 135272
rect 589332 135260 589338 135312
rect 578234 134240 578240 134292
rect 578292 134280 578298 134292
rect 585778 134280 585784 134292
rect 578292 134252 585784 134280
rect 578292 134240 578298 134252
rect 585778 134240 585784 134252
rect 585836 134240 585842 134292
rect 585962 133900 585968 133952
rect 586020 133940 586026 133952
rect 589458 133940 589464 133952
rect 586020 133912 589464 133940
rect 586020 133900 586026 133912
rect 589458 133900 589464 133912
rect 589516 133900 589522 133952
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 579246 133152 579252 133204
rect 579304 133192 579310 133204
rect 589090 133192 589096 133204
rect 579304 133164 589096 133192
rect 579304 133152 579310 133164
rect 589090 133152 589096 133164
rect 589148 133152 589154 133204
rect 582374 131724 582380 131776
rect 582432 131764 582438 131776
rect 589918 131764 589924 131776
rect 582432 131736 589924 131764
rect 582432 131724 582438 131736
rect 589918 131724 589924 131736
rect 589976 131724 589982 131776
rect 579522 129684 579528 129736
rect 579580 129724 579586 129736
rect 582374 129724 582380 129736
rect 579580 129696 582380 129724
rect 579580 129684 579586 129696
rect 582374 129684 582380 129696
rect 582432 129684 582438 129736
rect 583018 128324 583024 128376
rect 583076 128364 583082 128376
rect 589458 128364 589464 128376
rect 583076 128336 589464 128364
rect 583076 128324 583082 128336
rect 589458 128324 589464 128336
rect 589516 128324 589522 128376
rect 578326 128256 578332 128308
rect 578384 128296 578390 128308
rect 580258 128296 580264 128308
rect 578384 128268 580264 128296
rect 578384 128256 578390 128268
rect 580258 128256 580264 128268
rect 580316 128256 580322 128308
rect 580442 126964 580448 127016
rect 580500 127004 580506 127016
rect 589458 127004 589464 127016
rect 580500 126976 589464 127004
rect 580500 126964 580506 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 668210 125128 668216 125180
rect 668268 125168 668274 125180
rect 669774 125168 669780 125180
rect 668268 125140 669780 125168
rect 668268 125128 668274 125140
rect 669774 125128 669780 125140
rect 669832 125128 669838 125180
rect 585778 124176 585784 124228
rect 585836 124216 585842 124228
rect 589458 124216 589464 124228
rect 585836 124188 589464 124216
rect 585836 124176 585842 124188
rect 589458 124176 589464 124188
rect 589516 124176 589522 124228
rect 579246 124108 579252 124160
rect 579304 124148 579310 124160
rect 584398 124148 584404 124160
rect 579304 124120 584404 124148
rect 579304 124108 579310 124120
rect 584398 124108 584404 124120
rect 584456 124108 584462 124160
rect 579246 122816 579252 122868
rect 579304 122856 579310 122868
rect 589458 122856 589464 122868
rect 579304 122828 589464 122856
rect 579304 122816 579310 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 584398 121456 584404 121508
rect 584456 121496 584462 121508
rect 589458 121496 589464 121508
rect 584456 121468 589464 121496
rect 584456 121456 584462 121468
rect 589458 121456 589464 121468
rect 589516 121456 589522 121508
rect 579062 121116 579068 121168
rect 579120 121156 579126 121168
rect 581638 121156 581644 121168
rect 579120 121128 581644 121156
rect 579120 121116 579126 121128
rect 581638 121116 581644 121128
rect 581696 121116 581702 121168
rect 582006 120708 582012 120760
rect 582064 120748 582070 120760
rect 590102 120748 590108 120760
rect 582064 120720 590108 120748
rect 582064 120708 582070 120720
rect 590102 120708 590108 120720
rect 590160 120708 590166 120760
rect 578510 118600 578516 118652
rect 578568 118640 578574 118652
rect 587158 118640 587164 118652
rect 578568 118612 587164 118640
rect 578568 118600 578574 118612
rect 587158 118600 587164 118612
rect 587216 118600 587222 118652
rect 668026 117648 668032 117700
rect 668084 117688 668090 117700
rect 670326 117688 670332 117700
rect 668084 117660 670332 117688
rect 668084 117648 668090 117660
rect 670326 117648 670332 117660
rect 670384 117648 670390 117700
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 682378 117280 682384 117292
rect 675904 117252 682384 117280
rect 675904 117240 675910 117252
rect 682378 117240 682384 117252
rect 682436 117240 682442 117292
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 585962 116940 585968 116952
rect 579580 116912 585968 116940
rect 579580 116900 579586 116912
rect 585962 116900 585968 116912
rect 586020 116900 586026 116952
rect 587802 115948 587808 116000
rect 587860 115988 587866 116000
rect 589458 115988 589464 116000
rect 587860 115960 589464 115988
rect 587860 115948 587866 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 585134 115336 585140 115388
rect 585192 115376 585198 115388
rect 590286 115376 590292 115388
rect 585192 115348 590292 115376
rect 585192 115336 585198 115348
rect 590286 115336 590292 115348
rect 590344 115336 590350 115388
rect 579062 115200 579068 115252
rect 579120 115240 579126 115252
rect 587802 115240 587808 115252
rect 579120 115212 587808 115240
rect 579120 115200 579126 115212
rect 587802 115200 587808 115212
rect 587860 115200 587866 115252
rect 587158 114520 587164 114572
rect 587216 114560 587222 114572
rect 589642 114560 589648 114572
rect 587216 114532 589648 114560
rect 587216 114520 587222 114532
rect 589642 114520 589648 114532
rect 589700 114520 589706 114572
rect 579522 114384 579528 114436
rect 579580 114424 579586 114436
rect 591298 114424 591304 114436
rect 579580 114396 591304 114424
rect 579580 114384 579586 114396
rect 591298 114384 591304 114396
rect 591356 114384 591362 114436
rect 668210 114248 668216 114300
rect 668268 114288 668274 114300
rect 669590 114288 669596 114300
rect 668268 114260 669596 114288
rect 668268 114248 668274 114260
rect 669590 114248 669596 114260
rect 669648 114248 669654 114300
rect 579522 113092 579528 113144
rect 579580 113132 579586 113144
rect 588538 113132 588544 113144
rect 579580 113104 588544 113132
rect 579580 113092 579586 113104
rect 588538 113092 588544 113104
rect 588596 113092 588602 113144
rect 588538 110440 588544 110492
rect 588596 110480 588602 110492
rect 589642 110480 589648 110492
rect 588596 110452 589648 110480
rect 588596 110440 588602 110452
rect 589642 110440 589648 110452
rect 589700 110440 589706 110492
rect 579430 110236 579436 110288
rect 579488 110276 579494 110288
rect 582006 110276 582012 110288
rect 579488 110248 582012 110276
rect 579488 110236 579494 110248
rect 582006 110236 582012 110248
rect 582064 110236 582070 110288
rect 581822 109692 581828 109744
rect 581880 109732 581886 109744
rect 589458 109732 589464 109744
rect 581880 109704 589464 109732
rect 581880 109692 581886 109704
rect 589458 109692 589464 109704
rect 589516 109692 589522 109744
rect 578326 108332 578332 108384
rect 578384 108372 578390 108384
rect 585134 108372 585140 108384
rect 578384 108344 585140 108372
rect 578384 108332 578390 108344
rect 585134 108332 585140 108344
rect 585192 108332 585198 108384
rect 589458 107692 589464 107704
rect 579632 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 579632 107624 579660 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 579660 107624
rect 578936 107584 578942 107596
rect 580258 106904 580264 106956
rect 580316 106944 580322 106956
rect 589274 106944 589280 106956
rect 580316 106916 589280 106944
rect 580316 106904 580322 106916
rect 589274 106904 589280 106916
rect 589332 106904 589338 106956
rect 578326 106496 578332 106548
rect 578384 106536 578390 106548
rect 580442 106536 580448 106548
rect 578384 106508 580448 106536
rect 578384 106496 578390 106508
rect 580442 106496 580448 106508
rect 580500 106496 580506 106548
rect 580626 106292 580632 106344
rect 580684 106332 580690 106344
rect 589458 106332 589464 106344
rect 580684 106304 589464 106332
rect 580684 106292 580690 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 667198 106156 667204 106208
rect 667256 106196 667262 106208
rect 670694 106196 670700 106208
rect 667256 106168 670700 106196
rect 667256 106156 667262 106168
rect 670694 106156 670700 106168
rect 670752 106156 670758 106208
rect 581638 104864 581644 104916
rect 581696 104904 581702 104916
rect 589458 104904 589464 104916
rect 581696 104876 589464 104904
rect 581696 104864 581702 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 579522 103300 579528 103352
rect 579580 103340 579586 103352
rect 583018 103340 583024 103352
rect 579580 103312 583024 103340
rect 579580 103300 579586 103312
rect 583018 103300 583024 103312
rect 583076 103300 583082 103352
rect 582374 102756 582380 102808
rect 582432 102796 582438 102808
rect 589918 102796 589924 102808
rect 582432 102768 589924 102796
rect 582432 102756 582438 102768
rect 589918 102756 589924 102768
rect 589976 102756 589982 102808
rect 585962 100716 585968 100768
rect 586020 100756 586026 100768
rect 589458 100756 589464 100768
rect 586020 100728 589464 100756
rect 586020 100716 586026 100728
rect 589458 100716 589464 100728
rect 589516 100716 589522 100768
rect 615218 100104 615224 100156
rect 615276 100144 615282 100156
rect 668026 100144 668032 100156
rect 615276 100116 668032 100144
rect 615276 100104 615282 100116
rect 668026 100104 668032 100116
rect 668084 100104 668090 100156
rect 613378 99968 613384 100020
rect 613436 100008 613442 100020
rect 668486 100008 668492 100020
rect 613436 99980 668492 100008
rect 613436 99968 613442 99980
rect 668486 99968 668492 99980
rect 668544 99968 668550 100020
rect 577498 99288 577504 99340
rect 577556 99328 577562 99340
rect 595254 99328 595260 99340
rect 577556 99300 595260 99328
rect 577556 99288 577562 99300
rect 595254 99288 595260 99300
rect 595312 99288 595318 99340
rect 624602 99288 624608 99340
rect 624660 99328 624666 99340
rect 632974 99328 632980 99340
rect 624660 99300 632980 99328
rect 624660 99288 624666 99300
rect 632974 99288 632980 99300
rect 633032 99288 633038 99340
rect 579522 99152 579528 99204
rect 579580 99192 579586 99204
rect 585778 99192 585784 99204
rect 579580 99164 585784 99192
rect 579580 99152 579586 99164
rect 585778 99152 585784 99164
rect 585836 99152 585842 99204
rect 626810 99152 626816 99204
rect 626868 99192 626874 99204
rect 636378 99192 636384 99204
rect 626868 99164 636384 99192
rect 626868 99152 626874 99164
rect 636378 99152 636384 99164
rect 636436 99152 636442 99204
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 634078 99056 634084 99068
rect 625120 99028 634084 99056
rect 625120 99016 625126 99028
rect 634078 99016 634084 99028
rect 634136 99016 634142 99068
rect 629754 98880 629760 98932
rect 629812 98920 629818 98932
rect 640978 98920 640984 98932
rect 629812 98892 640984 98920
rect 629812 98880 629818 98892
rect 640978 98880 640984 98892
rect 641036 98880 641042 98932
rect 622302 98744 622308 98796
rect 622360 98784 622366 98796
rect 629478 98784 629484 98796
rect 622360 98756 629484 98784
rect 622360 98744 622366 98756
rect 629478 98744 629484 98756
rect 629536 98744 629542 98796
rect 630490 98744 630496 98796
rect 630548 98784 630554 98796
rect 642542 98784 642548 98796
rect 630548 98756 642548 98784
rect 630548 98744 630554 98756
rect 642542 98744 642548 98756
rect 642600 98744 642606 98796
rect 623682 98608 623688 98660
rect 623740 98648 623746 98660
rect 632146 98648 632152 98660
rect 623740 98620 632152 98648
rect 623740 98608 623746 98620
rect 632146 98608 632152 98620
rect 632204 98608 632210 98660
rect 637850 98608 637856 98660
rect 637908 98648 637914 98660
rect 660390 98648 660396 98660
rect 637908 98620 660396 98648
rect 637908 98608 637914 98620
rect 660390 98608 660396 98620
rect 660448 98608 660454 98660
rect 605466 97928 605472 97980
rect 605524 97968 605530 97980
rect 606478 97968 606484 97980
rect 605524 97940 606484 97968
rect 605524 97928 605530 97940
rect 606478 97928 606484 97940
rect 606536 97928 606542 97980
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625614 97968 625620 97980
rect 618772 97940 625620 97968
rect 618772 97928 618778 97940
rect 625614 97928 625620 97940
rect 625672 97928 625678 97980
rect 629018 97928 629024 97980
rect 629076 97968 629082 97980
rect 639874 97968 639880 97980
rect 629076 97940 639880 97968
rect 629076 97928 629082 97940
rect 639874 97928 639880 97940
rect 639932 97928 639938 97980
rect 643002 97928 643008 97980
rect 643060 97968 643066 97980
rect 643060 97940 657952 97968
rect 643060 97928 643066 97940
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 643278 97832 643284 97844
rect 632756 97804 643284 97832
rect 632756 97792 632762 97804
rect 643278 97792 643284 97804
rect 643336 97792 643342 97844
rect 657538 97832 657544 97844
rect 655256 97804 657544 97832
rect 623130 97656 623136 97708
rect 623188 97696 623194 97708
rect 630858 97696 630864 97708
rect 623188 97668 630864 97696
rect 623188 97656 623194 97668
rect 630858 97656 630864 97668
rect 630916 97656 630922 97708
rect 633342 97656 633348 97708
rect 633400 97696 633406 97708
rect 643462 97696 643468 97708
rect 633400 97668 643468 97696
rect 633400 97656 633406 97668
rect 643462 97656 643468 97668
rect 643520 97656 643526 97708
rect 647142 97656 647148 97708
rect 647200 97696 647206 97708
rect 655256 97696 655284 97804
rect 657538 97792 657544 97804
rect 657596 97792 657602 97844
rect 657924 97832 657952 97940
rect 658182 97928 658188 97980
rect 658240 97968 658246 97980
rect 663058 97968 663064 97980
rect 658240 97940 663064 97968
rect 658240 97928 658246 97940
rect 663058 97928 663064 97940
rect 663116 97928 663122 97980
rect 659746 97832 659752 97844
rect 657924 97804 659752 97832
rect 659746 97792 659752 97804
rect 659804 97792 659810 97844
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665174 97832 665180 97844
rect 659988 97804 665180 97832
rect 659988 97792 659994 97804
rect 665174 97792 665180 97804
rect 665232 97792 665238 97844
rect 647200 97668 655284 97696
rect 647200 97656 647206 97668
rect 655422 97656 655428 97708
rect 655480 97696 655486 97708
rect 655480 97668 659056 97696
rect 655480 97656 655486 97668
rect 615034 97520 615040 97572
rect 615092 97560 615098 97572
rect 616138 97560 616144 97572
rect 615092 97532 616144 97560
rect 615092 97520 615098 97532
rect 616138 97520 616144 97532
rect 616196 97520 616202 97572
rect 621658 97520 621664 97572
rect 621716 97560 621722 97572
rect 628374 97560 628380 97572
rect 621716 97532 628380 97560
rect 621716 97520 621722 97532
rect 628374 97520 628380 97532
rect 628432 97520 628438 97572
rect 631870 97520 631876 97572
rect 631928 97560 631934 97572
rect 644934 97560 644940 97572
rect 631928 97532 644940 97560
rect 631928 97520 631934 97532
rect 644934 97520 644940 97532
rect 644992 97520 644998 97572
rect 658826 97560 658832 97572
rect 654474 97532 658832 97560
rect 579522 97452 579528 97504
rect 579580 97492 579586 97504
rect 584398 97492 584404 97504
rect 579580 97464 584404 97492
rect 579580 97452 579586 97464
rect 584398 97452 584404 97464
rect 584456 97452 584462 97504
rect 627546 97384 627552 97436
rect 627604 97424 627610 97436
rect 637574 97424 637580 97436
rect 627604 97396 637580 97424
rect 627604 97384 627610 97396
rect 637574 97384 637580 97396
rect 637632 97384 637638 97436
rect 644290 97384 644296 97436
rect 644348 97424 644354 97436
rect 654474 97424 654502 97532
rect 658826 97520 658832 97532
rect 658884 97520 658890 97572
rect 659028 97560 659056 97668
rect 659194 97656 659200 97708
rect 659252 97696 659258 97708
rect 663886 97696 663892 97708
rect 659252 97668 663892 97696
rect 659252 97656 659258 97668
rect 663886 97656 663892 97668
rect 663944 97656 663950 97708
rect 662506 97560 662512 97572
rect 659028 97532 662512 97560
rect 662506 97520 662512 97532
rect 662564 97520 662570 97572
rect 644348 97396 654502 97424
rect 644348 97384 644354 97396
rect 654594 97384 654600 97436
rect 654652 97424 654658 97436
rect 659562 97424 659568 97436
rect 654652 97396 659568 97424
rect 654652 97384 654658 97396
rect 659562 97384 659568 97396
rect 659620 97384 659626 97436
rect 612642 97248 612648 97300
rect 612700 97288 612706 97300
rect 620278 97288 620284 97300
rect 612700 97260 620284 97288
rect 612700 97248 612706 97260
rect 620278 97248 620284 97260
rect 620336 97248 620342 97300
rect 628190 97248 628196 97300
rect 628248 97288 628254 97300
rect 639046 97288 639052 97300
rect 628248 97260 639052 97288
rect 628248 97248 628254 97260
rect 639046 97248 639052 97260
rect 639104 97248 639110 97300
rect 643738 97248 643744 97300
rect 643796 97288 643802 97300
rect 650822 97288 650828 97300
rect 643796 97260 650828 97288
rect 643796 97248 643802 97260
rect 650822 97248 650828 97260
rect 650880 97248 650886 97300
rect 651098 97248 651104 97300
rect 651156 97288 651162 97300
rect 655054 97288 655060 97300
rect 651156 97260 655060 97288
rect 651156 97248 651162 97260
rect 655054 97248 655060 97260
rect 655112 97248 655118 97300
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 620094 97112 620100 97164
rect 620152 97152 620158 97164
rect 626258 97152 626264 97164
rect 620152 97124 626264 97152
rect 620152 97112 620158 97124
rect 626258 97112 626264 97124
rect 626316 97112 626322 97164
rect 634262 97112 634268 97164
rect 634320 97152 634326 97164
rect 644750 97152 644756 97164
rect 634320 97124 644756 97152
rect 634320 97112 634326 97124
rect 644750 97112 644756 97124
rect 644808 97112 644814 97164
rect 650362 97112 650368 97164
rect 650420 97152 650426 97164
rect 658274 97152 658280 97164
rect 650420 97124 658280 97152
rect 650420 97112 650426 97124
rect 658274 97112 658280 97124
rect 658332 97112 658338 97164
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 643738 97016 643744 97028
rect 634780 96988 643744 97016
rect 634780 96976 634786 96988
rect 643738 96976 643744 96988
rect 643796 96976 643802 97028
rect 651834 96976 651840 97028
rect 651892 97016 651898 97028
rect 654594 97016 654600 97028
rect 651892 96988 654600 97016
rect 651892 96976 651898 96988
rect 654594 96976 654600 96988
rect 654652 96976 654658 97028
rect 597646 96908 597652 96960
rect 597704 96948 597710 96960
rect 598198 96948 598204 96960
rect 597704 96920 598204 96948
rect 597704 96908 597710 96920
rect 598198 96908 598204 96920
rect 598256 96908 598262 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 618898 96948 618904 96960
rect 615828 96920 618904 96948
rect 615828 96908 615834 96920
rect 618898 96908 618904 96920
rect 618956 96908 618962 96960
rect 645210 96908 645216 96960
rect 645268 96948 645274 96960
rect 649258 96948 649264 96960
rect 645268 96920 649264 96948
rect 645268 96908 645274 96920
rect 649258 96908 649264 96920
rect 649316 96908 649322 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 660666 96908 660672 96960
rect 660724 96948 660730 96960
rect 663426 96948 663432 96960
rect 660724 96920 663432 96948
rect 660724 96908 660730 96920
rect 663426 96908 663432 96920
rect 663484 96908 663490 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 626074 96840 626080 96892
rect 626132 96880 626138 96892
rect 635274 96880 635280 96892
rect 626132 96852 635280 96880
rect 626132 96840 626138 96852
rect 635274 96840 635280 96852
rect 635332 96840 635338 96892
rect 653950 96772 653956 96824
rect 654008 96812 654014 96824
rect 655238 96812 655244 96824
rect 654008 96784 655244 96812
rect 654008 96772 654014 96784
rect 655238 96772 655244 96784
rect 655296 96772 655302 96824
rect 657538 96772 657544 96824
rect 657596 96812 657602 96824
rect 661954 96812 661960 96824
rect 657596 96784 661960 96812
rect 657596 96772 657602 96784
rect 661954 96772 661960 96784
rect 662012 96772 662018 96824
rect 606202 96704 606208 96756
rect 606260 96744 606266 96756
rect 611998 96744 612004 96756
rect 606260 96716 612004 96744
rect 606260 96704 606266 96716
rect 611998 96704 612004 96716
rect 612056 96704 612062 96756
rect 617242 96704 617248 96756
rect 617300 96744 617306 96756
rect 618162 96744 618168 96756
rect 617300 96716 618168 96744
rect 617300 96704 617306 96716
rect 618162 96704 618168 96716
rect 618220 96704 618226 96756
rect 646682 96704 646688 96756
rect 646740 96744 646746 96756
rect 647878 96744 647884 96756
rect 646740 96716 647884 96744
rect 646740 96704 646746 96716
rect 647878 96704 647884 96716
rect 647936 96704 647942 96756
rect 631226 96568 631232 96620
rect 631284 96608 631290 96620
rect 643186 96608 643192 96620
rect 631284 96580 643192 96608
rect 631284 96568 631290 96580
rect 643186 96568 643192 96580
rect 643244 96568 643250 96620
rect 644474 96608 644480 96620
rect 643388 96580 644480 96608
rect 642266 96432 642272 96484
rect 642324 96472 642330 96484
rect 643388 96472 643416 96580
rect 644474 96568 644480 96580
rect 644532 96568 644538 96620
rect 649626 96568 649632 96620
rect 649684 96608 649690 96620
rect 650638 96608 650644 96620
rect 649684 96580 650644 96608
rect 649684 96568 649690 96580
rect 650638 96568 650644 96580
rect 650696 96568 650702 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 665358 96608 665364 96620
rect 652628 96580 665364 96608
rect 652628 96568 652634 96580
rect 665358 96568 665364 96580
rect 665416 96568 665422 96620
rect 647694 96472 647700 96484
rect 642324 96444 643416 96472
rect 643480 96444 647700 96472
rect 642324 96432 642330 96444
rect 609146 96296 609152 96348
rect 609204 96336 609210 96348
rect 621658 96336 621664 96348
rect 609204 96308 621664 96336
rect 609204 96296 609210 96308
rect 621658 96296 621664 96308
rect 621716 96296 621722 96348
rect 640058 96296 640064 96348
rect 640116 96336 640122 96348
rect 643480 96336 643508 96444
rect 647694 96432 647700 96444
rect 647752 96432 647758 96484
rect 648154 96432 648160 96484
rect 648212 96472 648218 96484
rect 652018 96472 652024 96484
rect 648212 96444 652024 96472
rect 648212 96432 648218 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 653858 96472 653864 96484
rect 652220 96444 653864 96472
rect 640116 96308 643508 96336
rect 640116 96296 640122 96308
rect 643922 96296 643928 96348
rect 643980 96336 643986 96348
rect 652220 96336 652248 96444
rect 653858 96432 653864 96444
rect 653916 96432 653922 96484
rect 643980 96308 652248 96336
rect 643980 96296 643986 96308
rect 653306 96296 653312 96348
rect 653364 96336 653370 96348
rect 664162 96336 664168 96348
rect 653364 96308 664168 96336
rect 653364 96296 653370 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 610618 96160 610624 96212
rect 610676 96200 610682 96212
rect 623038 96200 623044 96212
rect 610676 96172 623044 96200
rect 610676 96160 610682 96172
rect 623038 96160 623044 96172
rect 623096 96160 623102 96212
rect 640794 96160 640800 96212
rect 640852 96200 640858 96212
rect 663702 96200 663708 96212
rect 640852 96172 663708 96200
rect 640852 96160 640858 96172
rect 663702 96160 663708 96172
rect 663760 96160 663766 96212
rect 583018 96024 583024 96076
rect 583076 96064 583082 96076
rect 600406 96064 600412 96076
rect 583076 96036 600412 96064
rect 583076 96024 583082 96036
rect 600406 96024 600412 96036
rect 600464 96024 600470 96076
rect 607674 96024 607680 96076
rect 607732 96064 607738 96076
rect 620462 96064 620468 96076
rect 607732 96036 620468 96064
rect 607732 96024 607738 96036
rect 620462 96024 620468 96036
rect 620520 96024 620526 96076
rect 620922 96024 620928 96076
rect 620980 96064 620986 96076
rect 626442 96064 626448 96076
rect 620980 96036 626448 96064
rect 620980 96024 620986 96036
rect 626442 96024 626448 96036
rect 626500 96024 626506 96076
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 663242 96064 663248 96076
rect 641588 96036 663248 96064
rect 641588 96024 641594 96036
rect 663242 96024 663248 96036
rect 663300 96024 663306 96076
rect 577498 95888 577504 95940
rect 577556 95928 577562 95940
rect 598934 95928 598940 95940
rect 577556 95900 598940 95928
rect 577556 95888 577562 95900
rect 598934 95888 598940 95900
rect 598992 95888 598998 95940
rect 613562 95888 613568 95940
rect 613620 95928 613626 95940
rect 613620 95900 625154 95928
rect 613620 95888 613626 95900
rect 625126 95656 625154 95900
rect 635458 95888 635464 95940
rect 635516 95928 635522 95940
rect 635516 95900 638632 95928
rect 635516 95888 635522 95900
rect 638604 95792 638632 95900
rect 639322 95888 639328 95940
rect 639380 95928 639386 95940
rect 643922 95928 643928 95940
rect 639380 95900 643928 95928
rect 639380 95888 639386 95900
rect 643922 95888 643928 95900
rect 643980 95888 643986 95940
rect 647694 95888 647700 95940
rect 647752 95928 647758 95940
rect 653398 95928 653404 95940
rect 647752 95900 653404 95928
rect 647752 95888 647758 95900
rect 653398 95888 653404 95900
rect 653456 95888 653462 95940
rect 664622 95928 664628 95940
rect 654106 95900 664628 95928
rect 646038 95792 646044 95804
rect 638604 95764 646044 95792
rect 646038 95752 646044 95764
rect 646096 95752 646102 95804
rect 648890 95752 648896 95804
rect 648948 95792 648954 95804
rect 654106 95792 654134 95900
rect 664622 95888 664628 95900
rect 664680 95888 664686 95940
rect 648948 95764 654134 95792
rect 648948 95752 648954 95764
rect 638126 95656 638132 95668
rect 625126 95628 638132 95656
rect 638126 95616 638132 95628
rect 638184 95616 638190 95668
rect 638310 95616 638316 95668
rect 638368 95616 638374 95668
rect 638586 95616 638592 95668
rect 638644 95656 638650 95668
rect 646222 95656 646228 95668
rect 638644 95628 646228 95656
rect 638644 95616 638650 95628
rect 646222 95616 646228 95628
rect 646280 95616 646286 95668
rect 638328 95452 638356 95616
rect 648522 95520 648528 95532
rect 640306 95492 648528 95520
rect 640306 95452 640334 95492
rect 648522 95480 648528 95492
rect 648580 95480 648586 95532
rect 638328 95424 640334 95452
rect 579522 95004 579528 95056
rect 579580 95044 579586 95056
rect 582374 95044 582380 95056
rect 579580 95016 582380 95044
rect 579580 95004 579586 95016
rect 582374 95004 582380 95016
rect 582432 95004 582438 95056
rect 616506 94596 616512 94648
rect 616564 94636 616570 94648
rect 625338 94636 625344 94648
rect 616564 94608 625344 94636
rect 616564 94596 616570 94608
rect 625338 94596 625344 94608
rect 625396 94596 625402 94648
rect 584398 94460 584404 94512
rect 584456 94500 584462 94512
rect 601878 94500 601884 94512
rect 584456 94472 601884 94500
rect 584456 94460 584462 94472
rect 601878 94460 601884 94472
rect 601936 94460 601942 94512
rect 608410 94460 608416 94512
rect 608468 94500 608474 94512
rect 624418 94500 624424 94512
rect 608468 94472 624424 94500
rect 608468 94460 608474 94472
rect 624418 94460 624424 94472
rect 624476 94460 624482 94512
rect 578510 93780 578516 93832
rect 578568 93820 578574 93832
rect 588722 93820 588728 93832
rect 578568 93792 588728 93820
rect 578568 93780 578574 93792
rect 588722 93780 588728 93792
rect 588780 93780 588786 93832
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 644474 93780 644480 93832
rect 644532 93820 644538 93832
rect 654870 93820 654876 93832
rect 644532 93792 654876 93820
rect 644532 93780 644538 93792
rect 654870 93780 654876 93792
rect 654928 93780 654934 93832
rect 580442 93100 580448 93152
rect 580500 93140 580506 93152
rect 590102 93140 590108 93152
rect 580500 93112 590108 93140
rect 580500 93100 580506 93112
rect 590102 93100 590108 93112
rect 590160 93100 590166 93152
rect 664438 92488 664444 92540
rect 664496 92528 664502 92540
rect 668302 92528 668308 92540
rect 664496 92500 668308 92528
rect 664496 92488 664502 92500
rect 668302 92488 668308 92500
rect 668360 92488 668366 92540
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 625430 92460 625436 92472
rect 618036 92432 625436 92460
rect 618036 92420 618042 92432
rect 625430 92420 625436 92432
rect 625488 92420 625494 92472
rect 648522 92420 648528 92472
rect 648580 92460 648586 92472
rect 655422 92460 655428 92472
rect 648580 92432 655428 92460
rect 648580 92420 648586 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 617334 91032 617340 91044
rect 611320 91004 617340 91032
rect 611320 90992 611326 91004
rect 617334 90992 617340 91004
rect 617392 90992 617398 91044
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 579062 89700 579068 89752
rect 579120 89740 579126 89752
rect 580626 89740 580632 89752
rect 579120 89712 580632 89740
rect 579120 89700 579126 89712
rect 580626 89700 580632 89712
rect 580684 89700 580690 89752
rect 620462 89632 620468 89684
rect 620520 89672 620526 89684
rect 626442 89672 626448 89684
rect 620520 89644 626448 89672
rect 620520 89632 620526 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 645762 88748 645768 88800
rect 645820 88788 645826 88800
rect 657446 88788 657452 88800
rect 645820 88760 657452 88788
rect 645820 88748 645826 88760
rect 657446 88748 657452 88760
rect 657504 88748 657510 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 579522 88272 579528 88324
rect 579580 88312 579586 88324
rect 587158 88312 587164 88324
rect 579580 88284 587164 88312
rect 579580 88272 579586 88284
rect 587158 88272 587164 88284
rect 587216 88272 587222 88324
rect 607214 88272 607220 88324
rect 607272 88312 607278 88324
rect 626442 88312 626448 88324
rect 607272 88284 626448 88312
rect 607272 88272 607278 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655054 88272 655060 88324
rect 655112 88312 655118 88324
rect 658458 88312 658464 88324
rect 655112 88284 658464 88312
rect 655112 88272 655118 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 617334 88136 617340 88188
rect 617392 88176 617398 88188
rect 625614 88176 625620 88188
rect 617392 88148 625620 88176
rect 617392 88136 617398 88148
rect 625614 88136 625620 88148
rect 625672 88136 625678 88188
rect 647878 87116 647884 87168
rect 647936 87156 647942 87168
rect 657170 87156 657176 87168
rect 647936 87128 657176 87156
rect 647936 87116 647942 87128
rect 657170 87116 657176 87128
rect 657228 87116 657234 87168
rect 650822 86980 650828 87032
rect 650880 87020 650886 87032
rect 661402 87020 661408 87032
rect 650880 86992 661408 87020
rect 650880 86980 650886 86992
rect 661402 86980 661408 86992
rect 661460 86980 661466 87032
rect 649258 86844 649264 86896
rect 649316 86884 649322 86896
rect 660666 86884 660672 86896
rect 649316 86856 660672 86884
rect 649316 86844 649322 86856
rect 660666 86844 660672 86856
rect 660724 86844 660730 86896
rect 578510 86708 578516 86760
rect 578568 86748 578574 86760
rect 580258 86748 580264 86760
rect 578568 86720 580264 86748
rect 578568 86708 578574 86720
rect 580258 86708 580264 86720
rect 580316 86708 580322 86760
rect 650638 86708 650644 86760
rect 650696 86748 650702 86760
rect 658826 86748 658832 86760
rect 650696 86720 658832 86748
rect 650696 86708 650702 86720
rect 658826 86708 658832 86720
rect 658884 86708 658890 86760
rect 659562 86708 659568 86760
rect 659620 86748 659626 86760
rect 663426 86748 663432 86760
rect 659620 86720 663432 86748
rect 659620 86708 659626 86720
rect 663426 86708 663432 86720
rect 663484 86708 663490 86760
rect 652018 86572 652024 86624
rect 652076 86612 652082 86624
rect 662506 86612 662512 86624
rect 652076 86584 662512 86612
rect 652076 86572 652082 86584
rect 662506 86572 662512 86584
rect 662564 86572 662570 86624
rect 623038 86436 623044 86488
rect 623096 86476 623102 86488
rect 626442 86476 626448 86488
rect 623096 86448 626448 86476
rect 623096 86436 623102 86448
rect 626442 86436 626448 86448
rect 626500 86436 626506 86488
rect 653398 86436 653404 86488
rect 653456 86476 653462 86488
rect 660114 86476 660120 86488
rect 653456 86448 660120 86476
rect 653456 86436 653462 86448
rect 660114 86436 660120 86448
rect 660172 86436 660178 86488
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 621658 84124 621664 84176
rect 621716 84164 621722 84176
rect 625614 84164 625620 84176
rect 621716 84136 625620 84164
rect 621716 84124 621722 84136
rect 625614 84124 625620 84136
rect 625672 84124 625678 84176
rect 579338 83988 579344 84040
rect 579396 84028 579402 84040
rect 581822 84028 581828 84040
rect 579396 84000 581828 84028
rect 579396 83988 579402 84000
rect 581822 83988 581828 84000
rect 581880 83988 581886 84040
rect 579246 82764 579252 82816
rect 579304 82804 579310 82816
rect 588538 82804 588544 82816
rect 579304 82776 588544 82804
rect 579304 82764 579310 82776
rect 588538 82764 588544 82776
rect 588596 82764 588602 82816
rect 628650 80928 628656 80980
rect 628708 80968 628714 80980
rect 642450 80968 642456 80980
rect 628708 80940 642456 80968
rect 628708 80928 628714 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 614022 80792 614028 80844
rect 614080 80832 614086 80844
rect 647326 80832 647332 80844
rect 614080 80804 647332 80832
rect 614080 80792 614086 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636102 80696 636108 80708
rect 595496 80668 636108 80696
rect 595496 80656 595502 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 579246 80044 579252 80096
rect 579304 80084 579310 80096
rect 585962 80084 585968 80096
rect 579304 80056 585968 80084
rect 579304 80044 579310 80056
rect 585962 80044 585968 80056
rect 586020 80044 586026 80096
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 638862 79472 638868 79484
rect 629260 79444 638868 79472
rect 629260 79432 629266 79444
rect 638862 79432 638868 79444
rect 638920 79432 638926 79484
rect 616138 79296 616144 79348
rect 616196 79336 616202 79348
rect 648982 79336 648988 79348
rect 616196 79308 648988 79336
rect 616196 79296 616202 79308
rect 648982 79296 648988 79308
rect 649040 79296 649046 79348
rect 638862 78276 638868 78328
rect 638920 78316 638926 78328
rect 645302 78316 645308 78328
rect 638920 78288 645308 78316
rect 638920 78276 638926 78288
rect 645302 78276 645308 78288
rect 645360 78276 645366 78328
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 639046 78112 639052 78124
rect 631100 78084 639052 78112
rect 631100 78072 631106 78084
rect 639046 78072 639052 78084
rect 639104 78072 639110 78124
rect 612642 77936 612648 77988
rect 612700 77976 612706 77988
rect 647510 77976 647516 77988
rect 612700 77948 647516 77976
rect 612700 77936 612706 77948
rect 647510 77936 647516 77948
rect 647568 77936 647574 77988
rect 628190 77528 628196 77580
rect 628248 77568 628254 77580
rect 633894 77568 633900 77580
rect 628248 77540 633900 77568
rect 628248 77528 628254 77540
rect 633894 77528 633900 77540
rect 633952 77528 633958 77580
rect 578878 77392 578884 77444
rect 578936 77432 578942 77444
rect 631042 77432 631048 77444
rect 578936 77404 631048 77432
rect 578936 77392 578942 77404
rect 631042 77392 631048 77404
rect 631100 77392 631106 77444
rect 589918 77256 589924 77308
rect 589976 77296 589982 77308
rect 628190 77296 628196 77308
rect 589976 77268 628196 77296
rect 589976 77256 589982 77268
rect 628190 77256 628196 77268
rect 628248 77256 628254 77308
rect 628374 77256 628380 77308
rect 628432 77296 628438 77308
rect 631502 77296 631508 77308
rect 628432 77268 631508 77296
rect 628432 77256 628438 77268
rect 631502 77256 631508 77268
rect 631560 77256 631566 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 649166 76820 649172 76832
rect 620336 76792 649172 76820
rect 620336 76780 620342 76792
rect 649166 76780 649172 76792
rect 649224 76780 649230 76832
rect 611998 76644 612004 76696
rect 612056 76684 612062 76696
rect 647050 76684 647056 76696
rect 612056 76656 647056 76684
rect 612056 76644 612062 76656
rect 647050 76644 647056 76656
rect 647108 76644 647114 76696
rect 606478 76508 606484 76560
rect 606536 76548 606542 76560
rect 662414 76548 662420 76560
rect 606536 76520 662420 76548
rect 606536 76508 606542 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 579246 75556 579252 75608
rect 579304 75596 579310 75608
rect 581638 75596 581644 75608
rect 579304 75568 581644 75596
rect 579304 75556 579310 75568
rect 581638 75556 581644 75568
rect 581696 75556 581702 75608
rect 618898 75148 618904 75200
rect 618956 75188 618962 75200
rect 646866 75188 646872 75200
rect 618956 75160 646872 75188
rect 618956 75148 618962 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 588538 74808 588544 74860
rect 588596 74848 588602 74860
rect 628006 74848 628012 74860
rect 588596 74820 628012 74848
rect 588596 74808 588602 74820
rect 628006 74808 628012 74820
rect 628064 74808 628070 74860
rect 578602 73108 578608 73160
rect 578660 73148 578666 73160
rect 580442 73148 580448 73160
rect 578660 73120 580448 73148
rect 578660 73108 578666 73120
rect 580442 73108 580448 73120
rect 580500 73108 580506 73160
rect 579522 67600 579528 67652
rect 579580 67640 579586 67652
rect 624418 67640 624424 67652
rect 579580 67612 624424 67640
rect 579580 67600 579586 67612
rect 624418 67600 624424 67612
rect 624476 67600 624482 67652
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 605834 66280 605840 66292
rect 579580 66252 605840 66280
rect 579580 66240 579586 66252
rect 605834 66240 605840 66252
rect 605892 66240 605898 66292
rect 581638 65492 581644 65544
rect 581696 65532 581702 65544
rect 603074 65532 603080 65544
rect 581696 65504 603080 65532
rect 581696 65492 581702 65504
rect 603074 65492 603080 65504
rect 603132 65492 603138 65544
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 613378 64852 613384 64864
rect 579580 64824 613384 64852
rect 579580 64812 579586 64824
rect 613378 64812 613384 64824
rect 613436 64812 613442 64864
rect 580258 62772 580264 62824
rect 580316 62812 580322 62824
rect 601878 62812 601884 62824
rect 580316 62784 601884 62812
rect 580316 62772 580322 62784
rect 601878 62772 601884 62784
rect 601936 62772 601942 62824
rect 578510 62024 578516 62076
rect 578568 62064 578574 62076
rect 664438 62064 664444 62076
rect 578568 62036 664444 62064
rect 578568 62024 578574 62036
rect 664438 62024 664444 62036
rect 664496 62024 664502 62076
rect 579522 60664 579528 60716
rect 579580 60704 579586 60716
rect 614850 60704 614856 60716
rect 579580 60676 614856 60704
rect 579580 60664 579586 60676
rect 614850 60664 614856 60676
rect 614908 60664 614914 60716
rect 579062 58624 579068 58676
rect 579120 58664 579126 58676
rect 600498 58664 600504 58676
rect 579120 58636 600504 58664
rect 579120 58624 579126 58636
rect 600498 58624 600504 58636
rect 600556 58624 600562 58676
rect 605834 58624 605840 58676
rect 605892 58664 605898 58676
rect 663794 58664 663800 58676
rect 605892 58636 663800 58664
rect 605892 58624 605898 58636
rect 663794 58624 663800 58636
rect 663852 58624 663858 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 666554 57916 666560 57928
rect 579580 57888 666560 57916
rect 579580 57876 579586 57888
rect 666554 57876 666560 57888
rect 666612 57876 666618 57928
rect 579522 56516 579528 56568
rect 579580 56556 579586 56568
rect 588538 56556 588544 56568
rect 579580 56528 588544 56556
rect 579580 56516 579586 56528
rect 588538 56516 588544 56528
rect 588596 56516 588602 56568
rect 574922 56108 574928 56160
rect 574980 56148 574986 56160
rect 596450 56148 596456 56160
rect 574980 56120 596456 56148
rect 574980 56108 574986 56120
rect 596450 56108 596456 56120
rect 596508 56108 596514 56160
rect 574554 55972 574560 56024
rect 574612 56012 574618 56024
rect 596174 56012 596180 56024
rect 574612 55984 596180 56012
rect 574612 55972 574618 55984
rect 596174 55972 596180 55984
rect 596232 55972 596238 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 599118 55876 599124 55888
rect 574796 55848 599124 55876
rect 574796 55836 574802 55848
rect 599118 55836 599124 55848
rect 599176 55836 599182 55888
rect 624418 55836 624424 55888
rect 624476 55876 624482 55888
rect 663978 55876 663984 55888
rect 624476 55848 663984 55876
rect 624476 55836 624482 55848
rect 663978 55836 663984 55848
rect 664036 55836 664042 55888
rect 465046 55576 478874 55604
rect 465046 55196 465074 55576
rect 459480 55168 465074 55196
rect 465644 55440 478184 55468
rect 459480 53644 459508 55168
rect 465644 55060 465672 55440
rect 465000 55032 465672 55060
rect 465736 55304 474596 55332
rect 465000 54720 465028 55032
rect 464908 54692 465028 54720
rect 459462 53592 459468 53644
rect 459520 53592 459526 53644
rect 464908 53632 464936 54692
rect 465736 53644 465764 55304
rect 474568 55060 474596 55304
rect 478156 55060 478184 55440
rect 478846 55196 478874 55576
rect 577498 55196 577504 55208
rect 478846 55168 577504 55196
rect 577498 55156 577504 55168
rect 577556 55156 577562 55208
rect 585778 55060 585784 55072
rect 469784 55032 474504 55060
rect 474568 55032 474734 55060
rect 478156 55032 585784 55060
rect 465166 53632 465172 53644
rect 464908 53604 465172 53632
rect 465166 53592 465172 53604
rect 465224 53592 465230 53644
rect 465718 53592 465724 53644
rect 465776 53592 465782 53644
rect 465902 53592 465908 53644
rect 465960 53632 465966 53644
rect 469784 53632 469812 55032
rect 474476 54788 474504 55032
rect 474706 54924 474734 55032
rect 585778 55020 585784 55032
rect 585836 55020 585842 55072
rect 583018 54924 583024 54936
rect 474706 54896 583024 54924
rect 583018 54884 583024 54896
rect 583076 54884 583082 54936
rect 589918 54788 589924 54800
rect 469968 54760 474412 54788
rect 474476 54760 589924 54788
rect 469968 53644 469996 54760
rect 474384 54652 474412 54760
rect 589918 54748 589924 54760
rect 589976 54748 589982 54800
rect 597830 54652 597836 54664
rect 474384 54624 597836 54652
rect 597830 54612 597836 54624
rect 597888 54612 597894 54664
rect 597646 54516 597652 54528
rect 470152 54488 597652 54516
rect 470152 53644 470180 54488
rect 597646 54476 597652 54488
rect 597704 54476 597710 54528
rect 578878 54380 578884 54392
rect 474200 54352 578884 54380
rect 474200 54312 474228 54352
rect 578878 54340 578884 54352
rect 578936 54340 578942 54392
rect 474108 54284 474228 54312
rect 474108 53904 474136 54284
rect 579062 54244 579068 54256
rect 470428 53876 474136 53904
rect 477972 54216 579068 54244
rect 470428 53644 470456 53876
rect 470612 53740 473354 53768
rect 465960 53604 469812 53632
rect 465960 53592 465966 53604
rect 469950 53592 469956 53644
rect 470008 53592 470014 53644
rect 470134 53592 470140 53644
rect 470192 53592 470198 53644
rect 470410 53592 470416 53644
rect 470468 53592 470474 53644
rect 461302 53456 461308 53508
rect 461360 53496 461366 53508
rect 470612 53496 470640 53740
rect 473326 53632 473354 53740
rect 477972 53644 478000 54216
rect 579062 54204 579068 54216
rect 579120 54204 579126 54256
rect 574738 54108 574744 54120
rect 478156 54080 574744 54108
rect 473326 53604 474320 53632
rect 461360 53468 470640 53496
rect 474292 53496 474320 53604
rect 477954 53592 477960 53644
rect 478012 53592 478018 53644
rect 478156 53496 478184 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 574554 53972 574560 53984
rect 481744 53944 574560 53972
rect 481744 53644 481772 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 482986 53808 574928 53836
rect 481726 53592 481732 53644
rect 481784 53592 481790 53644
rect 482002 53592 482008 53644
rect 482060 53632 482066 53644
rect 482986 53632 483014 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 482060 53604 483014 53632
rect 482060 53592 482066 53604
rect 474292 53468 478184 53496
rect 461360 53456 461366 53468
rect 50522 53320 50528 53372
rect 50580 53360 50586 53372
rect 128998 53360 129004 53372
rect 50580 53332 129004 53360
rect 50580 53320 50586 53332
rect 128998 53320 129004 53332
rect 129056 53320 129062 53372
rect 463602 53320 463608 53372
rect 463660 53360 463666 53372
rect 470134 53360 470140 53372
rect 463660 53332 470140 53360
rect 463660 53320 463666 53332
rect 470134 53320 470140 53332
rect 470192 53320 470198 53372
rect 47762 53184 47768 53236
rect 47820 53224 47826 53236
rect 130378 53224 130384 53236
rect 47820 53196 130384 53224
rect 47820 53184 47826 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 463142 53184 463148 53236
rect 463200 53224 463206 53236
rect 477954 53224 477960 53236
rect 463200 53196 477960 53224
rect 463200 53184 463206 53196
rect 477954 53184 477960 53196
rect 478012 53184 478018 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 130562 53088 130568 53100
rect 46256 53060 130568 53088
rect 46256 53048 46262 53060
rect 130562 53048 130568 53060
rect 130620 53048 130626 53100
rect 464890 53048 464896 53100
rect 464948 53088 464954 53100
rect 481726 53088 481732 53100
rect 464948 53060 481732 53088
rect 464948 53048 464954 53060
rect 481726 53048 481732 53060
rect 481784 53048 481790 53100
rect 464062 52912 464068 52964
rect 464120 52952 464126 52964
rect 482002 52952 482008 52964
rect 464120 52924 482008 52952
rect 464120 52912 464126 52924
rect 482002 52912 482008 52924
rect 482060 52912 482066 52964
rect 460060 52776 460066 52828
rect 460118 52816 460124 52828
rect 460118 52788 462314 52816
rect 460118 52776 460124 52788
rect 462286 52680 462314 52788
rect 464200 52776 464206 52828
rect 464258 52816 464264 52828
rect 469950 52816 469956 52828
rect 464258 52788 469956 52816
rect 464258 52776 464264 52788
rect 469950 52776 469956 52788
rect 470008 52776 470014 52828
rect 470410 52680 470416 52692
rect 462286 52652 470416 52680
rect 470410 52640 470416 52652
rect 470468 52640 470474 52692
rect 145374 52436 145380 52488
rect 145432 52476 145438 52488
rect 306006 52476 306012 52488
rect 145432 52448 306012 52476
rect 145432 52436 145438 52448
rect 306006 52436 306012 52448
rect 306064 52436 306070 52488
rect 50706 51960 50712 52012
rect 50764 52000 50770 52012
rect 130746 52000 130752 52012
rect 50764 51972 130752 52000
rect 50764 51960 50770 51972
rect 130746 51960 130752 51972
rect 130804 51960 130810 52012
rect 49142 51824 49148 51876
rect 49200 51864 49206 51876
rect 127158 51864 127164 51876
rect 49200 51836 127164 51864
rect 49200 51824 49206 51836
rect 127158 51824 127164 51836
rect 127216 51824 127222 51876
rect 48958 51688 48964 51740
rect 49016 51728 49022 51740
rect 129458 51728 129464 51740
rect 49016 51700 129464 51728
rect 49016 51688 49022 51700
rect 129458 51688 129464 51700
rect 129516 51688 129522 51740
rect 127158 50736 127164 50788
rect 127216 50776 127222 50788
rect 129274 50776 129280 50788
rect 127216 50748 129280 50776
rect 127216 50736 127222 50748
rect 129274 50736 129280 50748
rect 129332 50736 129338 50788
rect 50338 50464 50344 50516
rect 50396 50504 50402 50516
rect 128630 50504 128636 50516
rect 50396 50476 128636 50504
rect 50396 50464 50402 50476
rect 128630 50464 128636 50476
rect 128688 50464 128694 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 128998 50368 129004 50380
rect 45520 50340 129004 50368
rect 45520 50328 45526 50340
rect 128998 50328 129004 50340
rect 129056 50328 129062 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 128446 49144 128452 49156
rect 51776 49116 128452 49144
rect 51776 49104 51782 49116
rect 128446 49104 128452 49116
rect 128504 49104 128510 49156
rect 47578 48968 47584 49020
rect 47636 49008 47642 49020
rect 129642 49008 129648 49020
rect 47636 48980 129648 49008
rect 47636 48968 47642 48980
rect 129642 48968 129648 48980
rect 129700 48968 129706 49020
rect 128630 47812 128636 47864
rect 128688 47852 128694 47864
rect 132126 47852 132132 47864
rect 128688 47824 132132 47852
rect 128688 47812 128694 47824
rect 132126 47812 132132 47824
rect 132184 47812 132190 47864
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 130856 45064 131146 45076
rect 129608 45048 131146 45064
rect 129608 45036 130884 45048
rect 129608 45024 129614 45036
rect 131316 44964 131376 44992
rect 129734 44888 129740 44940
rect 129792 44928 129798 44940
rect 131316 44928 131344 44964
rect 129792 44900 131344 44928
rect 129792 44888 129798 44900
rect 131500 44880 131560 44908
rect 131500 44860 131528 44880
rect 131454 44832 131528 44860
rect 131454 44824 131482 44832
rect 128446 44752 128452 44804
rect 128504 44792 128510 44804
rect 131362 44796 131482 44824
rect 131684 44796 131790 44824
rect 131362 44792 131390 44796
rect 131684 44792 131712 44796
rect 128504 44764 131390 44792
rect 131592 44764 131712 44792
rect 128504 44752 128510 44764
rect 129366 44548 129372 44600
rect 129424 44588 129430 44600
rect 131592 44588 131620 44764
rect 131960 44724 131988 44726
rect 129424 44560 131620 44588
rect 131868 44696 131988 44724
rect 131868 44572 131896 44696
rect 129424 44548 129430 44560
rect 131776 44544 131896 44572
rect 129182 44412 129188 44464
rect 129240 44452 129246 44464
rect 131776 44452 131804 44544
rect 132236 44520 132264 44642
rect 132144 44500 132264 44520
rect 129240 44424 131804 44452
rect 132126 44448 132132 44500
rect 132184 44492 132264 44500
rect 132184 44448 132190 44492
rect 132420 44464 132448 44558
rect 129240 44412 129246 44424
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 130746 44276 130752 44328
rect 130804 44316 130810 44328
rect 132604 44316 132632 44474
rect 130804 44288 132632 44316
rect 130804 44276 130810 44288
rect 128998 44140 129004 44192
rect 129056 44180 129062 44192
rect 132218 44180 132224 44192
rect 129056 44152 132224 44180
rect 129056 44140 129062 44152
rect 132218 44140 132224 44152
rect 132276 44140 132282 44192
rect 132788 44180 132816 44362
rect 132420 44152 132816 44180
rect 130562 44004 130568 44056
rect 130620 44044 130626 44056
rect 132420 44044 132448 44152
rect 130620 44016 132448 44044
rect 130620 44004 130626 44016
rect 130378 43868 130384 43920
rect 130436 43908 130442 43920
rect 132972 43908 133000 44250
rect 130436 43880 133000 43908
rect 130436 43868 130442 43880
rect 43438 42780 43444 42832
rect 43496 42820 43502 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43496 42792 133184 42820
rect 43496 42780 43502 42792
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 307352 42724 369256 42752
rect 307352 42712 307358 42724
rect 369228 42616 369256 42724
rect 369394 42712 369400 42764
rect 369452 42752 369458 42764
rect 431218 42752 431224 42764
rect 369452 42724 431224 42752
rect 369452 42712 369458 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 464338 42752 464344 42764
rect 456116 42724 464344 42752
rect 456116 42712 456122 42724
rect 464338 42712 464344 42724
rect 464396 42712 464402 42764
rect 427078 42616 427084 42628
rect 369228 42588 427084 42616
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 455874 42576 455880 42628
rect 455932 42616 455938 42628
rect 463970 42616 463976 42628
rect 455932 42588 463976 42616
rect 455932 42576 455938 42588
rect 463970 42576 463976 42588
rect 464028 42576 464034 42628
rect 361758 42440 361764 42492
rect 361816 42480 361822 42492
rect 369394 42480 369400 42492
rect 361816 42452 369400 42480
rect 361816 42440 361822 42452
rect 369394 42440 369400 42452
rect 369452 42440 369458 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 308950 42173 308956 42225
rect 309008 42173 309014 42225
rect 427078 42032 427084 42084
rect 427136 42072 427142 42084
rect 427136 42044 427814 42072
rect 427136 42032 427142 42044
rect 427786 41936 427814 42044
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 455874 41936 455880 41948
rect 427786 41908 455880 41936
rect 455874 41896 455880 41908
rect 455932 41896 455938 41948
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 106832 1007292 106884 1007344
rect 113824 1007360 113876 1007412
rect 425520 1007088 425572 1007140
rect 359740 1006952 359792 1007004
rect 371240 1006952 371292 1007004
rect 428372 1006884 428424 1006936
rect 359372 1006816 359424 1006868
rect 367376 1006816 367428 1006868
rect 429200 1006748 429252 1006800
rect 431868 1006748 431920 1006800
rect 440240 1006748 440292 1006800
rect 161756 1006680 161808 1006732
rect 164884 1006680 164936 1006732
rect 361396 1006680 361448 1006732
rect 376024 1006680 376076 1006732
rect 94504 1006544 94556 1006596
rect 101956 1006544 102008 1006596
rect 145564 1006544 145616 1006596
rect 153752 1006544 153804 1006596
rect 157432 1006544 157484 1006596
rect 162308 1006544 162360 1006596
rect 162492 1006544 162544 1006596
rect 173164 1006544 173216 1006596
rect 101588 1006408 101640 1006460
rect 104808 1006408 104860 1006460
rect 145748 1006408 145800 1006460
rect 152924 1006408 152976 1006460
rect 158260 1006408 158312 1006460
rect 171784 1006408 171836 1006460
rect 247868 1006408 247920 1006460
rect 256148 1006408 256200 1006460
rect 301504 1006408 301556 1006460
rect 307760 1006408 307812 1006460
rect 360568 1006408 360620 1006460
rect 367008 1006408 367060 1006460
rect 402244 1006408 402296 1006460
rect 431684 1006612 431736 1006664
rect 507860 1006884 507912 1006936
rect 520924 1006816 520976 1006868
rect 505008 1006680 505060 1006732
rect 518164 1006680 518216 1006732
rect 555976 1006680 556028 1006732
rect 558828 1006680 558880 1006732
rect 467104 1006544 467156 1006596
rect 501328 1006544 501380 1006596
rect 514760 1006544 514812 1006596
rect 556804 1006544 556856 1006596
rect 567844 1006544 567896 1006596
rect 429200 1006408 429252 1006460
rect 93124 1006272 93176 1006324
rect 100300 1006272 100352 1006324
rect 144276 1006272 144328 1006324
rect 93308 1006136 93360 1006188
rect 94688 1006000 94740 1006052
rect 98276 1006000 98328 1006052
rect 101404 1006136 101456 1006188
rect 103980 1006136 104032 1006188
rect 106004 1006136 106056 1006188
rect 124864 1006136 124916 1006188
rect 144736 1006136 144788 1006188
rect 151268 1006136 151320 1006188
rect 158628 1006272 158680 1006324
rect 162492 1006272 162544 1006324
rect 255964 1006272 256016 1006324
rect 259000 1006272 259052 1006324
rect 300492 1006272 300544 1006324
rect 306932 1006272 306984 1006324
rect 314660 1006272 314712 1006324
rect 319444 1006272 319496 1006324
rect 354864 1006272 354916 1006324
rect 360844 1006272 360896 1006324
rect 367376 1006272 367428 1006324
rect 380164 1006272 380216 1006324
rect 423496 1006272 423548 1006324
rect 429108 1006272 429160 1006324
rect 152096 1006136 152148 1006188
rect 160284 1006136 160336 1006188
rect 161756 1006136 161808 1006188
rect 162308 1006136 162360 1006188
rect 175924 1006136 175976 1006188
rect 210424 1006136 210476 1006188
rect 228364 1006136 228416 1006188
rect 262680 1006136 262732 1006188
rect 269764 1006136 269816 1006188
rect 298744 1006136 298796 1006188
rect 304908 1006136 304960 1006188
rect 357716 1006136 357768 1006188
rect 362224 1006136 362276 1006188
rect 365076 1006136 365128 1006188
rect 367744 1006136 367796 1006188
rect 553124 1006408 553176 1006460
rect 431868 1006340 431920 1006392
rect 505376 1006272 505428 1006324
rect 102324 1006000 102376 1006052
rect 108488 1006000 108540 1006052
rect 126244 1006000 126296 1006052
rect 148876 1006000 148928 1006052
rect 150072 1006000 150124 1006052
rect 153936 1006000 153988 1006052
rect 158260 1006000 158312 1006052
rect 159456 1006000 159508 1006052
rect 177304 1006000 177356 1006052
rect 198188 1006000 198240 1006052
rect 201040 1006000 201092 1006052
rect 208400 1006000 208452 1006052
rect 229744 1006000 229796 1006052
rect 249064 1006000 249116 1006052
rect 257344 1006000 257396 1006052
rect 261852 1006000 261904 1006052
rect 279424 1006000 279476 1006052
rect 298928 1006000 298980 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 311808 1006000 311860 1006052
rect 314660 1006000 314712 1006052
rect 320824 1006000 320876 1006052
rect 355692 1006000 355744 1006052
rect 359464 1006000 359516 1006052
rect 363420 1006000 363472 1006052
rect 382924 1006000 382976 1006052
rect 400864 1006000 400916 1006052
rect 469864 1006136 469916 1006188
rect 507032 1006136 507084 1006188
rect 509700 1006136 509752 1006188
rect 552296 1006272 552348 1006324
rect 558184 1006272 558236 1006324
rect 570604 1006272 570656 1006324
rect 519544 1006136 519596 1006188
rect 551468 1006136 551520 1006188
rect 557448 1006136 557500 1006188
rect 558828 1006136 558880 1006188
rect 571984 1006136 572036 1006188
rect 423496 1006000 423548 1006052
rect 430304 1006000 430356 1006052
rect 431684 1006000 431736 1006052
rect 471244 1006000 471296 1006052
rect 496728 1006000 496780 1006052
rect 498844 1006000 498896 1006052
rect 502524 1006000 502576 1006052
rect 505744 1006000 505796 1006052
rect 506204 1006000 506256 1006052
rect 509056 1006000 509108 1006052
rect 509240 1006000 509292 1006052
rect 522304 1006000 522356 1006052
rect 555976 1006000 556028 1006052
rect 573364 1006000 573416 1006052
rect 429476 1005796 429528 1005848
rect 426348 1005660 426400 1005712
rect 431868 1005796 431920 1005848
rect 453304 1005796 453356 1005848
rect 509240 1005728 509292 1005780
rect 514024 1005728 514076 1005780
rect 367008 1005524 367060 1005576
rect 377404 1005524 377456 1005576
rect 425520 1005524 425572 1005576
rect 445024 1005660 445076 1005712
rect 360568 1005388 360620 1005440
rect 378784 1005388 378836 1005440
rect 424324 1005388 424376 1005440
rect 429476 1005388 429528 1005440
rect 457444 1005524 457496 1005576
rect 462964 1005388 463016 1005440
rect 552296 1005388 552348 1005440
rect 566648 1005388 566700 1005440
rect 102784 1005252 102836 1005304
rect 108856 1005252 108908 1005304
rect 204904 1005252 204956 1005304
rect 212080 1005252 212132 1005304
rect 356520 1005252 356572 1005304
rect 373264 1005252 373316 1005304
rect 425152 1005252 425204 1005304
rect 468484 1005252 468536 1005304
rect 498844 1005252 498896 1005304
rect 516784 1005252 516836 1005304
rect 551468 1005252 551520 1005304
rect 569224 1005252 569276 1005304
rect 304264 1005184 304316 1005236
rect 307300 1005184 307352 1005236
rect 429108 1005116 429160 1005168
rect 447784 1005116 447836 1005168
rect 149888 1005048 149940 1005100
rect 152924 1005048 152976 1005100
rect 305828 1005048 305880 1005100
rect 308956 1005048 309008 1005100
rect 365076 1005048 365128 1005100
rect 370504 1005048 370556 1005100
rect 508228 1005048 508280 1005100
rect 511264 1005048 511316 1005100
rect 428004 1004980 428056 1005032
rect 431868 1004980 431920 1005032
rect 151084 1004912 151136 1004964
rect 153752 1004912 153804 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 263048 1004912 263100 1004964
rect 268384 1004912 268436 1004964
rect 353208 1004912 353260 1004964
rect 355692 1004912 355744 1004964
rect 361396 1004912 361448 1004964
rect 364984 1004912 365036 1004964
rect 497924 1004912 497976 1004964
rect 500500 1004912 500552 1004964
rect 149704 1004776 149756 1004828
rect 151728 1004776 151780 1004828
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 211252 1004776 211304 1004828
rect 215944 1004776 215996 1004828
rect 258172 1004776 258224 1004828
rect 259460 1004776 259512 1004828
rect 305644 1004776 305696 1004828
rect 308128 1004776 308180 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 354588 1004776 354640 1004828
rect 356520 1004776 356572 1004828
rect 362592 1004776 362644 1004828
rect 365168 1004776 365220 1004828
rect 420828 1004776 420880 1004828
rect 422668 1004776 422720 1004828
rect 498108 1004776 498160 1004828
rect 499672 1004776 499724 1004828
rect 508228 1004776 508280 1004828
rect 510804 1004776 510856 1004828
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 151268 1004640 151320 1004692
rect 154120 1004640 154172 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 304908 1004640 304960 1004692
rect 306932 1004640 306984 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 432880 1004640 432932 1004692
rect 438124 1004640 438176 1004692
rect 499488 1004640 499540 1004692
rect 500500 1004640 500552 1004692
rect 507400 1004640 507452 1004692
rect 509240 1004640 509292 1004692
rect 560852 1004640 560904 1004692
rect 566464 1004640 566516 1004692
rect 504548 1004368 504600 1004420
rect 510988 1004368 511040 1004420
rect 426348 1004028 426400 1004080
rect 455880 1004028 455932 1004080
rect 92296 1003892 92348 1003944
rect 103152 1003892 103204 1003944
rect 247316 1003892 247368 1003944
rect 255320 1003892 255372 1003944
rect 421840 1003892 421892 1003944
rect 464344 1003892 464396 1003944
rect 557172 1003892 557224 1003944
rect 571248 1003892 571300 1003944
rect 300308 1003280 300360 1003332
rect 305276 1003280 305328 1003332
rect 501696 1003280 501748 1003332
rect 504732 1003280 504784 1003332
rect 371240 1002940 371292 1002992
rect 374368 1002940 374420 1002992
rect 253112 1002668 253164 1002720
rect 256148 1002668 256200 1002720
rect 98644 1002600 98696 1002652
rect 101956 1002600 102008 1002652
rect 302240 1002600 302292 1002652
rect 304908 1002600 304960 1002652
rect 246580 1002532 246632 1002584
rect 254124 1002532 254176 1002584
rect 440240 1002532 440292 1002584
rect 466368 1002532 466420 1002584
rect 97448 1002464 97500 1002516
rect 100300 1002464 100352 1002516
rect 261024 1002464 261076 1002516
rect 264244 1002464 264296 1002516
rect 560852 1002464 560904 1002516
rect 565084 1002464 565136 1002516
rect 96068 1002328 96120 1002380
rect 99104 1002328 99156 1002380
rect 107660 1002328 107712 1002380
rect 109500 1002328 109552 1002380
rect 148508 1002328 148560 1002380
rect 150900 1002328 150952 1002380
rect 251824 1002328 251876 1002380
rect 254492 1002328 254544 1002380
rect 260196 1002328 260248 1002380
rect 262864 1002328 262916 1002380
rect 503352 1002328 503404 1002380
rect 506480 1002328 506532 1002380
rect 551928 1002328 551980 1002380
rect 553952 1002328 554004 1002380
rect 560484 1002328 560536 1002380
rect 563060 1002328 563112 1002380
rect 98828 1002192 98880 1002244
rect 101128 1002192 101180 1002244
rect 105636 1002192 105688 1002244
rect 107844 1002192 107896 1002244
rect 108028 1002192 108080 1002244
rect 110420 1002192 110472 1002244
rect 155776 1002192 155828 1002244
rect 157340 1002192 157392 1002244
rect 203340 1002192 203392 1002244
rect 206376 1002192 206428 1002244
rect 206744 1002192 206796 1002244
rect 208584 1002192 208636 1002244
rect 254584 1002192 254636 1002244
rect 256516 1002192 256568 1002244
rect 259828 1002192 259880 1002244
rect 262220 1002192 262272 1002244
rect 303252 1002192 303304 1002244
rect 306104 1002192 306156 1002244
rect 308404 1002192 308456 1002244
rect 310612 1002192 310664 1002244
rect 355324 1002192 355376 1002244
rect 358544 1002192 358596 1002244
rect 553308 1002192 553360 1002244
rect 555148 1002192 555200 1002244
rect 97264 1002056 97316 1002108
rect 99472 1002056 99524 1002108
rect 100024 1002056 100076 1002108
rect 103152 1002056 103204 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111800 1002056 111852 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 152464 1002056 152516 1002108
rect 154580 1002056 154632 1002108
rect 157800 1002056 157852 1002108
rect 160100 1002056 160152 1002108
rect 205088 1002056 205140 1002108
rect 207204 1002056 207256 1002108
rect 210884 1002056 210936 1002108
rect 213184 1002056 213236 1002108
rect 253388 1002056 253440 1002108
rect 255320 1002056 255372 1002108
rect 261024 1002056 261076 1002108
rect 95884 1001920 95936 1001972
rect 98276 1001920 98328 1001972
rect 99012 1001920 99064 1001972
rect 101128 1001920 101180 1001972
rect 106004 1001920 106056 1001972
rect 107752 1001920 107804 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 156604 1001920 156656 1001972
rect 158720 1001920 158772 1001972
rect 195152 1001920 195204 1001972
rect 202696 1001920 202748 1001972
rect 203708 1001920 203760 1001972
rect 205548 1001920 205600 1001972
rect 212540 1001920 212592 1001972
rect 214564 1001920 214616 1001972
rect 254768 1001920 254820 1001972
rect 256976 1001920 257028 1001972
rect 260196 1001920 260248 1001972
rect 260932 1001920 260984 1001972
rect 263508 1002056 263560 1002108
rect 265624 1002056 265676 1002108
rect 300124 1002056 300176 1002108
rect 304080 1002056 304132 1002108
rect 355784 1002056 355836 1002108
rect 357716 1002056 357768 1002108
rect 503352 1002056 503404 1002108
rect 506296 1002056 506348 1002108
rect 509884 1002056 509936 1002108
rect 515404 1002056 515456 1002108
rect 427544 1001988 427596 1002040
rect 431868 1001988 431920 1002040
rect 263600 1001920 263652 1001972
rect 263876 1001920 263928 1001972
rect 267004 1001920 267056 1001972
rect 302884 1001920 302936 1001972
rect 306104 1001920 306156 1001972
rect 307024 1001920 307076 1001972
rect 308956 1001920 309008 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 360200 1001920 360252 1001972
rect 363604 1001920 363656 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 423588 1001920 423640 1001972
rect 424324 1001920 424376 1001972
rect 500868 1001920 500920 1001972
rect 501696 1001920 501748 1001972
rect 502156 1001920 502208 1001972
rect 504180 1001920 504232 1001972
rect 505376 1001920 505428 1001972
rect 508504 1001920 508556 1001972
rect 510344 1001920 510396 1001972
rect 512644 1001920 512696 1001972
rect 552664 1001920 552716 1001972
rect 554320 1001920 554372 1001972
rect 561680 1001920 561732 1001972
rect 563704 1001920 563756 1001972
rect 551100 1001308 551152 1001360
rect 568488 1001308 568540 1001360
rect 195520 1001172 195572 1001224
rect 203892 1001172 203944 1001224
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 423588 1001172 423640 1001224
rect 440240 1001172 440292 1001224
rect 498108 1001172 498160 1001224
rect 521292 1001172 521344 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 298284 1000492 298336 1000544
rect 305828 1000492 305880 1000544
rect 427176 1000492 427228 1000544
rect 430488 1000492 430540 1000544
rect 247132 999744 247184 999796
rect 254768 999744 254820 999796
rect 430304 999744 430356 999796
rect 443644 999744 443696 999796
rect 514760 999268 514812 999320
rect 95148 999132 95200 999184
rect 99012 999132 99064 999184
rect 506480 999132 506532 999184
rect 517428 999132 517480 999184
rect 555148 999132 555200 999184
rect 556160 999132 556212 999184
rect 618168 999132 618220 999184
rect 625252 999132 625304 999184
rect 523500 999064 523552 999116
rect 457444 998928 457496 998980
rect 472624 998928 472676 998980
rect 504732 998928 504784 998980
rect 517704 998928 517756 998980
rect 92296 998792 92348 998844
rect 92940 998792 92992 998844
rect 428372 998792 428424 998844
rect 436100 998792 436152 998844
rect 453304 998792 453356 998844
rect 472440 998792 472492 998844
rect 517244 998792 517296 998844
rect 522120 998792 522172 998844
rect 196808 998656 196860 998708
rect 204352 998656 204404 998708
rect 357440 998656 357492 998708
rect 383292 998724 383344 998776
rect 502156 998724 502208 998776
rect 516876 998724 516928 998776
rect 430488 998656 430540 998708
rect 456800 998656 456852 998708
rect 467104 998656 467156 998708
rect 471980 998656 472032 998708
rect 517428 998656 517480 998708
rect 523684 998656 523736 998708
rect 378784 998588 378836 998640
rect 383568 998588 383620 998640
rect 196624 998520 196676 998572
rect 203524 998520 203576 998572
rect 351828 998520 351880 998572
rect 378600 998520 378652 998572
rect 430856 998520 430908 998572
rect 433984 998520 434036 998572
rect 436100 998520 436152 998572
rect 472440 998520 472492 998572
rect 500868 998520 500920 998572
rect 517520 998520 517572 998572
rect 557448 998520 557500 998572
rect 92388 998384 92440 998436
rect 100024 998384 100076 998436
rect 144000 998384 144052 998436
rect 155960 998384 156012 998436
rect 247500 998384 247552 998436
rect 200856 998316 200908 998368
rect 203524 998316 203576 998368
rect 246764 998248 246816 998300
rect 252468 998248 252520 998300
rect 200028 998180 200080 998232
rect 202696 998180 202748 998232
rect 250628 998112 250680 998164
rect 253664 998112 253716 998164
rect 197360 998044 197412 998096
rect 201868 998044 201920 998096
rect 202328 998044 202380 998096
rect 205548 998044 205600 998096
rect 92756 997976 92808 998028
rect 93492 997840 93544 997892
rect 94688 997840 94740 997892
rect 198004 997908 198056 997960
rect 200672 997908 200724 997960
rect 202144 997908 202196 997960
rect 204720 997908 204772 997960
rect 250444 997908 250496 997960
rect 253664 997908 253716 997960
rect 121736 997840 121788 997892
rect 195704 997772 195756 997824
rect 226340 997772 226392 997824
rect 247684 997772 247736 997824
rect 252468 997772 252520 997824
rect 355324 998384 355376 998436
rect 383476 998384 383528 998436
rect 431868 998384 431920 998436
rect 471796 998384 471848 998436
rect 497924 998384 497976 998436
rect 524052 998384 524104 998436
rect 555424 998384 555476 998436
rect 558828 998384 558880 998436
rect 572720 998384 572772 998436
rect 378600 998248 378652 998300
rect 382280 998248 382332 998300
rect 430028 998248 430080 998300
rect 432604 998248 432656 998300
rect 506296 998248 506348 998300
rect 517244 998248 517296 998300
rect 518164 998248 518216 998300
rect 523868 998248 523920 998300
rect 558000 998248 558052 998300
rect 560944 998248 560996 998300
rect 431224 998112 431276 998164
rect 433524 998112 433576 998164
rect 558828 998112 558880 998164
rect 562508 998112 562560 998164
rect 489276 998044 489328 998096
rect 493968 998044 494020 998096
rect 591304 998044 591356 998096
rect 625620 998044 625672 998096
rect 432052 997976 432104 998028
rect 436744 997976 436796 998028
rect 558000 997976 558052 998028
rect 560300 997976 560352 998028
rect 591120 997908 591172 997960
rect 625804 997908 625856 997960
rect 557632 997840 557684 997892
rect 559564 997840 559616 997892
rect 560024 997840 560076 997892
rect 562324 997840 562376 997892
rect 113824 997704 113876 997756
rect 117136 997704 117188 997756
rect 143816 997704 143868 997756
rect 160100 997704 160152 997756
rect 430028 997772 430080 997824
rect 432052 997772 432104 997824
rect 553952 997772 554004 997824
rect 555608 997772 555660 997824
rect 592040 997772 592092 997824
rect 625436 997772 625488 997824
rect 279240 997704 279292 997756
rect 298468 997704 298520 997756
rect 311900 997704 311952 997756
rect 355784 997704 355836 997756
rect 372344 997704 372396 997756
rect 433984 997704 434036 997756
rect 439688 997704 439740 997756
rect 489092 997704 489144 997756
rect 509240 997704 509292 997756
rect 509700 997704 509752 997756
rect 517060 997704 517112 997756
rect 558184 997704 558236 997756
rect 562692 997704 562744 997756
rect 566648 997704 566700 997756
rect 92572 997636 92624 997688
rect 101588 997636 101640 997688
rect 248052 997636 248104 997688
rect 259460 997636 259512 997688
rect 399944 997636 399996 997688
rect 432052 997636 432104 997688
rect 552664 997636 552716 997688
rect 109500 997568 109552 997620
rect 116124 997568 116176 997620
rect 144828 997568 144880 997620
rect 153936 997568 153988 997620
rect 299204 997568 299256 997620
rect 310520 997568 310572 997620
rect 365168 997568 365220 997620
rect 372528 997568 372580 997620
rect 432604 997568 432656 997620
rect 439872 997568 439924 997620
rect 488908 997568 488960 997620
rect 510804 997568 510856 997620
rect 618168 997636 618220 997688
rect 562140 997568 562192 997620
rect 246948 997500 247000 997552
rect 255964 997500 256016 997552
rect 540888 997500 540940 997552
rect 555424 997500 555476 997552
rect 508504 997432 508556 997484
rect 516692 997432 516744 997484
rect 571800 997568 571852 997620
rect 553308 997364 553360 997416
rect 562692 997432 562744 997484
rect 571616 997432 571668 997484
rect 571984 997432 572036 997484
rect 592040 997432 592092 997484
rect 562140 997296 562192 997348
rect 591304 997296 591356 997348
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 440240 997160 440292 997212
rect 445668 997160 445720 997212
rect 555608 997160 555660 997212
rect 570420 997160 570472 997212
rect 571800 997160 571852 997212
rect 590568 997160 590620 997212
rect 320824 997024 320876 997076
rect 332600 997024 332652 997076
rect 356060 997024 356112 997076
rect 372712 997024 372764 997076
rect 443644 997024 443696 997076
rect 453856 997024 453908 997076
rect 502984 997024 503036 997076
rect 516876 997024 516928 997076
rect 551928 997024 551980 997076
rect 623688 997024 623740 997076
rect 143724 996888 143776 996940
rect 151268 996888 151320 996940
rect 568488 996888 568540 996940
rect 571064 996888 571116 996940
rect 571616 996888 571668 996940
rect 572904 996888 572956 996940
rect 573364 996888 573416 996940
rect 591120 996888 591172 996940
rect 153016 996820 153068 996872
rect 158720 996820 158772 996872
rect 200212 996820 200264 996872
rect 203708 996820 203760 996872
rect 571248 996752 571300 996804
rect 590384 996752 590436 996804
rect 143816 996616 143868 996668
rect 149888 996616 149940 996668
rect 570604 996616 570656 996668
rect 144552 996480 144604 996532
rect 149060 996480 149112 996532
rect 590568 996412 590620 996464
rect 195244 996344 195296 996396
rect 198004 996344 198056 996396
rect 549444 996344 549496 996396
rect 550640 996344 550692 996396
rect 262864 996276 262916 996328
rect 270408 996276 270460 996328
rect 556160 996276 556212 996328
rect 590568 996208 590620 996260
rect 171784 996072 171836 996124
rect 211160 996072 211212 996124
rect 228364 996072 228416 996124
rect 263600 996072 263652 996124
rect 264244 996072 264296 996124
rect 299020 996072 299072 996124
rect 382924 996004 382976 996056
rect 169392 995936 169444 995988
rect 171692 995936 171744 995988
rect 213184 995936 213236 995988
rect 261116 995936 261168 995988
rect 269764 995936 269816 995988
rect 316040 995936 316092 995988
rect 354588 995936 354640 995988
rect 381544 995936 381596 995988
rect 433524 996072 433576 996124
rect 511264 996072 511316 996124
rect 563060 996072 563112 996124
rect 522304 995936 522356 995988
rect 560300 995936 560352 995988
rect 202972 995868 203024 995920
rect 205088 995868 205140 995920
rect 140780 995800 140832 995852
rect 144000 995800 144052 995852
rect 170680 995800 170732 995852
rect 171232 995800 171284 995852
rect 229744 995800 229796 995852
rect 262220 995800 262272 995852
rect 364984 995800 365036 995852
rect 400864 995800 400916 995852
rect 170864 995528 170916 995580
rect 246212 995528 246264 995580
rect 247132 995528 247184 995580
rect 297824 995528 297876 995580
rect 299388 995528 299440 995580
rect 380164 995528 380216 995580
rect 383108 995528 383160 995580
rect 383292 995528 383344 995580
rect 384764 995528 384816 995580
rect 385408 995528 385460 995580
rect 386972 995528 387024 995580
rect 472716 995528 472768 995580
rect 474004 995528 474056 995580
rect 493968 995528 494020 995580
rect 511080 995528 511132 995580
rect 524052 995528 524104 995580
rect 526076 995528 526128 995580
rect 625804 995528 625856 995580
rect 626540 995528 626592 995580
rect 194876 995460 194928 995512
rect 195520 995460 195572 995512
rect 475936 995460 475988 995512
rect 476396 995460 476448 995512
rect 476948 995460 477000 995512
rect 478972 995460 479024 995512
rect 211804 995392 211856 995444
rect 260932 995392 260984 995444
rect 171692 995277 171744 995329
rect 180708 995324 180760 995376
rect 202328 995324 202380 995376
rect 290648 995324 290700 995376
rect 296168 995256 296220 995308
rect 298652 995256 298704 995308
rect 171508 995165 171560 995217
rect 182962 995188 183014 995240
rect 208584 995188 208636 995240
rect 236230 995188 236282 995240
rect 251824 995188 251876 995240
rect 290832 995188 290884 995240
rect 295524 995188 295576 995240
rect 366364 995392 366416 995444
rect 402244 995392 402296 995444
rect 415400 995392 415452 995444
rect 402796 995324 402848 995376
rect 402980 995324 403032 995376
rect 362224 995256 362276 995308
rect 394608 995256 394660 995308
rect 307024 995188 307076 995240
rect 416136 995235 416188 995287
rect 171232 995053 171284 995105
rect 180156 995052 180208 995104
rect 206284 995052 206336 995104
rect 231584 995052 231636 995104
rect 257344 995052 257396 995104
rect 283472 995052 283524 995104
rect 305644 995052 305696 995104
rect 363604 994984 363656 995036
rect 384304 995120 384356 995172
rect 374368 994984 374420 995036
rect 392124 995120 392176 995172
rect 537760 995120 537812 995172
rect 538404 995120 538456 995172
rect 455880 995052 455932 995104
rect 487804 995052 487856 995104
rect 517704 995052 517756 995104
rect 533712 995052 533764 995104
rect 572720 995052 572772 995104
rect 635832 995052 635884 995104
rect 638868 995052 638920 995104
rect 640800 995052 640852 995104
rect 660304 995095 660356 995147
rect 384672 994984 384724 995036
rect 387800 994984 387852 995036
rect 387984 994984 388036 995036
rect 389364 994984 389416 995036
rect 389548 994984 389600 995036
rect 398840 994984 398892 995036
rect 183836 994916 183888 994968
rect 202144 994916 202196 994968
rect 232228 994916 232280 994968
rect 254584 994916 254636 994968
rect 284116 994916 284168 994968
rect 308404 994916 308456 994968
rect 420828 994916 420880 994968
rect 78312 994780 78364 994832
rect 104164 994780 104216 994832
rect 128452 994780 128504 994832
rect 157340 994780 157392 994832
rect 170496 994712 170548 994764
rect 171232 994829 171284 994881
rect 360844 994848 360896 994900
rect 402980 994848 403032 994900
rect 243268 994780 243320 994832
rect 246672 994780 246724 994832
rect 293224 994780 293276 994832
rect 298468 994780 298520 994832
rect 453856 994780 453908 994832
rect 489920 994780 489972 994832
rect 496728 994780 496780 994832
rect 538220 994780 538272 994832
rect 567844 994780 567896 994832
rect 639052 994780 639104 994832
rect 171048 994712 171100 994764
rect 243084 994712 243136 994764
rect 372712 994712 372764 994764
rect 393320 994712 393372 994764
rect 397644 994712 397696 994764
rect 402796 994712 402848 994764
rect 81348 994644 81400 994696
rect 98644 994644 98696 994696
rect 129096 994644 129148 994696
rect 142114 994644 142166 994696
rect 419448 994644 419500 994696
rect 660304 994644 660356 994696
rect 77668 994508 77720 994560
rect 93308 994508 93360 994560
rect 129740 994508 129792 994560
rect 134892 994508 134944 994560
rect 132408 994372 132460 994424
rect 149704 994576 149756 994628
rect 170864 994576 170916 994628
rect 300124 994576 300176 994628
rect 377404 994576 377456 994628
rect 397000 994576 397052 994628
rect 660764 994576 660816 994628
rect 472256 994508 472308 994560
rect 474924 994508 474976 994560
rect 481640 994508 481692 994560
rect 489736 994508 489788 994560
rect 499488 994508 499540 994560
rect 538588 994508 538640 994560
rect 571064 994508 571116 994560
rect 639512 994508 639564 994560
rect 660948 994508 661000 994560
rect 134892 994236 134944 994288
rect 153016 994440 153068 994492
rect 170680 994440 170732 994492
rect 250444 994440 250496 994492
rect 383108 994440 383160 994492
rect 389548 994440 389600 994492
rect 279240 994372 279292 994424
rect 316408 994372 316460 994424
rect 468484 994372 468536 994424
rect 484124 994372 484176 994424
rect 505744 994372 505796 994424
rect 149060 994304 149112 994356
rect 186136 994304 186188 994356
rect 186274 994304 186326 994356
rect 195796 994304 195848 994356
rect 226340 994236 226392 994288
rect 251456 994236 251508 994288
rect 294512 994236 294564 994288
rect 381176 994236 381228 994288
rect 414480 994236 414532 994288
rect 446128 994236 446180 994288
rect 471612 994236 471664 994288
rect 476304 994236 476356 994288
rect 519544 994372 519596 994424
rect 538404 994372 538456 994424
rect 572904 994372 572956 994424
rect 590568 994372 590620 994424
rect 625252 994372 625304 994424
rect 631508 994372 631560 994424
rect 528744 994236 528796 994288
rect 169392 994168 169444 994220
rect 142344 994100 142396 994152
rect 151084 994100 151136 994152
rect 298836 994100 298888 994152
rect 471796 994100 471848 994152
rect 475936 994100 475988 994152
rect 522120 994100 522172 994152
rect 539232 994236 539284 994288
rect 550640 994236 550692 994288
rect 572720 994236 572772 994288
rect 574100 994032 574152 994084
rect 141976 993964 142028 994016
rect 142344 993964 142396 994016
rect 181444 993964 181496 994016
rect 184296 993964 184348 994016
rect 184480 993964 184532 994016
rect 186136 993964 186188 994016
rect 186274 993964 186326 994016
rect 137560 993828 137612 993880
rect 141792 993828 141844 993880
rect 187608 993828 187660 993880
rect 190736 993828 190788 993880
rect 171232 993760 171284 993812
rect 187424 993760 187476 993812
rect 191104 993964 191156 994016
rect 203524 993964 203576 994016
rect 232872 993964 232924 994016
rect 258080 993964 258132 994016
rect 471980 993964 472032 994016
rect 477316 993964 477368 994016
rect 569224 993896 569276 993948
rect 207020 993828 207072 993880
rect 243084 993828 243136 993880
rect 247684 993828 247736 993880
rect 521292 993760 521344 993812
rect 660948 993760 661000 993812
rect 195934 993692 195986 993744
rect 196808 993692 196860 993744
rect 170496 993624 170548 993676
rect 190552 993488 190604 993540
rect 194876 993488 194928 993540
rect 197360 993624 197412 993676
rect 517244 993624 517296 993676
rect 660764 993624 660816 993676
rect 50344 993148 50396 993200
rect 107752 993148 107804 993200
rect 44824 993012 44876 993064
rect 109040 993012 109092 993064
rect 318064 993012 318116 993064
rect 349160 993012 349212 993064
rect 562508 993012 562560 993064
rect 660304 993012 660356 993064
rect 54484 992876 54536 992928
rect 148324 992876 148376 992928
rect 319444 992876 319496 992928
rect 364984 992876 365036 992928
rect 560944 992876 560996 992928
rect 667204 992876 667256 992928
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 51724 991584 51776 991636
rect 110420 991584 110472 991636
rect 138296 991584 138348 991636
rect 163136 991584 163188 991636
rect 369124 991584 369176 991636
rect 414112 991584 414164 991636
rect 55864 991448 55916 991500
rect 146944 991448 146996 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 367744 991448 367796 991500
rect 430304 991448 430356 991500
rect 435364 991448 435416 991500
rect 478972 991448 479024 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 214564 991176 214616 991228
rect 219440 991176 219492 991228
rect 164884 990836 164936 990888
rect 170772 990836 170824 990888
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 572720 990836 572772 990888
rect 576308 990836 576360 990888
rect 53288 990224 53340 990276
rect 95884 990224 95936 990276
rect 48964 990088 49016 990140
rect 108120 990088 108172 990140
rect 512644 990088 512696 990140
rect 543832 990088 543884 990140
rect 562324 990088 562376 990140
rect 668584 990088 668636 990140
rect 563704 987368 563756 987420
rect 608784 987368 608836 987420
rect 203156 986620 203208 986672
rect 204904 986620 204956 986672
rect 89628 986076 89680 986128
rect 111800 986076 111852 986128
rect 438124 986076 438176 986128
rect 462780 986076 462832 986128
rect 515404 986076 515456 986128
rect 527640 986076 527692 986128
rect 566464 986076 566516 986128
rect 592500 986076 592552 986128
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 370504 985940 370556 985992
rect 397828 985940 397880 985992
rect 436744 985940 436796 985992
rect 495164 985940 495216 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 664444 975672 664496 975724
rect 46204 961868 46256 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952348 36596 952400
rect 41696 952348 41748 952400
rect 33784 951464 33836 951516
rect 41512 951464 41564 951516
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 663064 948064 663116 948116
rect 676036 947996 676088 948048
rect 681004 947996 681056 948048
rect 45560 945956 45612 946008
rect 62120 945956 62172 946008
rect 28724 945276 28776 945328
rect 31760 945276 31812 945328
rect 35808 942556 35860 942608
rect 41696 942556 41748 942608
rect 35808 941196 35860 941248
rect 41696 941128 41748 941180
rect 35808 939768 35860 939820
rect 41512 939768 41564 939820
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 661684 921816 661736 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 663064 909440 663116 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 671344 895636 671396 895688
rect 44088 892712 44140 892764
rect 42938 892270 42990 892322
rect 43076 892202 43128 892254
rect 44088 891896 44140 891948
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 652392 855584 652444 855636
rect 664444 855584 664496 855636
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 35808 817028 35860 817080
rect 41696 817028 41748 817080
rect 35808 815600 35860 815652
rect 41604 815600 41656 815652
rect 651472 815600 651524 815652
rect 669964 815600 670016 815652
rect 35808 814240 35860 814292
rect 41420 814240 41472 814292
rect 41328 811588 41380 811640
rect 41696 811588 41748 811640
rect 40776 808936 40828 808988
rect 41604 808936 41656 808988
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 35164 802408 35216 802460
rect 41696 802408 41748 802460
rect 35900 802272 35952 802324
rect 41696 802272 41748 802324
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 651472 775548 651524 775600
rect 668768 775548 668820 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35808 768952 35860 769004
rect 41328 768952 41380 769004
rect 35624 768816 35676 768868
rect 41696 768816 41748 768868
rect 35440 768680 35492 768732
rect 40040 768680 40092 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35532 767320 35584 767372
rect 37924 767320 37976 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 37096 763240 37148 763292
rect 39304 763240 39356 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 37924 759024 37976 759076
rect 39488 759024 39540 759076
rect 35164 758412 35216 758464
rect 41696 758412 41748 758464
rect 42064 758344 42116 758396
rect 31024 758208 31076 758260
rect 40684 758140 40736 758192
rect 42064 758004 42116 758056
rect 39304 757596 39356 757648
rect 41696 757596 41748 757648
rect 676036 757120 676088 757172
rect 683120 757120 683172 757172
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 652576 735564 652628 735616
rect 671344 735564 671396 735616
rect 673552 732096 673604 732148
rect 674012 732096 674064 732148
rect 35808 730192 35860 730244
rect 41696 730192 41748 730244
rect 35624 730056 35676 730108
rect 41696 730056 41748 730108
rect 673828 728560 673880 728612
rect 673368 728424 673420 728476
rect 673000 728084 673052 728136
rect 674150 728084 674202 728136
rect 41328 725908 41380 725960
rect 41696 725908 41748 725960
rect 41328 724480 41380 724532
rect 41696 724480 41748 724532
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 31024 716796 31076 716848
rect 41604 716796 41656 716848
rect 33784 715640 33836 715692
rect 41512 715640 41564 715692
rect 33048 715504 33100 715556
rect 41696 715504 41748 715556
rect 36544 715368 36596 715420
rect 41604 715028 41656 715080
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 652576 709316 652628 709368
rect 664444 709316 664496 709368
rect 672448 707208 672500 707260
rect 673000 707208 673052 707260
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 652392 696940 652444 696992
rect 661684 696940 661736 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 35808 687216 35860 687268
rect 41696 687216 41748 687268
rect 35808 683136 35860 683188
rect 41512 683136 41564 683188
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35808 681708 35860 681760
rect 41328 681708 41380 681760
rect 35440 681028 35492 681080
rect 41604 681028 41656 681080
rect 35808 680620 35860 680672
rect 37924 680620 37976 680672
rect 35624 680348 35676 680400
rect 36544 680348 36596 680400
rect 51724 674840 51776 674892
rect 62120 674840 62172 674892
rect 35164 672732 35216 672784
rect 40500 672732 40552 672784
rect 36544 672052 36596 672104
rect 41604 672052 41656 672104
rect 39948 671440 40000 671492
rect 41696 671440 41748 671492
rect 651472 669332 651524 669384
rect 661868 669332 661920 669384
rect 671068 666204 671120 666256
rect 673368 666204 673420 666256
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651472 656888 651524 656940
rect 670148 656888 670200 656940
rect 54484 647844 54536 647896
rect 62120 647844 62172 647896
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639140 35860 639192
rect 41696 639072 41748 639124
rect 35808 638936 35860 638988
rect 40040 638936 40092 638988
rect 35808 637576 35860 637628
rect 41328 637576 41380 637628
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651472 629280 651524 629332
rect 667204 629280 667256 629332
rect 675852 626560 675904 626612
rect 676496 626560 676548 626612
rect 48964 623772 49016 623824
rect 62120 623772 62172 623824
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 43536 612892 43588 612944
rect 43371 612688 43423 612740
rect 43720 612484 43772 612536
rect 43582 612280 43634 612332
rect 46388 612348 46440 612400
rect 671896 612280 671948 612332
rect 671436 612144 671488 612196
rect 45560 611872 45612 611924
rect 46940 611668 46992 611720
rect 44042 611464 44094 611516
rect 45744 611260 45796 611312
rect 47216 611056 47268 611108
rect 44824 610920 44876 610972
rect 44379 610852 44431 610904
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 664628 603100 664680 603152
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 41236 594668 41288 594720
rect 41512 594668 41564 594720
rect 41328 593376 41380 593428
rect 41696 593376 41748 593428
rect 40500 592356 40552 592408
rect 41696 592356 41748 592408
rect 41052 592016 41104 592068
rect 41696 592016 41748 592068
rect 675944 591336 675996 591388
rect 679624 591336 679676 591388
rect 676128 591200 676180 591252
rect 682384 591200 682436 591252
rect 651472 590656 651524 590708
rect 662052 590656 662104 590708
rect 35164 585896 35216 585948
rect 41696 585896 41748 585948
rect 32404 585760 32456 585812
rect 41696 585760 41748 585812
rect 36544 585148 36596 585200
rect 41420 585148 41472 585200
rect 51724 583720 51776 583772
rect 62120 583720 62172 583772
rect 671068 578008 671120 578060
rect 671712 578008 671764 578060
rect 651472 576852 651524 576904
rect 666008 576852 666060 576904
rect 672264 571956 672316 572008
rect 672816 571956 672868 572008
rect 679624 571276 679676 571328
rect 683120 571276 683172 571328
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 35808 557540 35860 557592
rect 41512 557540 41564 557592
rect 35808 554752 35860 554804
rect 41696 554752 41748 554804
rect 35808 553528 35860 553580
rect 41696 553528 41748 553580
rect 35624 553392 35676 553444
rect 41328 553392 41380 553444
rect 41328 552032 41380 552084
rect 41604 552032 41656 552084
rect 41328 550740 41380 550792
rect 41604 550740 41656 550792
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 675852 547544 675904 547596
rect 678244 547544 678296 547596
rect 31760 547408 31812 547460
rect 37096 547408 37148 547460
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 33784 542988 33836 543040
rect 41512 542988 41564 543040
rect 37096 542308 37148 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669964 536800 670016 536852
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 672264 531972 672316 532024
rect 672632 531972 672684 532024
rect 673184 530408 673236 530460
rect 673828 530408 673880 530460
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 675852 518780 675904 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 675852 503616 675904 503668
rect 679624 503616 679676 503668
rect 676036 503480 676088 503532
rect 682384 503480 682436 503532
rect 675852 502324 675904 502376
rect 676864 502324 676916 502376
rect 676036 500896 676088 500948
rect 681004 500896 681056 500948
rect 652576 494708 652628 494760
rect 665824 494708 665876 494760
rect 676036 492668 676088 492720
rect 683396 492668 683448 492720
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 673368 488656 673420 488708
rect 673368 488248 673420 488300
rect 651472 484440 651524 484492
rect 668768 484372 668820 484424
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 651472 470568 651524 470620
rect 663064 470568 663116 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 652392 456764 652444 456816
rect 667204 456764 667256 456816
rect 673948 456152 674000 456204
rect 673828 456016 673880 456068
rect 673460 455812 673512 455864
rect 673598 455608 673650 455660
rect 673506 455336 673558 455388
rect 673388 455132 673440 455184
rect 671988 455064 672040 455116
rect 673164 454792 673216 454844
rect 673046 454588 673098 454640
rect 672954 454316 673006 454368
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672816 454044 672868 454096
rect 672264 453908 672316 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 671344 430584 671396 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 41328 423648 41380 423700
rect 41696 423648 41748 423700
rect 651840 416780 651892 416832
rect 661684 416780 661736 416832
rect 49148 415420 49200 415472
rect 62120 415420 62172 415472
rect 36544 415352 36596 415404
rect 41696 415352 41748 415404
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 41144 387064 41196 387116
rect 41696 387064 41748 387116
rect 41328 382372 41380 382424
rect 41512 382372 41564 382424
rect 35808 379652 35860 379704
rect 41696 379652 41748 379704
rect 40224 378496 40276 378548
rect 41696 378496 41748 378548
rect 35808 375368 35860 375420
rect 41696 375368 41748 375420
rect 51724 375368 51776 375420
rect 62120 375368 62172 375420
rect 37924 373260 37976 373312
rect 41696 373260 41748 373312
rect 651656 364352 651708 364404
rect 663248 364352 663300 364404
rect 46388 362924 46440 362976
rect 62120 362924 62172 362976
rect 45008 355784 45060 355836
rect 45652 355784 45704 355836
rect 44640 355648 44692 355700
rect 44575 354832 44627 354884
rect 44575 354628 44627 354680
rect 44799 354424 44851 354476
rect 44686 354288 44738 354340
rect 45652 354016 45704 354068
rect 45928 353744 45980 353796
rect 45560 353200 45612 353252
rect 651472 350548 651524 350600
rect 667388 350548 667440 350600
rect 28908 345040 28960 345092
rect 38292 345040 38344 345092
rect 35808 339464 35860 339516
rect 37924 339464 37976 339516
rect 35808 338104 35860 338156
rect 36544 338104 36596 338156
rect 651472 338104 651524 338156
rect 666192 338104 666244 338156
rect 50344 336744 50396 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 667756 324300 667808 324352
rect 54484 310496 54536 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667204 310496 667256 310548
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675944 298052 675996 298104
rect 678980 298052 679032 298104
rect 676128 297848 676180 297900
rect 681004 297848 681056 297900
rect 41328 285064 41380 285116
rect 41696 285064 41748 285116
rect 32404 284928 32456 284980
rect 41696 284928 41748 284980
rect 651472 284316 651524 284368
rect 667572 284316 667624 284368
rect 522948 276224 523000 276276
rect 526904 276224 526956 276276
rect 524880 276088 524932 276140
rect 88340 275952 88392 276004
rect 143356 275952 143408 276004
rect 156880 275952 156932 276004
rect 193864 275952 193916 276004
rect 201776 275952 201828 276004
rect 222108 275952 222160 276004
rect 389180 275952 389232 276004
rect 393320 275952 393372 276004
rect 400588 275952 400640 276004
rect 415768 275952 415820 276004
rect 427820 275952 427872 276004
rect 443000 275952 443052 276004
rect 443736 275952 443788 276004
rect 453580 275952 453632 276004
rect 456984 275952 457036 276004
rect 486700 275952 486752 276004
rect 486884 275952 486936 276004
rect 494704 275952 494756 276004
rect 495440 275952 495492 276004
rect 504364 275952 504416 276004
rect 504916 275952 504968 276004
rect 507032 275952 507084 276004
rect 508044 275952 508096 276004
rect 514024 275952 514076 276004
rect 95424 275816 95476 275868
rect 104808 275816 104860 275868
rect 113180 275816 113232 275868
rect 169944 275816 169996 275868
rect 181720 275816 181772 275868
rect 218888 275816 218940 275868
rect 393596 275816 393648 275868
rect 412272 275816 412324 275868
rect 415308 275816 415360 275868
rect 425244 275816 425296 275868
rect 432972 275816 433024 275868
rect 487896 275816 487948 275868
rect 498200 275816 498252 275868
rect 505652 275816 505704 275868
rect 507216 275816 507268 275868
rect 512736 275816 512788 275868
rect 512920 275816 512972 275868
rect 519820 275952 519872 276004
rect 520004 275952 520056 276004
rect 515496 275816 515548 275868
rect 81256 275680 81308 275732
rect 88984 275680 89036 275732
rect 103704 275680 103756 275732
rect 160100 275680 160152 275732
rect 178132 275680 178184 275732
rect 216864 275680 216916 275732
rect 299940 275680 299992 275732
rect 300768 275680 300820 275732
rect 370504 275680 370556 275732
rect 388628 275680 388680 275732
rect 410064 275680 410116 275732
rect 428832 275680 428884 275732
rect 429200 275680 429252 275732
rect 446496 275680 446548 275732
rect 76472 275544 76524 275596
rect 86868 275544 86920 275596
rect 96620 275544 96672 275596
rect 156604 275544 156656 275596
rect 163964 275544 164016 275596
rect 202144 275544 202196 275596
rect 221924 275544 221976 275596
rect 233884 275544 233936 275596
rect 236092 275544 236144 275596
rect 251088 275544 251140 275596
rect 350724 275544 350776 275596
rect 361396 275544 361448 275596
rect 362224 275544 362276 275596
rect 385040 275544 385092 275596
rect 388168 275544 388220 275596
rect 418160 275544 418212 275596
rect 418344 275544 418396 275596
rect 435916 275544 435968 275596
rect 445760 275544 445812 275596
rect 502064 275680 502116 275732
rect 502248 275680 502300 275732
rect 509148 275680 509200 275732
rect 512184 275680 512236 275732
rect 516232 275680 516284 275732
rect 516784 275816 516836 275868
rect 604920 275952 604972 276004
rect 524880 275816 524932 275868
rect 612004 275816 612056 275868
rect 519176 275680 519228 275732
rect 519360 275680 519412 275732
rect 449164 275544 449216 275596
rect 501788 275544 501840 275596
rect 85948 275408 86000 275460
rect 146668 275408 146720 275460
rect 160468 275408 160520 275460
rect 167736 275408 167788 275460
rect 171048 275408 171100 275460
rect 210792 275408 210844 275460
rect 218336 275408 218388 275460
rect 237472 275408 237524 275460
rect 244372 275408 244424 275460
rect 254584 275408 254636 275460
rect 260932 275408 260984 275460
rect 273536 275408 273588 275460
rect 273904 275408 273956 275460
rect 282920 275408 282972 275460
rect 326436 275408 326488 275460
rect 335360 275408 335412 275460
rect 341524 275408 341576 275460
rect 354312 275408 354364 275460
rect 298744 275340 298796 275392
rect 300032 275340 300084 275392
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 142712 275272 142764 275324
rect 183468 275272 183520 275324
rect 186412 275272 186464 275324
rect 187792 275272 187844 275324
rect 188804 275272 188856 275324
rect 222844 275272 222896 275324
rect 225420 275272 225472 275324
rect 245108 275272 245160 275324
rect 250260 275272 250312 275324
rect 266360 275272 266412 275324
rect 266820 275272 266872 275324
rect 276664 275272 276716 275324
rect 284576 275272 284628 275324
rect 290096 275272 290148 275324
rect 329472 275272 329524 275324
rect 338948 275272 339000 275324
rect 74080 275136 74132 275188
rect 77208 275136 77260 275188
rect 110788 275136 110840 275188
rect 162124 275136 162176 275188
rect 338948 275136 339000 275188
rect 353116 275272 353168 275324
rect 353944 275272 353996 275324
rect 360200 275408 360252 275460
rect 363052 275408 363104 275460
rect 367284 275408 367336 275460
rect 369124 275408 369176 275460
rect 377956 275408 378008 275460
rect 382004 275408 382056 275460
rect 414572 275408 414624 275460
rect 416412 275408 416464 275460
rect 463056 275408 463108 275460
rect 467656 275408 467708 275460
rect 519544 275544 519596 275596
rect 519728 275544 519780 275596
rect 522948 275544 523000 275596
rect 527364 275680 527416 275732
rect 619088 275680 619140 275732
rect 530492 275544 530544 275596
rect 530768 275544 530820 275596
rect 534908 275544 534960 275596
rect 538036 275544 538088 275596
rect 626172 275544 626224 275596
rect 504364 275408 504416 275460
rect 538220 275408 538272 275460
rect 356336 275272 356388 275324
rect 368480 275272 368532 275324
rect 375104 275272 375156 275324
rect 403992 275272 404044 275324
rect 411260 275272 411312 275324
rect 455972 275272 456024 275324
rect 456156 275272 456208 275324
rect 512184 275272 512236 275324
rect 420920 275136 420972 275188
rect 434720 275136 434772 275188
rect 437480 275136 437532 275188
rect 450084 275136 450136 275188
rect 456800 275136 456852 275188
rect 467840 275136 467892 275188
rect 468208 275136 468260 275188
rect 494520 275136 494572 275188
rect 494704 275136 494756 275188
rect 519360 275272 519412 275324
rect 519544 275272 519596 275324
rect 537576 275272 537628 275324
rect 537760 275272 537812 275324
rect 540980 275408 541032 275460
rect 541164 275408 541216 275460
rect 544292 275408 544344 275460
rect 544476 275408 544528 275460
rect 546040 275408 546092 275460
rect 546224 275408 546276 275460
rect 641628 275408 641680 275460
rect 538588 275272 538640 275324
rect 633348 275272 633400 275324
rect 224224 275068 224276 275120
rect 226156 275068 226208 275120
rect 294052 275068 294104 275120
rect 295156 275068 295208 275120
rect 135628 275000 135680 275052
rect 182088 275000 182140 275052
rect 449900 275000 449952 275052
rect 460664 275000 460716 275052
rect 488540 275000 488592 275052
rect 492588 275000 492640 275052
rect 494704 275000 494756 275052
rect 498568 275000 498620 275052
rect 505100 275000 505152 275052
rect 506848 275000 506900 275052
rect 507032 275000 507084 275052
rect 590752 275136 590804 275188
rect 611360 275136 611412 275188
rect 616788 275136 616840 275188
rect 619180 275136 619232 275188
rect 623872 275136 623924 275188
rect 514024 275000 514076 275052
rect 583668 275000 583720 275052
rect 71780 274932 71832 274984
rect 73804 274932 73856 274984
rect 277492 274932 277544 274984
rect 284300 274932 284352 274984
rect 129648 274864 129700 274916
rect 136548 274864 136600 274916
rect 149796 274864 149848 274916
rect 185584 274864 185636 274916
rect 289268 274864 289320 274916
rect 293408 274864 293460 274916
rect 471796 274864 471848 274916
rect 523132 274864 523184 274916
rect 523316 274864 523368 274916
rect 597836 274864 597888 274916
rect 283380 274796 283432 274848
rect 289084 274796 289136 274848
rect 404268 274796 404320 274848
rect 407488 274796 407540 274848
rect 426256 274796 426308 274848
rect 432328 274796 432380 274848
rect 106004 274728 106056 274780
rect 110420 274728 110472 274780
rect 140320 274728 140372 274780
rect 144644 274728 144696 274780
rect 146208 274728 146260 274780
rect 149888 274728 149940 274780
rect 435640 274728 435692 274780
rect 439412 274728 439464 274780
rect 453948 274728 454000 274780
rect 457168 274728 457220 274780
rect 464344 274728 464396 274780
rect 471336 274728 471388 274780
rect 482928 274728 482980 274780
rect 538680 274728 538732 274780
rect 539048 274728 539100 274780
rect 545856 274728 545908 274780
rect 546040 274728 546092 274780
rect 558828 274728 558880 274780
rect 570788 274728 570840 274780
rect 66996 274660 67048 274712
rect 71044 274660 71096 274712
rect 90640 274660 90692 274712
rect 95884 274660 95936 274712
rect 161572 274660 161624 274712
rect 163136 274660 163188 274712
rect 170128 274660 170180 274712
rect 173164 274660 173216 274712
rect 185216 274660 185268 274712
rect 187148 274660 187200 274712
rect 238484 274660 238536 274712
rect 239772 274660 239824 274712
rect 285772 274660 285824 274712
rect 286968 274660 287020 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 360292 274660 360344 274712
rect 363788 274660 363840 274712
rect 367100 274660 367152 274712
rect 369676 274660 369728 274712
rect 386052 274660 386104 274712
rect 389732 274660 389784 274712
rect 407120 274660 407172 274712
rect 411076 274660 411128 274712
rect 104808 274592 104860 274644
rect 157616 274592 157668 274644
rect 195888 274592 195940 274644
rect 206284 274592 206336 274644
rect 424968 274592 425020 274644
rect 474924 274592 474976 274644
rect 475384 274592 475436 274644
rect 538128 274592 538180 274644
rect 539048 274592 539100 274644
rect 570972 274592 571024 274644
rect 571800 274592 571852 274644
rect 121368 274456 121420 274508
rect 176752 274456 176804 274508
rect 182916 274456 182968 274508
rect 199660 274456 199712 274508
rect 210056 274456 210108 274508
rect 237840 274456 237892 274508
rect 392584 274456 392636 274508
rect 402796 274456 402848 274508
rect 406844 274456 406896 274508
rect 437480 274456 437532 274508
rect 440884 274456 440936 274508
rect 493784 274456 493836 274508
rect 496360 274456 496412 274508
rect 577780 274592 577832 274644
rect 585784 274456 585836 274508
rect 101312 274320 101364 274372
rect 160928 274320 160980 274372
rect 187792 274320 187844 274372
rect 220912 274320 220964 274372
rect 362868 274320 362920 274372
rect 386236 274320 386288 274372
rect 395896 274320 395948 274372
rect 420920 274320 420972 274372
rect 471244 274320 471296 274372
rect 491484 274320 491536 274372
rect 492496 274320 492548 274372
rect 570788 274320 570840 274372
rect 570972 274320 571024 274372
rect 586060 274320 586112 274372
rect 601424 274320 601476 274372
rect 84752 274184 84804 274236
rect 148324 274184 148376 274236
rect 160100 274184 160152 274236
rect 164240 274184 164292 274236
rect 176936 274184 176988 274236
rect 214656 274184 214708 274236
rect 220544 274184 220596 274236
rect 240600 274184 240652 274236
rect 342904 274184 342956 274236
rect 347228 274184 347280 274236
rect 366916 274184 366968 274236
rect 389180 274184 389232 274236
rect 390284 274184 390336 274236
rect 426440 274184 426492 274236
rect 438768 274184 438820 274236
rect 496176 274184 496228 274236
rect 501972 274184 502024 274236
rect 82360 274048 82412 274100
rect 145564 274048 145616 274100
rect 158076 274048 158128 274100
rect 200672 274048 200724 274100
rect 206560 274048 206612 274100
rect 235448 274048 235500 274100
rect 239588 274048 239640 274100
rect 258632 274048 258684 274100
rect 360108 274048 360160 274100
rect 383844 274048 383896 274100
rect 384948 274048 385000 274100
rect 419356 274048 419408 274100
rect 421564 274048 421616 274100
rect 458364 274048 458416 274100
rect 459376 274048 459428 274100
rect 516600 274048 516652 274100
rect 518440 274184 518492 274236
rect 602528 274184 602580 274236
rect 613384 274184 613436 274236
rect 615592 274184 615644 274236
rect 533896 274048 533948 274100
rect 534034 274048 534086 274100
rect 619180 274048 619232 274100
rect 77208 273912 77260 273964
rect 143540 273912 143592 273964
rect 145012 273912 145064 273964
rect 192484 273912 192536 273964
rect 193496 273912 193548 273964
rect 226340 273912 226392 273964
rect 234896 273912 234948 273964
rect 255504 273912 255556 273964
rect 256148 273912 256200 273964
rect 270592 273912 270644 273964
rect 271512 273912 271564 273964
rect 280804 273912 280856 273964
rect 346308 273912 346360 273964
rect 362592 273912 362644 273964
rect 377772 273912 377824 273964
rect 408684 273912 408736 273964
rect 413928 273912 413980 273964
rect 449900 273912 449952 273964
rect 451096 273912 451148 273964
rect 513840 273912 513892 273964
rect 517060 273912 517112 273964
rect 524236 273912 524288 273964
rect 524420 273912 524472 273964
rect 613200 273912 613252 273964
rect 123760 273776 123812 273828
rect 177488 273776 177540 273828
rect 426900 273776 426952 273828
rect 477224 273776 477276 273828
rect 491208 273776 491260 273828
rect 570604 273776 570656 273828
rect 280988 273708 281040 273760
rect 287520 273708 287572 273760
rect 134432 273640 134484 273692
rect 185032 273640 185084 273692
rect 460020 273640 460072 273692
rect 484308 273640 484360 273692
rect 487988 273640 488040 273692
rect 565912 273640 565964 273692
rect 570604 273640 570656 273692
rect 587164 273776 587216 273828
rect 144644 273504 144696 273556
rect 187792 273504 187844 273556
rect 429016 273504 429068 273556
rect 482008 273504 482060 273556
rect 487068 273504 487120 273556
rect 563520 273504 563572 273556
rect 481364 273368 481416 273420
rect 556436 273368 556488 273420
rect 347044 273232 347096 273284
rect 349620 273232 349672 273284
rect 350264 273232 350316 273284
rect 356336 273232 356388 273284
rect 409144 273232 409196 273284
rect 409880 273232 409932 273284
rect 114284 273164 114336 273216
rect 169024 273164 169076 273216
rect 104992 273028 105044 273080
rect 163320 273028 163372 273080
rect 167552 273028 167604 273080
rect 184204 273028 184256 273080
rect 187608 273028 187660 273080
rect 211988 273164 212040 273216
rect 419172 273164 419224 273216
rect 456800 273164 456852 273216
rect 463516 273164 463568 273216
rect 486884 273164 486936 273216
rect 493324 273164 493376 273216
rect 574192 273164 574244 273216
rect 578884 273164 578936 273216
rect 594340 273164 594392 273216
rect 211252 273028 211304 273080
rect 220084 273028 220136 273080
rect 382924 273028 382976 273080
rect 392124 273028 392176 273080
rect 403992 273028 404044 273080
rect 429200 273028 429252 273080
rect 434628 273028 434680 273080
rect 488724 273028 488776 273080
rect 496636 273028 496688 273080
rect 578516 273028 578568 273080
rect 580264 273028 580316 273080
rect 640432 273028 640484 273080
rect 78864 272892 78916 272944
rect 138664 272892 138716 272944
rect 141792 272892 141844 272944
rect 189816 272892 189868 272944
rect 191196 272892 191248 272944
rect 224868 272892 224920 272944
rect 288072 272892 288124 272944
rect 290464 272892 290516 272944
rect 373172 272892 373224 272944
rect 382648 272892 382700 272944
rect 94228 272756 94280 272808
rect 156052 272756 156104 272808
rect 180524 272756 180576 272808
rect 217232 272756 217284 272808
rect 228824 272756 228876 272808
rect 249064 272756 249116 272808
rect 352932 272756 352984 272808
rect 372988 272756 373040 272808
rect 380532 272756 380584 272808
rect 388628 272892 388680 272944
rect 391848 272892 391900 272944
rect 410064 272892 410116 272944
rect 412456 272892 412508 272944
rect 453948 272892 454000 272944
rect 458088 272892 458140 272944
rect 521844 272892 521896 272944
rect 87144 272620 87196 272672
rect 152004 272620 152056 272672
rect 168656 272620 168708 272672
rect 208492 272620 208544 272672
rect 217416 272620 217468 272672
rect 242164 272620 242216 272672
rect 242348 272620 242400 272672
rect 259552 272620 259604 272672
rect 331036 272620 331088 272672
rect 342444 272620 342496 272672
rect 368388 272620 368440 272672
rect 394516 272756 394568 272808
rect 397276 272756 397328 272808
rect 418344 272756 418396 272808
rect 426072 272756 426124 272808
rect 478420 272756 478472 272808
rect 482560 272756 482612 272808
rect 524374 272892 524426 272944
rect 524512 272892 524564 272944
rect 611360 272892 611412 272944
rect 388628 272620 388680 272672
rect 393596 272620 393648 272672
rect 393964 272620 394016 272672
rect 406292 272620 406344 272672
rect 408408 272620 408460 272672
rect 452476 272620 452528 272672
rect 453856 272620 453908 272672
rect 516416 272620 516468 272672
rect 516600 272620 516652 272672
rect 606116 272756 606168 272808
rect 524328 272620 524380 272672
rect 524512 272620 524564 272672
rect 524880 272620 524932 272672
rect 614396 272620 614448 272672
rect 77668 272484 77720 272536
rect 145104 272484 145156 272536
rect 152188 272484 152240 272536
rect 197544 272484 197596 272536
rect 199476 272484 199528 272536
rect 230572 272484 230624 272536
rect 231400 272484 231452 272536
rect 252744 272484 252796 272536
rect 252928 272484 252980 272536
rect 267740 272484 267792 272536
rect 268016 272484 268068 272536
rect 278780 272484 278832 272536
rect 279792 272484 279844 272536
rect 287152 272484 287204 272536
rect 338028 272484 338080 272536
rect 351920 272484 351972 272536
rect 358636 272484 358688 272536
rect 380348 272484 380400 272536
rect 380716 272484 380768 272536
rect 413376 272484 413428 272536
rect 415124 272484 415176 272536
rect 461860 272484 461912 272536
rect 463332 272484 463384 272536
rect 524512 272484 524564 272536
rect 524696 272484 524748 272536
rect 533988 272484 534040 272536
rect 534172 272484 534224 272536
rect 632152 272484 632204 272536
rect 127348 272348 127400 272400
rect 179880 272348 179932 272400
rect 439320 272348 439372 272400
rect 473728 272348 473780 272400
rect 474648 272348 474700 272400
rect 495440 272348 495492 272400
rect 501604 272348 501656 272400
rect 581276 272348 581328 272400
rect 139124 272212 139176 272264
rect 141424 272212 141476 272264
rect 143908 272212 143960 272264
rect 190736 272212 190788 272264
rect 451924 272212 451976 272264
rect 480812 272212 480864 272264
rect 488356 272212 488408 272264
rect 567108 272212 567160 272264
rect 153292 272076 153344 272128
rect 171784 272076 171836 272128
rect 473084 272076 473136 272128
rect 482928 272076 482980 272128
rect 483388 272076 483440 272128
rect 560024 272076 560076 272128
rect 478420 271940 478472 271992
rect 552480 271940 552532 271992
rect 552848 271940 552900 271992
rect 580080 271940 580132 271992
rect 110420 271804 110472 271856
rect 164976 271804 165028 271856
rect 175832 271804 175884 271856
rect 207664 271804 207716 271856
rect 214840 271804 214892 271856
rect 221464 271804 221516 271856
rect 222108 271804 222160 271856
rect 232136 271804 232188 271856
rect 356520 271804 356572 271856
rect 359004 271804 359056 271856
rect 394332 271804 394384 271856
rect 426256 271804 426308 271856
rect 427084 271804 427136 271856
rect 433524 271804 433576 271856
rect 447784 271804 447836 271856
rect 504548 271804 504600 271856
rect 504732 271804 504784 271856
rect 589556 271804 589608 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 93032 271668 93084 271720
rect 120724 271668 120776 271720
rect 120908 271668 120960 271720
rect 175280 271668 175332 271720
rect 192300 271668 192352 271720
rect 225512 271668 225564 271720
rect 237472 271668 237524 271720
rect 243728 271668 243780 271720
rect 355324 271668 355376 271720
rect 374368 271668 374420 271720
rect 387708 271668 387760 271720
rect 421380 271668 421432 271720
rect 421748 271668 421800 271720
rect 438216 271668 438268 271720
rect 442908 271668 442960 271720
rect 500500 271668 500552 271720
rect 500868 271668 500920 271720
rect 508044 271668 508096 271720
rect 508964 271668 509016 271720
rect 596640 271804 596692 271856
rect 591488 271668 591540 271720
rect 603724 271668 603776 271720
rect 111984 271532 112036 271584
rect 168380 271532 168432 271584
rect 173440 271532 173492 271584
rect 212632 271532 212684 271584
rect 226156 271532 226208 271584
rect 247224 271532 247276 271584
rect 259736 271532 259788 271584
rect 272616 271532 272668 271584
rect 372528 271532 372580 271584
rect 400404 271532 400456 271584
rect 409788 271532 409840 271584
rect 443736 271532 443788 271584
rect 453304 271532 453356 271584
rect 511540 271532 511592 271584
rect 511908 271532 511960 271584
rect 600228 271532 600280 271584
rect 607864 271532 607916 271584
rect 643928 271532 643980 271584
rect 89720 271396 89772 271448
rect 152648 271396 152700 271448
rect 165160 271396 165212 271448
rect 205732 271396 205784 271448
rect 223580 271396 223632 271448
rect 247408 271396 247460 271448
rect 247868 271396 247920 271448
rect 264336 271396 264388 271448
rect 334624 271396 334676 271448
rect 341340 271396 341392 271448
rect 342168 271396 342220 271448
rect 356704 271396 356756 271448
rect 360844 271396 360896 271448
rect 381544 271396 381596 271448
rect 397920 271396 397972 271448
rect 427084 271396 427136 271448
rect 427268 271396 427320 271448
rect 72976 271260 73028 271312
rect 142160 271260 142212 271312
rect 150992 271260 151044 271312
rect 195980 271260 196032 271312
rect 215944 271260 215996 271312
rect 242072 271260 242124 271312
rect 243176 271260 243228 271312
rect 261024 271260 261076 271312
rect 275100 271260 275152 271312
rect 283472 271260 283524 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 325516 271260 325568 271312
rect 334164 271260 334216 271312
rect 340604 271260 340656 271312
rect 355508 271260 355560 271312
rect 364156 271260 364208 271312
rect 386052 271260 386104 271312
rect 400128 271260 400180 271312
rect 435640 271260 435692 271312
rect 436928 271396 436980 271448
rect 454776 271396 454828 271448
rect 457444 271396 457496 271448
rect 511724 271396 511776 271448
rect 448888 271260 448940 271312
rect 454684 271260 454736 271312
rect 515128 271396 515180 271448
rect 515312 271396 515364 271448
rect 518624 271396 518676 271448
rect 520096 271396 520148 271448
rect 523960 271396 524012 271448
rect 524144 271396 524196 271448
rect 514484 271260 514536 271312
rect 529020 271260 529072 271312
rect 529388 271396 529440 271448
rect 610808 271396 610860 271448
rect 617984 271260 618036 271312
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 208860 271124 208912 271176
rect 237472 271124 237524 271176
rect 240784 271124 240836 271176
rect 259828 271124 259880 271176
rect 262128 271124 262180 271176
rect 274640 271124 274692 271176
rect 276296 271124 276348 271176
rect 284484 271124 284536 271176
rect 333888 271124 333940 271176
rect 344468 271124 344520 271176
rect 344652 271124 344704 271176
rect 350724 271124 350776 271176
rect 351828 271124 351880 271176
rect 372068 271124 372120 271176
rect 379428 271124 379480 271176
rect 407120 271124 407172 271176
rect 416596 271124 416648 271176
rect 463976 271124 464028 271176
rect 464528 271124 464580 271176
rect 524512 271124 524564 271176
rect 524696 271124 524748 271176
rect 529388 271124 529440 271176
rect 529572 271124 529624 271176
rect 532792 271124 532844 271176
rect 533160 271124 533212 271176
rect 621480 271124 621532 271176
rect 621664 271124 621716 271176
rect 636844 271124 636896 271176
rect 128544 270988 128596 271040
rect 181352 270988 181404 271040
rect 190000 270988 190052 271040
rect 216128 270988 216180 271040
rect 381544 270988 381596 271040
rect 399208 270988 399260 271040
rect 401324 270988 401376 271040
rect 130844 270852 130896 270904
rect 182456 270852 182508 270904
rect 200488 270852 200540 270904
rect 224224 270852 224276 270904
rect 389088 270852 389140 270904
rect 415308 270852 415360 270904
rect 425704 270988 425756 271040
rect 427268 270988 427320 271040
rect 431684 270988 431736 271040
rect 485504 270988 485556 271040
rect 488724 270988 488776 271040
rect 551744 270988 551796 271040
rect 552664 270988 552716 271040
rect 591488 270988 591540 271040
rect 427820 270852 427872 270904
rect 435364 270852 435416 270904
rect 436928 270852 436980 270904
rect 445024 270852 445076 270904
rect 497372 270852 497424 270904
rect 507676 270852 507728 270904
rect 522028 270852 522080 270904
rect 524788 270852 524840 270904
rect 593144 270852 593196 270904
rect 137928 270716 137980 270768
rect 187884 270716 187936 270768
rect 433156 270716 433208 270768
rect 456984 270716 457036 270768
rect 465724 270716 465776 270768
rect 526260 270716 526312 270768
rect 526444 270716 526496 270768
rect 528652 270716 528704 270768
rect 529020 270716 529072 270768
rect 116676 270580 116728 270632
rect 151084 270580 151136 270632
rect 237288 270580 237340 270632
rect 115848 270444 115900 270496
rect 171232 270444 171284 270496
rect 173164 270444 173216 270496
rect 210148 270444 210200 270496
rect 210792 270444 210844 270496
rect 211804 270444 211856 270496
rect 233148 270444 233200 270496
rect 237288 270444 237340 270496
rect 428464 270580 428516 270632
rect 466644 270580 466696 270632
rect 477500 270580 477552 270632
rect 538864 270580 538916 270632
rect 540520 270716 540572 270768
rect 543556 270716 543608 270768
rect 543694 270716 543746 270768
rect 607312 270716 607364 270768
rect 552664 270580 552716 270632
rect 252008 270444 252060 270496
rect 292856 270444 292908 270496
rect 296260 270444 296312 270496
rect 359740 270444 359792 270496
rect 376760 270444 376812 270496
rect 377588 270444 377640 270496
rect 394700 270444 394752 270496
rect 397092 270444 397144 270496
rect 423680 270444 423732 270496
rect 424600 270444 424652 270496
rect 476304 270444 476356 270496
rect 479248 270444 479300 270496
rect 552204 270444 552256 270496
rect 552388 270444 552440 270496
rect 564440 270444 564492 270496
rect 110236 270308 110288 270360
rect 167920 270308 167972 270360
rect 172428 270308 172480 270360
rect 208676 270308 208728 270360
rect 212448 270308 212500 270360
rect 239956 270308 240008 270360
rect 253848 270308 253900 270360
rect 265072 270308 265124 270360
rect 291660 270308 291712 270360
rect 295524 270308 295576 270360
rect 348424 270308 348476 270360
rect 363052 270308 363104 270360
rect 364984 270308 365036 270360
rect 390560 270308 390612 270360
rect 392308 270308 392360 270360
rect 429384 270308 429436 270360
rect 429568 270308 429620 270360
rect 483112 270308 483164 270360
rect 486700 270308 486752 270360
rect 490380 270308 490432 270360
rect 490564 270308 490616 270360
rect 560300 270308 560352 270360
rect 316960 270240 317012 270292
rect 321560 270240 321612 270292
rect 339316 270240 339368 270292
rect 341524 270240 341576 270292
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 166908 270172 166960 270224
rect 207388 270172 207440 270224
rect 213828 270172 213880 270224
rect 240508 270172 240560 270224
rect 249616 270172 249668 270224
rect 263324 270172 263376 270224
rect 269212 270172 269264 270224
rect 279700 270172 279752 270224
rect 321928 270172 321980 270224
rect 328460 270172 328512 270224
rect 341800 270172 341852 270224
rect 357440 270172 357492 270224
rect 369400 270172 369452 270224
rect 396080 270172 396132 270224
rect 403072 270172 403124 270224
rect 444380 270172 444432 270224
rect 446956 270172 447008 270224
rect 504180 270172 504232 270224
rect 504364 270172 504416 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 528928 270172 528980 270224
rect 533528 270172 533580 270224
rect 533988 270172 534040 270224
rect 626540 270172 626592 270224
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 146668 270036 146720 270088
rect 151360 270036 151412 270088
rect 75828 269900 75880 269952
rect 142620 269900 142672 269952
rect 143356 269900 143408 269952
rect 153844 270036 153896 270088
rect 159916 270036 159968 270088
rect 202696 270036 202748 270088
rect 205548 270036 205600 270088
rect 234988 270036 235040 270088
rect 239772 270036 239824 270088
rect 253204 270036 253256 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 323584 270036 323636 270088
rect 331220 270036 331272 270088
rect 354220 270036 354272 270088
rect 375380 270036 375432 270088
rect 376576 270036 376628 270088
rect 404268 270036 404320 270088
rect 417148 270036 417200 270088
rect 465080 270036 465132 270088
rect 466000 270036 466052 270088
rect 528468 270036 528520 270088
rect 538864 270036 538916 270088
rect 540980 270036 541032 270088
rect 541808 270036 541860 270088
rect 541992 270036 542044 270088
rect 633624 270036 633676 270088
rect 154488 269900 154540 269952
rect 198188 269900 198240 269952
rect 198648 269900 198700 269952
rect 230020 269900 230072 269952
rect 230388 269900 230440 269952
rect 252376 269900 252428 269952
rect 258448 269900 258500 269952
rect 272248 269900 272300 269952
rect 273076 269900 273128 269952
rect 282184 269900 282236 269952
rect 286784 269900 286836 269952
rect 292120 269900 292172 269952
rect 331680 269900 331732 269952
rect 336740 269900 336792 269952
rect 347596 269900 347648 269952
rect 365720 269900 365772 269952
rect 372344 269900 372396 269952
rect 401784 269900 401836 269952
rect 413008 269900 413060 269952
rect 459560 269900 459612 269952
rect 461860 269900 461912 269952
rect 528652 269900 528704 269952
rect 529756 269900 529808 269952
rect 530768 269900 530820 269952
rect 530952 269900 531004 269952
rect 532976 269900 533028 269952
rect 536564 269900 536616 269952
rect 630680 269900 630732 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 139952 269764 140004 269816
rect 181168 269764 181220 269816
rect 182088 269764 182140 269816
rect 186964 269764 187016 269816
rect 187332 269764 187384 269816
rect 191932 269764 191984 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 84108 269628 84160 269680
rect 119804 269628 119856 269680
rect 119068 269492 119120 269544
rect 173716 269628 173768 269680
rect 184756 269628 184808 269680
rect 213828 269628 213880 269680
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 251456 269764 251508 269816
rect 267280 269764 267332 269816
rect 270316 269764 270368 269816
rect 280528 269764 280580 269816
rect 314476 269764 314528 269816
rect 318800 269764 318852 269816
rect 326896 269764 326948 269816
rect 335912 269764 335964 269816
rect 336832 269764 336884 269816
rect 350540 269764 350592 269816
rect 356704 269764 356756 269816
rect 378140 269764 378192 269816
rect 385684 269764 385736 269816
rect 419540 269764 419592 269816
rect 420000 269764 420052 269816
rect 468024 269764 468076 269816
rect 470968 269764 471020 269816
rect 537484 269764 537536 269816
rect 538864 269764 538916 269816
rect 552296 269764 552348 269816
rect 552480 269764 552532 269816
rect 641904 269764 641956 269816
rect 253204 269628 253256 269680
rect 258172 269628 258224 269680
rect 329656 269628 329708 269680
rect 339500 269628 339552 269680
rect 351644 269628 351696 269680
rect 364340 269628 364392 269680
rect 384028 269628 384080 269680
rect 388168 269628 388220 269680
rect 394700 269628 394752 269680
rect 416780 269628 416832 269680
rect 427360 269628 427412 269680
rect 478880 269628 478932 269680
rect 484216 269628 484268 269680
rect 490564 269628 490616 269680
rect 490748 269628 490800 269680
rect 504364 269628 504416 269680
rect 504548 269628 504600 269680
rect 553032 269628 553084 269680
rect 558920 269628 558972 269680
rect 572720 269628 572772 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 187332 269492 187384 269544
rect 208308 269492 208360 269544
rect 230756 269492 230808 269544
rect 401600 269492 401652 269544
rect 430580 269492 430632 269544
rect 449900 269492 449952 269544
rect 471980 269492 472032 269544
rect 474280 269492 474332 269544
rect 118608 269356 118660 269408
rect 166908 269356 166960 269408
rect 335636 269356 335688 269408
rect 343824 269356 343876 269408
rect 404360 269356 404412 269408
rect 426624 269356 426676 269408
rect 457720 269356 457772 269408
rect 471796 269356 471848 269408
rect 476764 269356 476816 269408
rect 537484 269492 537536 269544
rect 540980 269492 541032 269544
rect 541348 269492 541400 269544
rect 552388 269492 552440 269544
rect 568580 269492 568632 269544
rect 136824 269220 136876 269272
rect 182180 269220 182232 269272
rect 264888 269220 264940 269272
rect 269120 269220 269172 269272
rect 321100 269220 321152 269272
rect 327908 269220 327960 269272
rect 468760 269220 468812 269272
rect 537024 269220 537076 269272
rect 546224 269356 546276 269408
rect 546408 269356 546460 269408
rect 551928 269356 551980 269408
rect 549444 269220 549496 269272
rect 549628 269220 549680 269272
rect 553032 269356 553084 269408
rect 557540 269356 557592 269408
rect 552296 269220 552348 269272
rect 607588 269220 607640 269272
rect 282736 269084 282788 269136
rect 288808 269084 288860 269136
rect 295340 269084 295392 269136
rect 297548 269084 297600 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 434444 269084 434496 269136
rect 489920 269084 489972 269136
rect 108948 269016 109000 269068
rect 166264 269016 166316 269068
rect 185584 269016 185636 269068
rect 196900 269016 196952 269068
rect 251088 269016 251140 269068
rect 256516 269016 256568 269068
rect 86868 268880 86920 268932
rect 144736 268880 144788 268932
rect 179328 268880 179380 268932
rect 215944 268880 215996 268932
rect 382372 268880 382424 268932
rect 400588 268880 400640 268932
rect 102508 268744 102560 268796
rect 162952 268744 163004 268796
rect 163136 268744 163188 268796
rect 203524 268744 203576 268796
rect 203984 268744 204036 268796
rect 227720 268744 227772 268796
rect 227904 268744 227956 268796
rect 250720 268744 250772 268796
rect 387340 268744 387392 268796
rect 422300 269016 422352 269068
rect 503260 269016 503312 269068
rect 581460 269016 581512 269068
rect 581644 269016 581696 269068
rect 584128 269016 584180 269068
rect 590660 269016 590712 269068
rect 418988 268880 419040 268932
rect 440240 268880 440292 268932
rect 443644 268880 443696 268932
rect 502432 268880 502484 268932
rect 503444 268880 503496 268932
rect 505100 268880 505152 268932
rect 508504 268880 508556 268932
rect 594800 268880 594852 268932
rect 422300 268744 422352 268796
rect 436100 268744 436152 268796
rect 441160 268744 441212 268796
rect 499580 268744 499632 268796
rect 500684 268744 500736 268796
rect 581276 268744 581328 268796
rect 581644 268744 581696 268796
rect 598848 268744 598900 268796
rect 99288 268608 99340 268660
rect 160468 268608 160520 268660
rect 162768 268608 162820 268660
rect 205180 268608 205232 268660
rect 219532 268608 219584 268660
rect 244924 268608 244976 268660
rect 363052 268608 363104 268660
rect 386420 268608 386472 268660
rect 400588 268608 400640 268660
rect 441620 268608 441672 268660
rect 442724 268608 442776 268660
rect 445760 268608 445812 268660
rect 446588 268608 446640 268660
rect 503444 268608 503496 268660
rect 504180 268608 504232 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 155868 268472 155920 268524
rect 200212 268472 200264 268524
rect 202972 268472 203024 268524
rect 233332 268472 233384 268524
rect 245568 268472 245620 268524
rect 263140 268472 263192 268524
rect 263508 268472 263560 268524
rect 275560 268472 275612 268524
rect 333520 268472 333572 268524
rect 345112 268472 345164 268524
rect 345940 268472 345992 268524
rect 360292 268472 360344 268524
rect 361028 268472 361080 268524
rect 369860 268472 369912 268524
rect 370320 268472 370372 268524
rect 397460 268472 397512 268524
rect 402244 268472 402296 268524
rect 443276 268472 443328 268524
rect 448612 268472 448664 268524
rect 504364 268472 504416 268524
rect 506112 268608 506164 268660
rect 514024 268608 514076 268660
rect 514208 268608 514260 268660
rect 590660 268608 590712 268660
rect 608692 268608 608744 268660
rect 66260 268336 66312 268388
rect 137284 268336 137336 268388
rect 147588 268336 147640 268388
rect 193588 268336 193640 268388
rect 197268 268336 197320 268388
rect 229192 268336 229244 268388
rect 233700 268336 233752 268388
rect 254860 268336 254912 268388
rect 255320 268336 255372 268388
rect 269764 268336 269816 268388
rect 322756 268336 322808 268388
rect 329840 268336 329892 268388
rect 335176 268336 335228 268388
rect 347780 268336 347832 268388
rect 350080 268336 350132 268388
rect 367100 268336 367152 268388
rect 374920 268336 374972 268388
rect 404544 268336 404596 268388
rect 407212 268336 407264 268388
rect 451464 268336 451516 268388
rect 461032 268336 461084 268388
rect 518900 268336 518952 268388
rect 519360 268472 519412 268524
rect 533896 268472 533948 268524
rect 534034 268472 534086 268524
rect 619640 268472 619692 268524
rect 520280 268336 520332 268388
rect 520464 268336 520516 268388
rect 526996 268336 527048 268388
rect 527180 268336 527232 268388
rect 547512 268336 547564 268388
rect 547696 268336 547748 268388
rect 638960 268336 639012 268388
rect 122748 268200 122800 268252
rect 176200 268200 176252 268252
rect 436192 268200 436244 268252
rect 480996 268200 481048 268252
rect 504180 268200 504232 268252
rect 504364 268200 504416 268252
rect 509608 268200 509660 268252
rect 510712 268200 510764 268252
rect 513840 268200 513892 268252
rect 514024 268200 514076 268252
rect 591028 268200 591080 268252
rect 133788 268064 133840 268116
rect 183652 268064 183704 268116
rect 420460 268064 420512 268116
rect 469036 268064 469088 268116
rect 469220 268064 469272 268116
rect 480444 268064 480496 268116
rect 488540 268064 488592 268116
rect 491484 268064 491536 268116
rect 494704 268064 494756 268116
rect 499120 268064 499172 268116
rect 579620 268064 579672 268116
rect 581460 268064 581512 268116
rect 587900 268064 587952 268116
rect 125508 267928 125560 267980
rect 147588 267928 147640 267980
rect 437848 267928 437900 267980
rect 468208 267928 468260 267980
rect 431960 267792 432012 267844
rect 447140 267792 447192 267844
rect 533896 267928 533948 267980
rect 534034 267928 534086 267980
rect 581644 267928 581696 267980
rect 95884 267656 95936 267708
rect 154672 267656 154724 267708
rect 162124 267656 162176 267708
rect 169576 267656 169628 267708
rect 171784 267656 171836 267708
rect 199384 267656 199436 267708
rect 207664 267656 207716 267708
rect 213460 267656 213512 267708
rect 216128 267656 216180 267708
rect 223396 267656 223448 267708
rect 368204 267656 368256 267708
rect 377588 267656 377640 267708
rect 388168 267656 388220 267708
rect 397092 267656 397144 267708
rect 398104 267656 398156 267708
rect 421748 267656 421800 267708
rect 430396 267656 430448 267708
rect 460020 267656 460072 267708
rect 460204 267656 460256 267708
rect 465540 267656 465592 267708
rect 466828 267656 466880 267708
rect 489184 267792 489236 267844
rect 567660 267792 567712 267844
rect 579620 267792 579672 267844
rect 582380 267792 582432 267844
rect 470140 267656 470192 267708
rect 518808 267656 518860 267708
rect 518992 267656 519044 267708
rect 533988 267656 534040 267708
rect 534172 267656 534224 267708
rect 537024 267656 537076 267708
rect 537208 267656 537260 267708
rect 539048 267656 539100 267708
rect 539692 267656 539744 267708
rect 543556 267656 543608 267708
rect 543694 267656 543746 267708
rect 546408 267656 546460 267708
rect 546592 267656 546644 267708
rect 580264 267656 580316 267708
rect 88984 267520 89036 267572
rect 144552 267520 144604 267572
rect 144920 267520 144972 267572
rect 150532 267520 150584 267572
rect 151084 267520 151136 267572
rect 172888 267520 172940 267572
rect 187148 267520 187200 267572
rect 221740 267520 221792 267572
rect 227720 267520 227772 267572
rect 234160 267520 234212 267572
rect 313648 267520 313700 267572
rect 317788 267520 317840 267572
rect 370780 267520 370832 267572
rect 381544 267520 381596 267572
rect 383200 267520 383252 267572
rect 394700 267520 394752 267572
rect 397092 267520 397144 267572
rect 422300 267520 422352 267572
rect 443460 267520 443512 267572
rect 449900 267520 449952 267572
rect 450084 267520 450136 267572
rect 481548 267520 481600 267572
rect 481732 267520 481784 267572
rect 503076 267520 503128 267572
rect 504180 267520 504232 267572
rect 107568 267384 107620 267436
rect 167092 267384 167144 267436
rect 167736 267384 167788 267436
rect 204352 267384 204404 267436
rect 211988 267384 212040 267436
rect 222568 267384 222620 267436
rect 224224 267384 224276 267436
rect 231676 267384 231728 267436
rect 233884 267384 233936 267436
rect 246580 267384 246632 267436
rect 334348 267384 334400 267436
rect 342904 267384 342956 267436
rect 350908 267384 350960 267436
rect 361028 267384 361080 267436
rect 365812 267384 365864 267436
rect 382924 267384 382976 267436
rect 390652 267384 390704 267436
rect 404360 267384 404412 267436
rect 409604 267384 409656 267436
rect 435364 267384 435416 267436
rect 440332 267384 440384 267436
rect 485734 267384 485786 267436
rect 485872 267384 485924 267436
rect 487068 267384 487120 267436
rect 487252 267384 487304 267436
rect 491484 267384 491536 267436
rect 491668 267384 491720 267436
rect 492496 267384 492548 267436
rect 492680 267384 492732 267436
rect 504364 267384 504416 267436
rect 506480 267520 506532 267572
rect 507216 267520 507268 267572
rect 507400 267520 507452 267572
rect 578884 267520 578936 267572
rect 552848 267384 552900 267436
rect 100668 267248 100720 267300
rect 159824 267248 159876 267300
rect 166908 267248 166960 267300
rect 174544 267248 174596 267300
rect 175096 267248 175148 267300
rect 214288 267248 214340 267300
rect 220084 267248 220136 267300
rect 239128 267248 239180 267300
rect 254584 267248 254636 267300
rect 262312 267248 262364 267300
rect 312820 267248 312872 267300
rect 316040 267248 316092 267300
rect 343456 267248 343508 267300
rect 353944 267248 353996 267300
rect 363328 267248 363380 267300
rect 370504 267248 370556 267300
rect 375748 267248 375800 267300
rect 393964 267248 394016 267300
rect 399760 267248 399812 267300
rect 418988 267248 419040 267300
rect 421288 267248 421340 267300
rect 464344 267248 464396 267300
rect 465172 267248 465224 267300
rect 480904 267248 480956 267300
rect 481088 267248 481140 267300
rect 518808 267248 518860 267300
rect 518992 267248 519044 267300
rect 533896 267248 533948 267300
rect 534034 267248 534086 267300
rect 538864 267248 538916 267300
rect 539048 267248 539100 267300
rect 621664 267248 621716 267300
rect 71044 267112 71096 267164
rect 138112 267112 138164 267164
rect 141424 267112 141476 267164
rect 73804 266976 73856 267028
rect 141424 266976 141476 267028
rect 144552 267112 144604 267164
rect 147404 267112 147456 267164
rect 147588 267112 147640 267164
rect 149060 267112 149112 267164
rect 149888 267112 149940 267164
rect 194416 267112 194468 267164
rect 199660 267112 199712 267164
rect 218428 267112 218480 267164
rect 221464 267112 221516 267164
rect 241612 267112 241664 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 336004 267112 336056 267164
rect 347044 267112 347096 267164
rect 355876 267112 355928 267164
rect 369124 267112 369176 267164
rect 373264 267112 373316 267164
rect 392584 267112 392636 267164
rect 404728 267112 404780 267164
rect 431960 267112 432012 267164
rect 439504 267112 439556 267164
rect 445024 267112 445076 267164
rect 445300 267112 445352 267164
rect 450084 267112 450136 267164
rect 450268 267112 450320 267164
rect 499580 267112 499632 267164
rect 499764 267112 499816 267164
rect 504180 267112 504232 267164
rect 504364 267112 504416 267164
rect 521752 267112 521804 267164
rect 184020 266976 184072 267028
rect 184204 266976 184256 267028
rect 132408 266840 132460 266892
rect 184480 266840 184532 266892
rect 193864 266976 193916 267028
rect 201868 266976 201920 267028
rect 206284 266976 206336 267028
rect 228364 266976 228416 267028
rect 237288 266976 237340 267028
rect 254032 266976 254084 267028
rect 271420 266976 271472 267028
rect 276664 266976 276716 267028
rect 278044 266976 278096 267028
rect 286968 266976 287020 267028
rect 291292 266976 291344 267028
rect 295156 266976 295208 267028
rect 297088 266976 297140 267028
rect 316132 266976 316184 267028
rect 320180 266976 320232 267028
rect 324412 266976 324464 267028
rect 332508 266976 332560 267028
rect 353392 266976 353444 267028
rect 355324 266976 355376 267028
rect 378232 266976 378284 267028
rect 409144 266976 409196 267028
rect 422116 266976 422168 267028
rect 443460 266976 443512 267028
rect 209320 266840 209372 266892
rect 257988 266840 258040 266892
rect 320272 266840 320324 266892
rect 327448 266840 327500 266892
rect 342628 266840 342680 266892
rect 356520 266840 356572 266892
rect 359188 266840 359240 266892
rect 265072 266772 265124 266824
rect 268936 266772 268988 266824
rect 331864 266772 331916 266824
rect 335636 266772 335688 266824
rect 120724 266704 120776 266756
rect 157156 266704 157208 266756
rect 169024 266704 169076 266756
rect 172060 266704 172112 266756
rect 184020 266704 184072 266756
rect 189448 266704 189500 266756
rect 240692 266704 240744 266756
rect 245752 266704 245804 266756
rect 249064 266704 249116 266756
rect 251548 266704 251600 266756
rect 358360 266704 358412 266756
rect 360844 266704 360896 266756
rect 330208 266636 330260 266688
rect 334624 266636 334676 266688
rect 393136 266840 393188 266892
rect 401600 266840 401652 266892
rect 405556 266840 405608 266892
rect 425704 266840 425756 266892
rect 412180 266704 412232 266756
rect 373080 266636 373132 266688
rect 138664 266568 138716 266620
rect 119804 266432 119856 266484
rect 144920 266432 144972 266484
rect 149060 266568 149112 266620
rect 179512 266568 179564 266620
rect 213828 266568 213880 266620
rect 220084 266568 220136 266620
rect 245108 266568 245160 266620
rect 249064 266568 249116 266620
rect 360844 266568 360896 266620
rect 362224 266568 362276 266620
rect 417976 266704 418028 266756
rect 428464 266840 428516 266892
rect 435180 266840 435232 266892
rect 439320 266840 439372 266892
rect 427912 266704 427964 266756
rect 451924 266976 451976 267028
rect 455236 266976 455288 267028
rect 460204 266976 460256 267028
rect 462320 266976 462372 267028
rect 464988 266976 465040 267028
rect 465540 266976 465592 267028
rect 512920 266976 512972 267028
rect 513380 266976 513432 267028
rect 518808 266976 518860 267028
rect 518992 266976 519044 267028
rect 520096 266976 520148 267028
rect 520280 266976 520332 267028
rect 585784 267112 585836 267164
rect 523132 266976 523184 267028
rect 524328 266976 524380 267028
rect 524788 266976 524840 267028
rect 525708 266976 525760 267028
rect 525892 266976 525944 267028
rect 613384 266976 613436 267028
rect 421564 266568 421616 266620
rect 422944 266568 422996 266620
rect 435180 266568 435232 266620
rect 435364 266568 435416 266620
rect 471244 266840 471296 266892
rect 449440 266704 449492 266756
rect 145564 266500 145616 266552
rect 148876 266500 148928 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 327724 266500 327776 266552
rect 331680 266500 331732 266552
rect 346768 266500 346820 266552
rect 351644 266500 351696 266552
rect 355048 266500 355100 266552
rect 359740 266500 359792 266552
rect 394792 266500 394844 266552
rect 397920 266500 397972 266552
rect 444472 266500 444524 266552
rect 447784 266500 447836 266552
rect 456432 266704 456484 266756
rect 462320 266704 462372 266756
rect 452752 266636 452804 266688
rect 456156 266636 456208 266688
rect 459192 266568 459244 266620
rect 464528 266704 464580 266756
rect 464988 266704 465040 266756
rect 469220 266704 469272 266756
rect 462688 266568 462740 266620
rect 463516 266568 463568 266620
rect 464344 266568 464396 266620
rect 465724 266568 465776 266620
rect 469312 266568 469364 266620
rect 471796 266704 471848 266756
rect 475384 266704 475436 266756
rect 473452 266568 473504 266620
rect 474648 266568 474700 266620
rect 480904 266840 480956 266892
rect 492680 266840 492732 266892
rect 497464 266840 497516 266892
rect 499764 266840 499816 266892
rect 499948 266840 500000 266892
rect 500868 266840 500920 266892
rect 501052 266840 501104 266892
rect 506388 266840 506440 266892
rect 506572 266840 506624 266892
rect 507676 266840 507728 266892
rect 507860 266840 507912 266892
rect 570604 266840 570656 266892
rect 622400 266976 622452 267028
rect 475936 266704 475988 266756
rect 481088 266704 481140 266756
rect 481548 266704 481600 266756
rect 492312 266704 492364 266756
rect 492496 266704 492548 266756
rect 477316 266568 477368 266620
rect 477592 266568 477644 266620
rect 485688 266568 485740 266620
rect 486056 266568 486108 266620
rect 488724 266568 488776 266620
rect 490012 266568 490064 266620
rect 534080 266568 534132 266620
rect 453304 266500 453356 266552
rect 454408 266500 454460 266552
rect 457444 266500 457496 266552
rect 159824 266432 159876 266484
rect 162124 266432 162176 266484
rect 208676 266432 208728 266484
rect 210976 266432 211028 266484
rect 361672 266432 361724 266484
rect 362776 266432 362828 266484
rect 460204 266432 460256 266484
rect 147220 266364 147272 266416
rect 148324 266364 148376 266416
rect 149704 266364 149756 266416
rect 156604 266364 156656 266416
rect 159640 266364 159692 266416
rect 182180 266364 182232 266416
rect 186136 266364 186188 266416
rect 202144 266364 202196 266416
rect 206836 266364 206888 266416
rect 222844 266364 222896 266416
rect 224224 266364 224276 266416
rect 230756 266364 230808 266416
rect 236644 266364 236696 266416
rect 242256 266364 242308 266416
rect 243268 266364 243320 266416
rect 252008 266364 252060 266416
rect 257344 266364 257396 266416
rect 263324 266364 263376 266416
rect 265624 266364 265676 266416
rect 269120 266364 269172 266416
rect 276388 266364 276440 266416
rect 278596 266364 278648 266416
rect 286324 266364 286376 266416
rect 290464 266364 290516 266416
rect 292948 266364 293000 266416
rect 297916 266364 297968 266416
rect 299572 266364 299624 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 312360 266364 312412 266416
rect 314660 266364 314712 266416
rect 317788 266364 317840 266416
rect 323124 266364 323176 266416
rect 328552 266364 328604 266416
rect 329472 266364 329524 266416
rect 332692 266364 332744 266416
rect 333888 266364 333940 266416
rect 340972 266364 341024 266416
rect 342168 266364 342220 266416
rect 345112 266364 345164 266416
rect 346308 266364 346360 266416
rect 349252 266364 349304 266416
rect 350264 266364 350316 266416
rect 357532 266364 357584 266416
rect 358636 266364 358688 266416
rect 367468 266364 367520 266416
rect 368388 266364 368440 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375104 266364 375156 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412456 266364 412508 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 423772 266364 423824 266416
rect 424968 266364 425020 266416
rect 425428 266364 425480 266416
rect 426900 266364 426952 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 433708 266364 433760 266416
rect 434628 266364 434680 266416
rect 437020 266364 437072 266416
rect 440884 266364 440936 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 447784 266364 447836 266416
rect 449164 266364 449216 266416
rect 451924 266364 451976 266416
rect 454684 266364 454736 266416
rect 456892 266364 456944 266416
rect 458088 266364 458140 266416
rect 458548 266364 458600 266416
rect 459376 266364 459428 266416
rect 498568 266296 498620 266348
rect 501604 266296 501656 266348
rect 502800 266296 502852 266348
rect 507860 266296 507912 266348
rect 512368 266432 512420 266484
rect 513380 266432 513432 266484
rect 517336 266432 517388 266484
rect 538680 266568 538732 266620
rect 538864 266568 538916 266620
rect 552848 266704 552900 266756
rect 558920 266568 558972 266620
rect 552848 266432 552900 266484
rect 514668 266364 514720 266416
rect 514852 266364 514904 266416
rect 516784 266364 516836 266416
rect 518808 266296 518860 266348
rect 520280 266296 520332 266348
rect 522672 266296 522724 266348
rect 525892 266296 525944 266348
rect 527640 266296 527692 266348
rect 533896 266296 533948 266348
rect 534080 266296 534132 266348
rect 549628 266364 549680 266416
rect 475108 266024 475160 266076
rect 547880 266024 547932 266076
rect 485044 265888 485096 265940
rect 561680 265888 561732 265940
rect 494980 265752 495032 265804
rect 575848 265752 575900 265804
rect 187700 265616 187752 265668
rect 188252 265616 188304 265668
rect 247224 265616 247276 265668
rect 247868 265616 247920 265668
rect 259552 265616 259604 265668
rect 260380 265616 260432 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 480076 265616 480128 265668
rect 554780 265616 554832 265668
rect 558184 265616 558236 265668
rect 647240 265616 647292 265668
rect 533068 265072 533120 265124
rect 536564 265072 536616 265124
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 567844 259428 567896 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 562324 256708 562376 256760
rect 554504 253376 554556 253428
rect 559564 253376 559616 253428
rect 35808 252832 35860 252884
rect 40684 252832 40736 252884
rect 35624 252696 35676 252748
rect 41696 252696 41748 252748
rect 35440 252560 35492 252612
rect 41328 252560 41380 252612
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 675852 251540 675904 251592
rect 678428 251540 678480 251592
rect 35808 251200 35860 251252
rect 36544 251200 36596 251252
rect 553492 251200 553544 251252
rect 555424 251200 555476 251252
rect 553676 249024 553728 249076
rect 571340 249024 571392 249076
rect 553860 246304 553912 246356
rect 632704 246304 632756 246356
rect 554412 245624 554464 245676
rect 591304 245624 591356 245676
rect 554504 244264 554556 244316
rect 624424 244264 624476 244316
rect 36544 242836 36596 242888
rect 41696 242836 41748 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553952 241476 554004 241528
rect 628564 241476 628616 241528
rect 553860 240116 553912 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672172 237804 672224 237856
rect 671344 237600 671396 237652
rect 668768 237328 668820 237380
rect 671528 237192 671580 237244
rect 671620 236988 671672 237040
rect 673184 236716 673236 236768
rect 673414 236852 673466 236904
rect 673528 236648 673580 236700
rect 673644 236512 673696 236564
rect 673368 236240 673420 236292
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 673304 236036 673356 236088
rect 670332 235696 670384 235748
rect 672448 235696 672500 235748
rect 591304 235220 591356 235272
rect 633624 235220 633676 235272
rect 674196 234948 674248 235000
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 669780 234540 669832 234592
rect 674380 234744 674432 234796
rect 672264 234336 672316 234388
rect 675852 234540 675904 234592
rect 679624 234540 679676 234592
rect 669596 234200 669648 234252
rect 674564 234200 674616 234252
rect 675852 234336 675904 234388
rect 679992 234336 680044 234388
rect 674886 234268 674938 234320
rect 675852 234200 675904 234252
rect 679808 234200 679860 234252
rect 669136 234064 669188 234116
rect 673000 233928 673052 233980
rect 674932 233928 674984 233980
rect 675852 233928 675904 233980
rect 683488 233928 683540 233980
rect 670792 233588 670844 233640
rect 675236 233656 675288 233708
rect 675852 233520 675904 233572
rect 677784 233520 677836 233572
rect 671068 233452 671120 233504
rect 668308 233180 668360 233232
rect 674196 233180 674248 233232
rect 670884 233044 670936 233096
rect 674748 233044 674800 233096
rect 652024 232500 652076 232552
rect 675484 232568 675536 232620
rect 675852 232500 675904 232552
rect 680176 232500 680228 232552
rect 662328 232296 662380 232348
rect 675346 232296 675398 232348
rect 665088 232160 665140 232212
rect 675346 232024 675398 232076
rect 675180 231752 675232 231804
rect 672264 231548 672316 231600
rect 673368 231548 673420 231600
rect 675070 231480 675122 231532
rect 674956 231276 675008 231328
rect 675852 231208 675904 231260
rect 677600 231208 677652 231260
rect 674840 231140 674892 231192
rect 674732 230868 674784 230920
rect 668124 230800 668176 230852
rect 669412 230800 669464 230852
rect 673092 230800 673144 230852
rect 144644 230528 144696 230580
rect 150532 230528 150584 230580
rect 150900 230528 150952 230580
rect 158260 230664 158312 230716
rect 90364 230392 90416 230444
rect 439320 230528 439372 230580
rect 161112 230392 161164 230444
rect 161296 230392 161348 230444
rect 215208 230392 215260 230444
rect 223396 230392 223448 230444
rect 271880 230392 271932 230444
rect 274180 230392 274232 230444
rect 307944 230392 307996 230444
rect 312544 230392 312596 230444
rect 315672 230392 315724 230444
rect 377404 230392 377456 230444
rect 378784 230392 378836 230444
rect 674518 230460 674570 230512
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 444472 230392 444524 230444
rect 447600 230392 447652 230444
rect 528008 230392 528060 230444
rect 529020 230392 529072 230444
rect 534632 230392 534684 230444
rect 544200 230392 544252 230444
rect 671804 230392 671856 230444
rect 404268 230324 404320 230376
rect 412272 230324 412324 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 448336 230324 448388 230376
rect 449164 230324 449216 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 475384 230324 475436 230376
rect 478328 230324 478380 230376
rect 480536 230324 480588 230376
rect 481548 230324 481600 230376
rect 492772 230324 492824 230376
rect 493968 230324 494020 230376
rect 513380 230324 513432 230376
rect 515404 230324 515456 230376
rect 520464 230324 520516 230376
rect 521568 230324 521620 230376
rect 526904 230324 526956 230376
rect 527824 230324 527876 230376
rect 118424 230256 118476 230308
rect 189448 230256 189500 230308
rect 190920 230256 190972 230308
rect 111064 230120 111116 230172
rect 184296 230120 184348 230172
rect 88248 229984 88300 230036
rect 166264 229984 166316 230036
rect 166632 229984 166684 230036
rect 181720 229984 181772 230036
rect 184204 229984 184256 230036
rect 191564 230120 191616 230172
rect 196992 230256 197044 230308
rect 202328 230120 202380 230172
rect 205364 230256 205416 230308
rect 256424 230256 256476 230308
rect 276296 230256 276348 230308
rect 313096 230256 313148 230308
rect 251272 230120 251324 230172
rect 261392 230120 261444 230172
rect 297640 230120 297692 230172
rect 308128 230120 308180 230172
rect 323400 230256 323452 230308
rect 436100 230256 436152 230308
rect 436836 230256 436888 230308
rect 497924 230256 497976 230308
rect 504364 230256 504416 230308
rect 528836 230256 528888 230308
rect 541624 230256 541676 230308
rect 408868 230188 408920 230240
rect 410984 230188 411036 230240
rect 443828 230188 443880 230240
rect 444656 230188 444708 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 454132 230188 454184 230240
rect 455236 230188 455288 230240
rect 470876 230188 470928 230240
rect 471888 230188 471940 230240
rect 476672 230188 476724 230240
rect 479708 230188 479760 230240
rect 493416 230188 493468 230240
rect 495164 230188 495216 230240
rect 511448 230188 511500 230240
rect 516508 230188 516560 230240
rect 668124 230188 668176 230240
rect 674104 230188 674156 230240
rect 315304 230120 315356 230172
rect 340144 230120 340196 230172
rect 302884 230052 302936 230104
rect 305368 230052 305420 230104
rect 345664 230052 345716 230104
rect 353024 230052 353076 230104
rect 453488 230052 453540 230104
rect 455788 230052 455840 230104
rect 476028 230052 476080 230104
rect 479524 230052 479576 230104
rect 490840 230052 490892 230104
rect 493784 230052 493836 230104
rect 494336 230052 494388 230104
rect 503260 230120 503312 230172
rect 521108 230120 521160 230172
rect 529940 230120 529992 230172
rect 536564 230120 536616 230172
rect 549260 230120 549312 230172
rect 674288 230052 674340 230104
rect 190184 229984 190236 230036
rect 246120 229984 246172 230036
rect 251732 229984 251784 230036
rect 292488 229984 292540 230036
rect 296996 229984 297048 230036
rect 302516 229984 302568 230036
rect 305644 229984 305696 230036
rect 334992 229984 335044 230036
rect 380440 229984 380492 230036
rect 389088 229984 389140 230036
rect 410892 229984 410944 230036
rect 417424 229984 417476 230036
rect 447048 229984 447100 230036
rect 449900 229984 449952 230036
rect 467012 229984 467064 230036
rect 474004 229984 474056 230036
rect 483112 229984 483164 230036
rect 484308 229984 484360 230036
rect 484768 229984 484820 230036
rect 490656 229984 490708 230036
rect 503720 229984 503772 230036
rect 506940 229984 506992 230036
rect 509516 229984 509568 230036
rect 518900 229984 518952 230036
rect 519176 229984 519228 230036
rect 528008 229984 528060 230036
rect 530768 229984 530820 230036
rect 547144 229984 547196 230036
rect 555424 229984 555476 230036
rect 569960 229984 570012 230036
rect 675852 229984 675904 230036
rect 676588 229984 676640 230036
rect 674172 229916 674224 229968
rect 74448 229848 74500 229900
rect 155960 229848 156012 229900
rect 156328 229848 156380 229900
rect 176568 229848 176620 229900
rect 177580 229848 177632 229900
rect 67548 229712 67600 229764
rect 144644 229712 144696 229764
rect 144828 229712 144880 229764
rect 140044 229576 140096 229628
rect 146944 229576 146996 229628
rect 148600 229712 148652 229764
rect 150900 229712 150952 229764
rect 151360 229712 151412 229764
rect 190920 229712 190972 229764
rect 191564 229848 191616 229900
rect 240968 229848 241020 229900
rect 245660 229848 245712 229900
rect 287336 229848 287388 229900
rect 300124 229848 300176 229900
rect 329840 229848 329892 229900
rect 334256 229848 334308 229900
rect 345296 229848 345348 229900
rect 352564 229848 352616 229900
rect 358176 229848 358228 229900
rect 364156 229848 364208 229900
rect 381360 229848 381412 229900
rect 384304 229848 384356 229900
rect 394240 229848 394292 229900
rect 468944 229848 468996 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 235816 229712 235868 229764
rect 236920 229712 236972 229764
rect 282184 229712 282236 229764
rect 285312 229712 285364 229764
rect 318248 229712 318300 229764
rect 324044 229712 324096 229764
rect 350448 229712 350500 229764
rect 210056 229576 210108 229628
rect 210240 229576 210292 229628
rect 261576 229576 261628 229628
rect 350540 229576 350592 229628
rect 371056 229712 371108 229764
rect 370964 229576 371016 229628
rect 386512 229712 386564 229764
rect 386972 229712 387024 229764
rect 396816 229712 396868 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 412456 229712 412508 229764
rect 419356 229712 419408 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 468300 229712 468352 229764
rect 469128 229712 469180 229764
rect 469588 229848 469640 229900
rect 476764 229848 476816 229900
rect 479248 229848 479300 229900
rect 484032 229848 484084 229900
rect 486332 229848 486384 229900
rect 500224 229848 500276 229900
rect 505652 229848 505704 229900
rect 516048 229848 516100 229900
rect 517428 229848 517480 229900
rect 522304 229848 522356 229900
rect 523040 229848 523092 229900
rect 534724 229848 534776 229900
rect 538496 229848 538548 229900
rect 556804 229848 556856 229900
rect 674058 229848 674110 229900
rect 675852 229848 675904 229900
rect 677232 229848 677284 229900
rect 475384 229712 475436 229764
rect 481824 229712 481876 229764
rect 489920 229712 489972 229764
rect 495992 229712 496044 229764
rect 509240 229712 509292 229764
rect 515680 229712 515732 229764
rect 525524 229712 525576 229764
rect 532700 229712 532752 229764
rect 555608 229712 555660 229764
rect 675852 229712 675904 229764
rect 676956 229712 677008 229764
rect 455420 229576 455472 229628
rect 457168 229576 457220 229628
rect 490656 229576 490708 229628
rect 497464 229576 497516 229628
rect 524972 229576 525024 229628
rect 532424 229576 532476 229628
rect 448980 229508 449032 229560
rect 451372 229508 451424 229560
rect 673948 229508 674000 229560
rect 131120 229440 131172 229492
rect 197176 229440 197228 229492
rect 203892 229440 203944 229492
rect 205364 229440 205416 229492
rect 231124 229440 231176 229492
rect 277032 229440 277084 229492
rect 499856 229440 499908 229492
rect 501328 229440 501380 229492
rect 673460 229440 673512 229492
rect 446404 229372 446456 229424
rect 448612 229372 448664 229424
rect 450912 229372 450964 229424
rect 453028 229372 453080 229424
rect 501788 229372 501840 229424
rect 507124 229372 507176 229424
rect 92480 229304 92532 229356
rect 146300 229304 146352 229356
rect 146944 229304 146996 229356
rect 153384 229304 153436 229356
rect 153844 229304 153896 229356
rect 163688 229304 163740 229356
rect 163872 229304 163924 229356
rect 166632 229304 166684 229356
rect 167644 229304 167696 229356
rect 220360 229304 220412 229356
rect 494704 229304 494756 229356
rect 496360 229304 496412 229356
rect 673092 229304 673144 229356
rect 358084 229236 358136 229288
rect 360752 229236 360804 229288
rect 360936 229236 360988 229288
rect 363328 229236 363380 229288
rect 419448 229236 419500 229288
rect 424508 229236 424560 229288
rect 450268 229236 450320 229288
rect 451832 229236 451884 229288
rect 479892 229236 479944 229288
rect 482284 229236 482336 229288
rect 483756 229236 483808 229288
rect 486792 229236 486844 229288
rect 115756 229168 115808 229220
rect 106188 229032 106240 229084
rect 122932 229168 122984 229220
rect 179144 229168 179196 229220
rect 181628 229168 181680 229220
rect 230664 229168 230716 229220
rect 669320 229168 669372 229220
rect 673276 229168 673328 229220
rect 675852 229168 675904 229220
rect 378968 229100 379020 229152
rect 383936 229100 383988 229152
rect 97908 228896 97960 228948
rect 82084 228624 82136 228676
rect 106648 228760 106700 228812
rect 107016 228896 107068 228948
rect 115572 228896 115624 228948
rect 116032 229032 116084 229084
rect 179788 229032 179840 229084
rect 180616 229032 180668 229084
rect 116400 228896 116452 228948
rect 184940 228896 184992 228948
rect 185676 229032 185728 229084
rect 190368 229032 190420 229084
rect 194600 229032 194652 229084
rect 195704 229032 195756 229084
rect 250628 229032 250680 229084
rect 259276 229032 259328 229084
rect 298284 229032 298336 229084
rect 413836 229032 413888 229084
rect 420000 229100 420052 229152
rect 420184 229100 420236 229152
rect 421932 229100 421984 229152
rect 424324 229100 424376 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 507584 229100 507636 229152
rect 511264 229100 511316 229152
rect 517888 229032 517940 229084
rect 540244 229032 540296 229084
rect 673460 229032 673512 229084
rect 675852 229032 675904 229084
rect 677048 229032 677100 229084
rect 677416 229032 677468 229084
rect 173992 228760 174044 228812
rect 174176 228760 174228 228812
rect 96252 228624 96304 228676
rect 172060 228624 172112 228676
rect 172244 228624 172296 228676
rect 175280 228624 175332 228676
rect 175740 228760 175792 228812
rect 188344 228760 188396 228812
rect 241612 228896 241664 228948
rect 251088 228896 251140 228948
rect 291200 228896 291252 228948
rect 319812 228896 319864 228948
rect 345940 228896 345992 228948
rect 350172 228896 350224 228948
rect 369124 228896 369176 228948
rect 507124 228896 507176 228948
rect 520188 228896 520240 228948
rect 526260 228896 526312 228948
rect 551652 228896 551704 228948
rect 673506 228828 673558 228880
rect 204720 228760 204772 228812
rect 204904 228760 204956 228812
rect 210700 228760 210752 228812
rect 214104 228760 214156 228812
rect 218428 228760 218480 228812
rect 219348 228760 219400 228812
rect 224040 228760 224092 228812
rect 231308 228760 231360 228812
rect 246304 228760 246356 228812
rect 253848 228760 253900 228812
rect 255136 228760 255188 228812
rect 295708 228760 295760 228812
rect 317972 228760 318024 228812
rect 344652 228760 344704 228812
rect 346216 228760 346268 228812
rect 366548 228760 366600 228812
rect 376576 228760 376628 228812
rect 389732 228760 389784 228812
rect 401416 228760 401468 228812
rect 408408 228760 408460 228812
rect 493784 228760 493836 228812
rect 506020 228760 506072 228812
rect 519820 228760 519872 228812
rect 543188 228760 543240 228812
rect 675852 228760 675904 228812
rect 676220 228760 676272 228812
rect 62764 228488 62816 228540
rect 140780 228488 140832 228540
rect 140964 228488 141016 228540
rect 66168 228352 66220 228404
rect 147634 228352 147686 228404
rect 153292 228488 153344 228540
rect 204904 228488 204956 228540
rect 205088 228488 205140 228540
rect 237104 228624 237156 228676
rect 239404 228624 239456 228676
rect 284116 228624 284168 228676
rect 292396 228624 292448 228676
rect 326620 228624 326672 228676
rect 333244 228624 333296 228676
rect 355600 228624 355652 228676
rect 157432 228352 157484 228404
rect 157800 228352 157852 228404
rect 214104 228352 214156 228404
rect 102048 228216 102100 228268
rect 171048 228216 171100 228268
rect 171232 228216 171284 228268
rect 222752 228352 222804 228404
rect 224040 228352 224092 228404
rect 267372 228488 267424 228540
rect 267556 228488 267608 228540
rect 307300 228488 307352 228540
rect 307668 228488 307720 228540
rect 335636 228488 335688 228540
rect 336648 228488 336700 228540
rect 358820 228488 358872 228540
rect 225696 228352 225748 228404
rect 273812 228352 273864 228404
rect 284116 228352 284168 228404
rect 320180 228352 320232 228404
rect 326896 228352 326948 228404
rect 351092 228352 351144 228404
rect 355232 228352 355284 228404
rect 369768 228624 369820 228676
rect 373816 228624 373868 228676
rect 387248 228624 387300 228676
rect 390284 228624 390336 228676
rect 400036 228624 400088 228676
rect 410892 228624 410944 228676
rect 416136 228624 416188 228676
rect 478788 228624 478840 228676
rect 483572 228624 483624 228676
rect 495348 228624 495400 228676
rect 511816 228624 511868 228676
rect 512092 228624 512144 228676
rect 366916 228488 366968 228540
rect 382004 228488 382056 228540
rect 362868 228352 362920 228404
rect 379428 228352 379480 228404
rect 381728 228352 381780 228404
rect 392952 228488 393004 228540
rect 393228 228488 393280 228540
rect 391848 228352 391900 228404
rect 400128 228488 400180 228540
rect 407764 228488 407816 228540
rect 482468 228488 482520 228540
rect 494612 228488 494664 228540
rect 502432 228488 502484 228540
rect 520924 228488 520976 228540
rect 214748 228216 214800 228268
rect 257068 228216 257120 228268
rect 277216 228216 277268 228268
rect 311808 228216 311860 228268
rect 402612 228352 402664 228404
rect 409788 228352 409840 228404
rect 415492 228352 415544 228404
rect 487620 228352 487672 228404
rect 501512 228352 501564 228404
rect 506296 228352 506348 228404
rect 525892 228352 525944 228404
rect 533988 228624 534040 228676
rect 561588 228624 561640 228676
rect 531412 228488 531464 228540
rect 558184 228488 558236 228540
rect 673388 228488 673440 228540
rect 672172 228420 672224 228472
rect 533896 228352 533948 228404
rect 537852 228352 537904 228404
rect 566372 228352 566424 228404
rect 403900 228216 403952 228268
rect 479708 228216 479760 228268
rect 487804 228216 487856 228268
rect 671804 228216 671856 228268
rect 112996 228080 113048 228132
rect 115756 228080 115808 228132
rect 115572 227944 115624 227996
rect 140964 228080 141016 228132
rect 141148 228080 141200 228132
rect 201040 228080 201092 228132
rect 201408 228080 201460 228132
rect 252560 228080 252612 228132
rect 288164 228080 288216 228132
rect 321468 228080 321520 228132
rect 484032 228080 484084 228132
rect 490564 228080 490616 228132
rect 122748 227944 122800 227996
rect 192668 227944 192720 227996
rect 197912 227944 197964 227996
rect 204536 227944 204588 227996
rect 205456 227944 205508 227996
rect 214748 227944 214800 227996
rect 222752 227944 222804 227996
rect 226156 227944 226208 227996
rect 134616 227808 134668 227860
rect 141148 227808 141200 227860
rect 141332 227808 141384 227860
rect 200396 227808 200448 227860
rect 226156 227808 226208 227860
rect 272524 227944 272576 227996
rect 369124 227876 369176 227928
rect 375564 227876 375616 227928
rect 407764 227876 407816 227928
rect 411628 227876 411680 227928
rect 471520 227876 471572 227928
rect 479340 227876 479392 227928
rect 673046 227876 673098 227928
rect 242716 227740 242768 227792
rect 245660 227740 245712 227792
rect 255964 227740 256016 227792
rect 259000 227740 259052 227792
rect 366364 227740 366416 227792
rect 372988 227740 373040 227792
rect 393964 227740 394016 227792
rect 395528 227740 395580 227792
rect 396632 227740 396684 227792
rect 397460 227740 397512 227792
rect 402244 227740 402296 227792
rect 403256 227740 403308 227792
rect 404084 227740 404136 227792
rect 408868 227740 408920 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416688 227740 416740 227792
rect 420644 227740 420696 227792
rect 475016 227740 475068 227792
rect 482928 227740 482980 227792
rect 110144 227672 110196 227724
rect 182364 227672 182416 227724
rect 186688 227672 186740 227724
rect 187240 227672 187292 227724
rect 191564 227672 191616 227724
rect 270132 227672 270184 227724
rect 306656 227672 306708 227724
rect 321376 227672 321428 227724
rect 346584 227672 346636 227724
rect 525524 227672 525576 227724
rect 537576 227672 537628 227724
rect 672954 227672 673006 227724
rect 248052 227604 248104 227656
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 100668 227536 100720 227588
rect 174636 227536 174688 227588
rect 179052 227536 179104 227588
rect 236460 227536 236512 227588
rect 252468 227536 252520 227588
rect 293132 227536 293184 227588
rect 299296 227536 299348 227588
rect 328552 227536 328604 227588
rect 359372 227536 359424 227588
rect 374920 227536 374972 227588
rect 515864 227536 515916 227588
rect 538864 227536 538916 227588
rect 663708 227536 663760 227588
rect 665548 227536 665600 227588
rect 672816 227468 672868 227520
rect 89628 227400 89680 227452
rect 159640 227400 159692 227452
rect 160008 227400 160060 227452
rect 166908 227400 166960 227452
rect 86868 227264 86920 227316
rect 151912 227264 151964 227316
rect 152924 227264 152976 227316
rect 164332 227264 164384 227316
rect 165436 227264 165488 227316
rect 175188 227400 175240 227452
rect 231952 227400 232004 227452
rect 248236 227400 248288 227452
rect 291844 227400 291896 227452
rect 293776 227400 293828 227452
rect 325332 227400 325384 227452
rect 340604 227400 340656 227452
rect 361396 227400 361448 227452
rect 227444 227264 227496 227316
rect 75828 227128 75880 227180
rect 150164 227128 150216 227180
rect 150348 227128 150400 227180
rect 57888 226992 57940 227044
rect 135260 226992 135312 227044
rect 135444 226992 135496 227044
rect 151912 226992 151964 227044
rect 152280 227128 152332 227180
rect 168840 227128 168892 227180
rect 169576 227128 169628 227180
rect 228732 227128 228784 227180
rect 213276 226992 213328 227044
rect 226892 226992 226944 227044
rect 233240 227264 233292 227316
rect 234528 227264 234580 227316
rect 278320 227264 278372 227316
rect 280712 227264 280764 227316
rect 312084 227264 312136 227316
rect 326344 227264 326396 227316
rect 352380 227264 352432 227316
rect 361212 227264 361264 227316
rect 377220 227400 377272 227452
rect 361764 227264 361816 227316
rect 372344 227264 372396 227316
rect 373264 227264 373316 227316
rect 383292 227400 383344 227452
rect 524328 227400 524380 227452
rect 547880 227400 547932 227452
rect 382924 227264 382976 227316
rect 391664 227264 391716 227316
rect 395988 227264 396040 227316
rect 406476 227264 406528 227316
rect 485044 227264 485096 227316
rect 498752 227264 498804 227316
rect 501328 227264 501380 227316
rect 517704 227264 517756 227316
rect 521752 227264 521804 227316
rect 545764 227264 545816 227316
rect 672724 227264 672776 227316
rect 672264 227196 672316 227248
rect 235908 227128 235960 227180
rect 280252 227128 280304 227180
rect 296444 227128 296496 227180
rect 329196 227128 329248 227180
rect 329748 227128 329800 227180
rect 353668 227128 353720 227180
rect 354588 227128 354640 227180
rect 373632 227128 373684 227180
rect 381912 227128 381964 227180
rect 396172 227128 396224 227180
rect 481180 227128 481232 227180
rect 492956 227128 493008 227180
rect 498568 227128 498620 227180
rect 515864 227128 515916 227180
rect 516048 227128 516100 227180
rect 525064 227128 525116 227180
rect 535920 227128 535972 227180
rect 564072 227128 564124 227180
rect 229054 226992 229106 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 308772 226992 308824 227044
rect 336280 226992 336332 227044
rect 336464 226992 336516 227044
rect 360108 226992 360160 227044
rect 369768 226992 369820 227044
rect 385868 226992 385920 227044
rect 386328 226992 386380 227044
rect 398748 226992 398800 227044
rect 472164 226992 472216 227044
rect 481180 226992 481232 227044
rect 497280 226992 497332 227044
rect 106924 226856 106976 226908
rect 125784 226856 125836 226908
rect 121092 226720 121144 226772
rect 190736 226856 190788 226908
rect 200028 226856 200080 226908
rect 251916 226856 251968 226908
rect 272432 226856 272484 226908
rect 284760 226856 284812 226908
rect 355508 226856 355560 226908
rect 361764 226856 361816 226908
rect 398472 226856 398524 226908
rect 408684 226856 408736 226908
rect 514024 226992 514076 227044
rect 536012 226992 536064 227044
rect 537208 226992 537260 227044
rect 565728 226992 565780 227044
rect 671068 226992 671120 227044
rect 514300 226856 514352 226908
rect 672264 226856 672316 226908
rect 119988 226584 120040 226636
rect 189724 226720 189776 226772
rect 195888 226720 195940 226772
rect 199292 226720 199344 226772
rect 212172 226720 212224 226772
rect 262220 226720 262272 226772
rect 125784 226448 125836 226500
rect 135444 226584 135496 226636
rect 135628 226584 135680 226636
rect 129372 226448 129424 226500
rect 137192 226448 137244 226500
rect 137560 226584 137612 226636
rect 197360 226584 197412 226636
rect 222016 226584 222068 226636
rect 269948 226584 270000 226636
rect 669412 226584 669464 226636
rect 142114 226448 142166 226500
rect 142252 226448 142304 226500
rect 205272 226448 205324 226500
rect 213184 226448 213236 226500
rect 217784 226448 217836 226500
rect 221832 226448 221884 226500
rect 229008 226448 229060 226500
rect 232504 226448 232556 226500
rect 266728 226448 266780 226500
rect 666836 226448 666888 226500
rect 291844 226380 291896 226432
rect 295064 226380 295116 226432
rect 83464 226244 83516 226296
rect 69572 226108 69624 226160
rect 143540 226108 143592 226160
rect 166954 226312 167006 226364
rect 221004 226312 221056 226364
rect 152832 226244 152884 226296
rect 161940 226244 161992 226296
rect 162308 226244 162360 226296
rect 166816 226244 166868 226296
rect 222476 226244 222528 226296
rect 225512 226244 225564 226296
rect 228732 226244 228784 226296
rect 275100 226244 275152 226296
rect 278504 226244 278556 226296
rect 315028 226244 315080 226296
rect 317328 226244 317380 226296
rect 334256 226244 334308 226296
rect 503260 226244 503312 226296
rect 510160 226244 510212 226296
rect 529940 226244 529992 226296
rect 544936 226244 544988 226296
rect 562324 226244 562376 226296
rect 568396 226244 568448 226296
rect 671068 226244 671120 226296
rect 157432 226108 157484 226160
rect 157616 226108 157668 226160
rect 215852 226108 215904 226160
rect 216496 226108 216548 226160
rect 264796 226108 264848 226160
rect 266268 226108 266320 226160
rect 303436 226108 303488 226160
rect 325424 226108 325476 226160
rect 349160 226108 349212 226160
rect 510804 226108 510856 226160
rect 531688 226108 531740 226160
rect 667020 226040 667072 226092
rect 93768 225972 93820 226024
rect 161572 225972 161624 226024
rect 161940 225972 161992 226024
rect 171048 225972 171100 226024
rect 171232 225972 171284 226024
rect 186274 225972 186326 226024
rect 186412 225972 186464 226024
rect 224224 225972 224276 226024
rect 95148 225836 95200 225888
rect 166816 225836 166868 225888
rect 166954 225836 167006 225888
rect 64788 225700 64840 225752
rect 92480 225700 92532 225752
rect 108304 225700 108356 225752
rect 171048 225700 171100 225752
rect 171232 225700 171284 225752
rect 175924 225700 175976 225752
rect 176292 225836 176344 225888
rect 176614 225836 176666 225888
rect 176752 225836 176804 225888
rect 181076 225836 181128 225888
rect 185952 225836 186004 225888
rect 186136 225836 186188 225888
rect 233884 225972 233936 226024
rect 243452 225972 243504 226024
rect 248696 225972 248748 226024
rect 267694 225972 267746 226024
rect 304080 225972 304132 226024
rect 313096 225972 313148 226024
rect 340788 225972 340840 226024
rect 181444 225700 181496 225752
rect 186688 225700 186740 225752
rect 186872 225700 186924 225752
rect 239036 225836 239088 225888
rect 249708 225836 249760 225888
rect 290556 225836 290608 225888
rect 294972 225836 295024 225888
rect 325976 225836 326028 225888
rect 340144 225836 340196 225888
rect 347872 225972 347924 226024
rect 349068 225972 349120 226024
rect 367192 225972 367244 226024
rect 518532 225972 518584 226024
rect 541440 225972 541492 226024
rect 544200 225972 544252 226024
rect 561956 225972 562008 226024
rect 347044 225836 347096 225888
rect 365904 225836 365956 225888
rect 367652 225836 367704 225888
rect 379612 225836 379664 225888
rect 488908 225836 488960 225888
rect 503076 225836 503128 225888
rect 528192 225836 528244 225888
rect 554044 225836 554096 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 61292 225564 61344 225616
rect 136824 225564 136876 225616
rect 137008 225564 137060 225616
rect 147036 225564 147088 225616
rect 147404 225564 147456 225616
rect 203892 225564 203944 225616
rect 204904 225564 204956 225616
rect 222476 225564 222528 225616
rect 224224 225564 224276 225616
rect 242900 225700 242952 225752
rect 257712 225700 257764 225752
rect 299572 225700 299624 225752
rect 304908 225700 304960 225752
rect 333704 225700 333756 225752
rect 335268 225700 335320 225752
rect 356888 225700 356940 225752
rect 379336 225700 379388 225752
rect 393596 225700 393648 225752
rect 394608 225700 394660 225752
rect 404544 225700 404596 225752
rect 491484 225700 491536 225752
rect 506848 225700 506900 225752
rect 507308 225700 507360 225752
rect 526352 225700 526404 225752
rect 527548 225700 527600 225752
rect 553308 225700 553360 225752
rect 671820 225700 671872 225752
rect 234344 225564 234396 225616
rect 281540 225564 281592 225616
rect 285496 225564 285548 225616
rect 318892 225564 318944 225616
rect 322848 225564 322900 225616
rect 349804 225564 349856 225616
rect 351184 225564 351236 225616
rect 370412 225564 370464 225616
rect 372528 225564 372580 225616
rect 388076 225564 388128 225616
rect 388444 225564 388496 225616
rect 399392 225564 399444 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 489184 225564 489236 225616
rect 495164 225564 495216 225616
rect 509700 225564 509752 225616
rect 510344 225564 510396 225616
rect 530952 225564 531004 225616
rect 532056 225564 532108 225616
rect 558920 225564 558972 225616
rect 671712 225496 671764 225548
rect 103428 225428 103480 225480
rect 108304 225428 108356 225480
rect 106004 225292 106056 225344
rect 127440 225428 127492 225480
rect 117228 225292 117280 225344
rect 181444 225428 181496 225480
rect 183284 225428 183336 225480
rect 185676 225428 185728 225480
rect 190736 225428 190788 225480
rect 242256 225428 242308 225480
rect 668400 225428 668452 225480
rect 127440 225156 127492 225208
rect 137008 225292 137060 225344
rect 128268 225156 128320 225208
rect 142114 225292 142166 225344
rect 142252 225292 142304 225344
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 203156 225292 203208 225344
rect 203892 225292 203944 225344
rect 207756 225292 207808 225344
rect 208032 225292 208084 225344
rect 260932 225292 260984 225344
rect 671068 225224 671120 225276
rect 126888 225020 126940 225072
rect 186872 225156 186924 225208
rect 187240 225156 187292 225208
rect 195888 225156 195940 225208
rect 199384 225156 199436 225208
rect 204904 225156 204956 225208
rect 205088 225156 205140 225208
rect 254492 225156 254544 225208
rect 137468 225020 137520 225072
rect 141516 225020 141568 225072
rect 141792 225020 141844 225072
rect 116768 224884 116820 224936
rect 122932 224884 122984 224936
rect 123484 224884 123536 224936
rect 142068 224884 142120 224936
rect 142436 225020 142488 225072
rect 162308 225020 162360 225072
rect 162492 225020 162544 225072
rect 166540 225020 166592 225072
rect 166724 225020 166776 225072
rect 169024 225020 169076 225072
rect 169208 225020 169260 225072
rect 170864 225020 170916 225072
rect 171048 225020 171100 225072
rect 223580 225020 223632 225072
rect 224868 225020 224920 225072
rect 270592 225020 270644 225072
rect 669412 225020 669464 225072
rect 275836 224952 275888 225004
rect 276296 224952 276348 225004
rect 282736 224952 282788 225004
rect 285312 224952 285364 225004
rect 489920 224952 489972 225004
rect 494796 224952 494848 225004
rect 509240 224952 509292 225004
rect 512644 224952 512696 225004
rect 209412 224884 209464 224936
rect 209688 224884 209740 224936
rect 259644 224884 259696 224936
rect 264152 224884 264204 224936
rect 269304 224884 269356 224936
rect 288348 224884 288400 224936
rect 322388 224884 322440 224936
rect 406752 224884 406804 224936
rect 414848 224884 414900 224936
rect 516508 224884 516560 224936
rect 531320 224884 531372 224936
rect 669412 224816 669464 224868
rect 118608 224748 118660 224800
rect 177212 224748 177264 224800
rect 177396 224748 177448 224800
rect 181260 224748 181312 224800
rect 115756 224612 115808 224664
rect 187056 224748 187108 224800
rect 187332 224748 187384 224800
rect 190736 224748 190788 224800
rect 194508 224748 194560 224800
rect 247408 224748 247460 224800
rect 282552 224748 282604 224800
rect 316316 224748 316368 224800
rect 532424 224748 532476 224800
rect 550456 224748 550508 224800
rect 460572 224680 460624 224732
rect 463148 224680 463200 224732
rect 60648 224476 60700 224528
rect 103612 224476 103664 224528
rect 108672 224476 108724 224528
rect 177028 224476 177080 224528
rect 177212 224476 177264 224528
rect 191380 224612 191432 224664
rect 192760 224612 192812 224664
rect 194324 224612 194376 224664
rect 195612 224612 195664 224664
rect 248880 224612 248932 224664
rect 249064 224612 249116 224664
rect 263876 224612 263928 224664
rect 271604 224612 271656 224664
rect 309876 224612 309928 224664
rect 315856 224612 315908 224664
rect 341432 224612 341484 224664
rect 344652 224612 344704 224664
rect 364616 224612 364668 224664
rect 514668 224612 514720 224664
rect 536656 224612 536708 224664
rect 668400 224612 668452 224664
rect 456064 224544 456116 224596
rect 459652 224544 459704 224596
rect 181720 224476 181772 224528
rect 183836 224476 183888 224528
rect 184020 224476 184072 224528
rect 233700 224476 233752 224528
rect 233884 224476 233936 224528
rect 246764 224476 246816 224528
rect 247684 224476 247736 224528
rect 289268 224476 289320 224528
rect 319996 224476 320048 224528
rect 347228 224476 347280 224528
rect 479524 224476 479576 224528
rect 486608 224476 486660 224528
rect 508228 224476 508280 224528
rect 528376 224476 528428 224528
rect 530124 224476 530176 224528
rect 556528 224476 556580 224528
rect 82728 224340 82780 224392
rect 123484 224340 123536 224392
rect 131304 224340 131356 224392
rect 193956 224340 194008 224392
rect 194140 224340 194192 224392
rect 204904 224340 204956 224392
rect 205088 224340 205140 224392
rect 255780 224340 255832 224392
rect 261852 224340 261904 224392
rect 300860 224340 300912 224392
rect 303252 224340 303304 224392
rect 333060 224340 333112 224392
rect 333888 224340 333940 224392
rect 356244 224340 356296 224392
rect 357348 224340 357400 224392
rect 374276 224340 374328 224392
rect 375288 224340 375340 224392
rect 387800 224340 387852 224392
rect 462504 224340 462556 224392
rect 469312 224340 469364 224392
rect 470232 224340 470284 224392
rect 479708 224340 479760 224392
rect 486792 224340 486844 224392
rect 496912 224340 496964 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525708 224340 525760 224392
rect 550640 224340 550692 224392
rect 58992 224204 59044 224256
rect 145196 224204 145248 224256
rect 145380 224204 145432 224256
rect 147220 224204 147272 224256
rect 147772 224204 147824 224256
rect 156696 224204 156748 224256
rect 157432 224204 157484 224256
rect 170956 224204 171008 224256
rect 171094 224204 171146 224256
rect 186872 224204 186924 224256
rect 187056 224204 187108 224256
rect 188804 224204 188856 224256
rect 188988 224204 189040 224256
rect 243820 224204 243872 224256
rect 246948 224204 247000 224256
rect 288624 224204 288676 224256
rect 289636 224204 289688 224256
rect 308128 224204 308180 224256
rect 308956 224204 309008 224256
rect 339500 224204 339552 224256
rect 342076 224204 342128 224256
rect 364800 224204 364852 224256
rect 364984 224204 365036 224256
rect 378140 224204 378192 224256
rect 389088 224204 389140 224256
rect 400956 224204 401008 224256
rect 416504 224204 416556 224256
rect 422208 224204 422260 224256
rect 423312 224204 423364 224256
rect 424324 224204 424376 224256
rect 451372 224204 451424 224256
rect 452200 224204 452252 224256
rect 474740 224204 474792 224256
rect 484584 224204 484636 224256
rect 485688 224204 485740 224256
rect 499396 224204 499448 224256
rect 508872 224204 508924 224256
rect 529204 224204 529256 224256
rect 535276 224204 535328 224256
rect 563704 224204 563756 224256
rect 104808 224068 104860 224120
rect 116768 224068 116820 224120
rect 116952 224068 117004 224120
rect 118424 224068 118476 224120
rect 121920 224068 121972 224120
rect 131304 224068 131356 224120
rect 131488 224068 131540 224120
rect 192760 224068 192812 224120
rect 192944 224068 192996 224120
rect 194140 224068 194192 224120
rect 194324 224068 194376 224120
rect 196532 224068 196584 224120
rect 201224 224068 201276 224120
rect 204720 224068 204772 224120
rect 204904 224068 204956 224120
rect 233884 224068 233936 224120
rect 76564 223932 76616 223984
rect 140964 223932 141016 223984
rect 142068 223932 142120 223984
rect 157064 223932 157116 223984
rect 157248 223932 157300 223984
rect 217140 223932 217192 223984
rect 217324 223932 217376 223984
rect 228088 223932 228140 223984
rect 231676 223932 231728 223984
rect 278964 224068 279016 224120
rect 286692 224068 286744 224120
rect 319536 224068 319588 224120
rect 670930 224272 670982 224324
rect 238668 223932 238720 223984
rect 282368 223932 282420 223984
rect 670700 223932 670752 223984
rect 125232 223796 125284 223848
rect 131488 223796 131540 223848
rect 134432 223796 134484 223848
rect 204260 223796 204312 223848
rect 205272 223796 205324 223848
rect 212632 223796 212684 223848
rect 215944 223796 215996 223848
rect 222936 223796 222988 223848
rect 233700 223796 233752 223848
rect 239680 223796 239732 223848
rect 241980 223796 242032 223848
rect 285036 223796 285088 223848
rect 126704 223660 126756 223712
rect 131120 223660 131172 223712
rect 132408 223660 132460 223712
rect 201684 223660 201736 223712
rect 87972 223524 88024 223576
rect 81348 223388 81400 223440
rect 157248 223388 157300 223440
rect 157432 223388 157484 223440
rect 159824 223388 159876 223440
rect 161940 223524 161992 223576
rect 167828 223524 167880 223576
rect 168288 223524 168340 223576
rect 226708 223524 226760 223576
rect 269028 223524 269080 223576
rect 298008 223524 298060 223576
rect 300124 223524 300176 223576
rect 426440 223592 426492 223644
rect 426992 223592 427044 223644
rect 306012 223524 306064 223576
rect 329104 223524 329156 223576
rect 342720 223524 342772 223576
rect 457996 223524 458048 223576
rect 460204 223524 460256 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 679256 223524 679308 223576
rect 680176 223524 680228 223576
rect 164976 223388 165028 223440
rect 165252 223388 165304 223440
rect 224040 223388 224092 223440
rect 260104 223388 260156 223440
rect 298928 223388 298980 223440
rect 302148 223388 302200 223440
rect 331128 223388 331180 223440
rect 518900 223388 518952 223440
rect 530032 223388 530084 223440
rect 92112 223252 92164 223304
rect 166816 223252 166868 223304
rect 166954 223252 167006 223304
rect 176108 223252 176160 223304
rect 176292 223252 176344 223304
rect 181444 223252 181496 223304
rect 181628 223252 181680 223304
rect 192024 223252 192076 223304
rect 203892 223252 203944 223304
rect 254860 223252 254912 223304
rect 264796 223252 264848 223304
rect 304724 223252 304776 223304
rect 306288 223252 306340 223304
rect 336924 223252 336976 223304
rect 343548 223252 343600 223304
rect 363972 223252 364024 223304
rect 489552 223252 489604 223304
rect 504364 223252 504416 223304
rect 505100 223252 505152 223304
rect 524236 223252 524288 223304
rect 529020 223252 529072 223304
rect 542452 223252 542504 223304
rect 78588 223116 78640 223168
rect 156880 223116 156932 223168
rect 157064 223116 157116 223168
rect 162124 223116 162176 223168
rect 164148 223116 164200 223168
rect 165252 223116 165304 223168
rect 165804 223116 165856 223168
rect 222292 223116 222344 223168
rect 224224 223116 224276 223168
rect 238392 223116 238444 223168
rect 245292 223116 245344 223168
rect 287612 223116 287664 223168
rect 290832 223116 290884 223168
rect 323676 223116 323728 223168
rect 330484 223116 330536 223168
rect 354956 223116 355008 223168
rect 357072 223116 357124 223168
rect 376208 223116 376260 223168
rect 490196 223116 490248 223168
rect 505652 223116 505704 223168
rect 513104 223116 513156 223168
rect 534172 223116 534224 223168
rect 534724 223116 534776 223168
rect 547420 223116 547472 223168
rect 89444 222980 89496 223032
rect 161940 222980 161992 223032
rect 112812 222844 112864 222896
rect 180892 222980 180944 223032
rect 181444 222980 181496 223032
rect 234804 222980 234856 223032
rect 235172 222980 235224 223032
rect 243268 222980 243320 223032
rect 250904 222980 250956 223032
rect 294420 222980 294472 223032
rect 300308 222980 300360 223032
rect 331772 222980 331824 223032
rect 337936 222980 337988 223032
rect 359188 222980 359240 223032
rect 370504 222980 370556 223032
rect 384580 222980 384632 223032
rect 387708 222980 387760 223032
rect 398104 222980 398156 223032
rect 501144 222980 501196 223032
rect 519268 222980 519320 223032
rect 523684 222980 523736 223032
rect 548064 222980 548116 223032
rect 549260 222980 549312 223032
rect 564808 222980 564860 223032
rect 162308 222844 162360 222896
rect 221648 222844 221700 222896
rect 233148 222844 233200 222896
rect 277676 222844 277728 222896
rect 283380 222844 283432 222896
rect 316960 222844 317012 222896
rect 317144 222844 317196 222896
rect 343364 222844 343416 222896
rect 347596 222844 347648 222896
rect 368480 222844 368532 222896
rect 375104 222844 375156 222896
rect 391020 222844 391072 222896
rect 397368 222844 397420 222896
rect 407120 222844 407172 222896
rect 408408 222844 408460 222896
rect 416872 222844 416924 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 478328 222844 478380 222896
rect 486148 222844 486200 222896
rect 486976 222844 487028 222896
rect 501052 222844 501104 222896
rect 504640 222844 504692 222896
rect 523408 222844 523460 222896
rect 533712 222844 533764 222896
rect 560760 222844 560812 222896
rect 562968 222844 563020 222896
rect 564624 222776 564676 222828
rect 569316 222776 569368 222828
rect 85488 222708 85540 222760
rect 161756 222708 161808 222760
rect 162124 222708 162176 222760
rect 99288 222572 99340 222624
rect 175556 222572 175608 222624
rect 176108 222708 176160 222760
rect 181628 222708 181680 222760
rect 192116 222708 192168 222760
rect 207480 222708 207532 222760
rect 209504 222708 209556 222760
rect 210240 222708 210292 222760
rect 213828 222708 213880 222760
rect 262864 222708 262916 222760
rect 263508 222708 263560 222760
rect 296996 222708 297048 222760
rect 564808 222640 564860 222692
rect 572168 222640 572220 222692
rect 133512 222436 133564 222488
rect 151360 222436 151412 222488
rect 154212 222436 154264 222488
rect 214380 222436 214432 222488
rect 214748 222572 214800 222624
rect 260288 222572 260340 222624
rect 562416 222504 562468 222556
rect 569132 222504 569184 222556
rect 219716 222436 219768 222488
rect 220084 222436 220136 222488
rect 268660 222436 268712 222488
rect 557356 222368 557408 222420
rect 562784 222368 562836 222420
rect 563428 222368 563480 222420
rect 571432 222368 571484 222420
rect 572352 222368 572404 222420
rect 573180 222368 573232 222420
rect 56508 222300 56560 222352
rect 142620 222300 142672 222352
rect 145012 222300 145064 222352
rect 208768 222300 208820 222352
rect 210976 222300 211028 222352
rect 214748 222300 214800 222352
rect 220452 222300 220504 222352
rect 268016 222300 268068 222352
rect 143448 222232 143500 222284
rect 144828 222232 144880 222284
rect 214932 222232 214984 222284
rect 216220 222232 216272 222284
rect 95424 221960 95476 222012
rect 117780 222096 117832 222148
rect 117964 222096 118016 222148
rect 171048 222096 171100 222148
rect 104532 221960 104584 222012
rect 174912 222164 174964 222216
rect 176292 222164 176344 222216
rect 180892 222164 180944 222216
rect 185216 222164 185268 222216
rect 482928 222164 482980 222216
rect 593972 222232 594024 222284
rect 176660 222096 176712 222148
rect 179972 222096 180024 222148
rect 176108 222028 176160 222080
rect 181628 222028 181680 222080
rect 240140 222096 240192 222148
rect 261024 222096 261076 222148
rect 301688 222096 301740 222148
rect 311532 222096 311584 222148
rect 338396 222096 338448 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 553216 222096 553268 222148
rect 558184 222096 558236 222148
rect 558368 222096 558420 222148
rect 562416 222096 562468 222148
rect 562968 222096 563020 222148
rect 567568 222096 567620 222148
rect 567752 222096 567804 222148
rect 572352 222096 572404 222148
rect 572628 222096 572680 222148
rect 71412 221824 71464 221876
rect 142804 221824 142856 221876
rect 142988 221824 143040 221876
rect 172980 221960 173032 222012
rect 176292 221960 176344 222012
rect 181444 221960 181496 222012
rect 185860 221960 185912 222012
rect 237564 221960 237616 222012
rect 243636 221960 243688 222012
rect 285956 221960 286008 222012
rect 309876 221960 309928 222012
rect 338212 221960 338264 222012
rect 500040 221960 500092 222012
rect 518440 221960 518492 222012
rect 525892 221960 525944 222012
rect 597468 221960 597520 222012
rect 340880 221892 340932 221944
rect 341616 221892 341668 221944
rect 171508 221824 171560 221876
rect 229652 221824 229704 221876
rect 230388 221824 230440 221876
rect 258724 221824 258776 221876
rect 267832 221824 267884 221876
rect 273996 221824 274048 221876
rect 285680 221824 285732 221876
rect 286324 221824 286376 221876
rect 304632 221824 304684 221876
rect 334072 221824 334124 221876
rect 515404 221824 515456 221876
rect 535000 221824 535052 221876
rect 542728 221824 542780 221876
rect 543188 221824 543240 221876
rect 600596 221960 600648 222012
rect 600964 222096 601016 222148
rect 607772 222096 607824 222148
rect 601148 221960 601200 222012
rect 597836 221824 597888 221876
rect 607312 221824 607364 221876
rect 68100 221688 68152 221740
rect 147496 221688 147548 221740
rect 147772 221688 147824 221740
rect 61476 221552 61528 221604
rect 137284 221552 137336 221604
rect 137468 221552 137520 221604
rect 64604 221416 64656 221468
rect 138296 221416 138348 221468
rect 138480 221416 138532 221468
rect 142436 221416 142488 221468
rect 142804 221552 142856 221604
rect 147312 221552 147364 221604
rect 161664 221688 161716 221740
rect 224408 221688 224460 221740
rect 227076 221688 227128 221740
rect 272708 221688 272760 221740
rect 204904 221552 204956 221604
rect 205088 221552 205140 221604
rect 142988 221416 143040 221468
rect 148416 221416 148468 221468
rect 211988 221416 212040 221468
rect 214656 221552 214708 221604
rect 258540 221552 258592 221604
rect 258724 221552 258776 221604
rect 275284 221688 275336 221740
rect 278320 221688 278372 221740
rect 313464 221688 313516 221740
rect 331404 221688 331456 221740
rect 353944 221688 353996 221740
rect 359556 221688 359608 221740
rect 376852 221688 376904 221740
rect 484308 221688 484360 221740
rect 496084 221688 496136 221740
rect 503444 221688 503496 221740
rect 521752 221688 521804 221740
rect 522856 221688 522908 221740
rect 546592 221688 546644 221740
rect 547144 221688 547196 221740
rect 275100 221552 275152 221604
rect 310888 221552 310940 221604
rect 314568 221552 314620 221604
rect 340880 221552 340932 221604
rect 341340 221552 341392 221604
rect 361948 221552 362000 221604
rect 377772 221552 377824 221604
rect 390008 221552 390060 221604
rect 456708 221552 456760 221604
rect 462136 221552 462188 221604
rect 496268 221552 496320 221604
rect 513380 221552 513432 221604
rect 529756 221552 529808 221604
rect 555424 221552 555476 221604
rect 556068 221688 556120 221740
rect 562968 221688 563020 221740
rect 563796 221688 563848 221740
rect 567384 221688 567436 221740
rect 567568 221688 567620 221740
rect 556344 221552 556396 221604
rect 556804 221552 556856 221604
rect 567476 221552 567528 221604
rect 567752 221552 567804 221604
rect 568120 221552 568172 221604
rect 597836 221552 597888 221604
rect 601332 221688 601384 221740
rect 606576 221688 606628 221740
rect 610256 221552 610308 221604
rect 655704 221552 655756 221604
rect 659568 221552 659620 221604
rect 232136 221416 232188 221468
rect 241152 221416 241204 221468
rect 285680 221416 285732 221468
rect 285956 221416 286008 221468
rect 289820 221416 289872 221468
rect 290004 221416 290056 221468
rect 321744 221416 321796 221468
rect 338856 221416 338908 221468
rect 117780 221280 117832 221332
rect 107844 221144 107896 221196
rect 117964 221144 118016 221196
rect 118424 221280 118476 221332
rect 177396 221280 177448 221332
rect 178224 221280 178276 221332
rect 181260 221280 181312 221332
rect 181444 221280 181496 221332
rect 195244 221280 195296 221332
rect 195428 221280 195480 221332
rect 245108 221280 245160 221332
rect 258540 221280 258592 221332
rect 265716 221280 265768 221332
rect 273444 221280 273496 221332
rect 309232 221280 309284 221332
rect 362040 221416 362092 221468
rect 379888 221416 379940 221468
rect 391020 221416 391072 221468
rect 400312 221416 400364 221468
rect 405096 221416 405148 221468
rect 414204 221416 414256 221468
rect 452568 221416 452620 221468
rect 456708 221416 456760 221468
rect 483756 221416 483808 221468
rect 538680 221416 538732 221468
rect 550640 221416 550692 221468
rect 600964 221416 601016 221468
rect 601148 221416 601200 221468
rect 610072 221416 610124 221468
rect 654140 221416 654192 221468
rect 655888 221416 655940 221468
rect 362316 221280 362368 221332
rect 548064 221212 548116 221264
rect 567752 221212 567804 221264
rect 567936 221212 567988 221264
rect 568948 221212 569000 221264
rect 569132 221212 569184 221264
rect 608692 221212 608744 221264
rect 137100 221144 137152 221196
rect 137284 221144 137336 221196
rect 144000 221144 144052 221196
rect 144184 221144 144236 221196
rect 203248 221144 203300 221196
rect 117780 221008 117832 221060
rect 187884 221008 187936 221060
rect 188160 221008 188212 221060
rect 195060 221008 195112 221060
rect 195244 221008 195296 221060
rect 205088 221144 205140 221196
rect 206008 221144 206060 221196
rect 258356 221144 258408 221196
rect 542084 221076 542136 221128
rect 549260 221076 549312 221128
rect 550456 221076 550508 221128
rect 554228 221076 554280 221128
rect 558184 221076 558236 221128
rect 608876 221076 608928 221128
rect 204904 221008 204956 221060
rect 211620 221008 211672 221060
rect 211988 221008 212040 221060
rect 214196 221008 214248 221060
rect 237104 221008 237156 221060
rect 280436 221008 280488 221060
rect 415032 221008 415084 221060
rect 420184 221008 420236 221060
rect 545764 220940 545816 220992
rect 601332 220940 601384 220992
rect 108028 220872 108080 220924
rect 97724 220736 97776 220788
rect 114468 220872 114520 220924
rect 118424 220872 118476 220924
rect 128544 220872 128596 220924
rect 198924 220872 198976 220924
rect 203248 220872 203300 220924
rect 206468 220872 206520 220924
rect 256056 220872 256108 220924
rect 261392 220872 261444 220924
rect 420644 220804 420696 220856
rect 423772 220804 423824 220856
rect 466092 220804 466144 220856
rect 471704 220804 471756 220856
rect 518440 220804 518492 220856
rect 600412 220804 600464 220856
rect 600596 220804 600648 220856
rect 606024 220940 606076 220992
rect 137284 220736 137336 220788
rect 137468 220736 137520 220788
rect 197728 220736 197780 220788
rect 198096 220736 198148 220788
rect 252744 220736 252796 220788
rect 253572 220736 253624 220788
rect 293316 220736 293368 220788
rect 296996 220736 297048 220788
rect 310704 220736 310756 220788
rect 311808 220736 311860 220788
rect 327080 220736 327132 220788
rect 329288 220736 329340 220788
rect 331956 220736 332008 220788
rect 414204 220736 414256 220788
rect 418252 220736 418304 220788
rect 455236 220736 455288 220788
rect 458824 220736 458876 220788
rect 475384 220736 475436 220788
rect 476212 220736 476264 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 601976 220736 602028 220788
rect 617248 220736 617300 220788
rect 91284 220600 91336 220652
rect 108028 220600 108080 220652
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 172704 220600 172756 220652
rect 177212 220600 177264 220652
rect 182640 220600 182692 220652
rect 183100 220600 183152 220652
rect 184204 220600 184256 220652
rect 184388 220600 184440 220652
rect 234068 220600 234120 220652
rect 240324 220600 240376 220652
rect 283012 220600 283064 220652
rect 296628 220600 296680 220652
rect 327448 220600 327500 220652
rect 328092 220600 328144 220652
rect 351368 220600 351420 220652
rect 474004 220600 474056 220652
rect 475384 220600 475436 220652
rect 493968 220600 494020 220652
rect 508504 220600 508556 220652
rect 511264 220600 511316 220652
rect 527548 220600 527600 220652
rect 541716 220600 541768 220652
rect 545948 220600 546000 220652
rect 83004 220464 83056 220516
rect 76380 220328 76432 220380
rect 150026 220328 150078 220380
rect 150900 220328 150952 220380
rect 152280 220328 152332 220380
rect 152648 220464 152700 220516
rect 167184 220464 167236 220516
rect 170772 220464 170824 220516
rect 229284 220464 229336 220516
rect 254400 220464 254452 220516
rect 296812 220464 296864 220516
rect 299940 220464 299992 220516
rect 330024 220464 330076 220516
rect 371148 220464 371200 220516
rect 385224 220464 385276 220516
rect 482284 220464 482336 220516
rect 491944 220464 491996 220516
rect 507032 220464 507084 220516
rect 522028 220464 522080 220516
rect 522304 220464 522356 220516
rect 539968 220464 540020 220516
rect 157340 220328 157392 220380
rect 157524 220328 157576 220380
rect 210240 220328 210292 220380
rect 66444 220192 66496 220244
rect 147496 220192 147548 220244
rect 147634 220192 147686 220244
rect 152648 220192 152700 220244
rect 152832 220192 152884 220244
rect 214012 220328 214064 220380
rect 229192 220328 229244 220380
rect 276112 220328 276164 220380
rect 280068 220328 280120 220380
rect 314108 220328 314160 220380
rect 323124 220328 323176 220380
rect 348148 220328 348200 220380
rect 352932 220328 352984 220380
rect 371424 220328 371476 220380
rect 436284 220328 436336 220380
rect 437020 220328 437072 220380
rect 469128 220328 469180 220380
rect 474556 220328 474608 220380
rect 481548 220328 481600 220380
rect 492772 220328 492824 220380
rect 496452 220328 496504 220380
rect 510988 220328 511040 220380
rect 517152 220328 517204 220380
rect 539140 220328 539192 220380
rect 543832 220464 543884 220516
rect 552388 220600 552440 220652
rect 557540 220600 557592 220652
rect 558552 220600 558604 220652
rect 559932 220600 559984 220652
rect 626632 220600 626684 220652
rect 546316 220464 546368 220516
rect 553492 220464 553544 220516
rect 554228 220464 554280 220516
rect 625252 220464 625304 220516
rect 622676 220328 622728 220380
rect 63132 220056 63184 220108
rect 140780 220056 140832 220108
rect 140964 220056 141016 220108
rect 147036 220056 147088 220108
rect 150716 220056 150768 220108
rect 211344 220192 211396 220244
rect 217140 220192 217192 220244
rect 265164 220192 265216 220244
rect 280896 220192 280948 220244
rect 317512 220192 317564 220244
rect 332232 220192 332284 220244
rect 357532 220192 357584 220244
rect 360384 220192 360436 220244
rect 377404 220192 377456 220244
rect 390100 220192 390152 220244
rect 401692 220192 401744 220244
rect 430120 220192 430172 220244
rect 432052 220192 432104 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 472992 220192 473044 220244
rect 482008 220192 482060 220244
rect 488448 220192 488500 220244
rect 502708 220192 502760 220244
rect 504180 220192 504232 220244
rect 515220 220192 515272 220244
rect 515956 220192 516008 220244
rect 521568 220192 521620 220244
rect 543832 220192 543884 220244
rect 544016 220192 544068 220244
rect 559380 220192 559432 220244
rect 559564 220192 559616 220244
rect 563244 220192 563296 220244
rect 566924 220192 566976 220244
rect 571248 220192 571300 220244
rect 571892 220192 571944 220244
rect 628012 220192 628064 220244
rect 563428 220124 563480 220176
rect 566740 220124 566792 220176
rect 211344 220056 211396 220108
rect 263048 220056 263100 220108
rect 263324 220056 263376 220108
rect 301044 220056 301096 220108
rect 318156 220056 318208 220108
rect 343732 220056 343784 220108
rect 345480 220056 345532 220108
rect 367376 220056 367428 220108
rect 367836 220056 367888 220108
rect 382464 220056 382516 220108
rect 382740 220056 382792 220108
rect 394792 220056 394844 220108
rect 397644 220056 397696 220108
rect 405832 220056 405884 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 431960 220056 432012 220108
rect 434812 220056 434864 220108
rect 478512 220056 478564 220108
rect 489460 220056 489512 220108
rect 492312 220056 492364 220108
rect 507676 220056 507728 220108
rect 527824 220056 527876 220108
rect 543694 220056 543746 220108
rect 549996 220056 550048 220108
rect 550456 220056 550508 220108
rect 553492 220056 553544 220108
rect 111248 219920 111300 219972
rect 177212 219920 177264 219972
rect 177396 219920 177448 219972
rect 184388 219920 184440 219972
rect 190644 219920 190696 219972
rect 244464 219920 244516 219972
rect 256884 219920 256936 219972
rect 295892 219920 295944 219972
rect 306748 219920 306800 219972
rect 320364 219920 320416 219972
rect 549444 219988 549496 220040
rect 554964 220056 555016 220108
rect 556068 220056 556120 220108
rect 556344 220056 556396 220108
rect 557356 220056 557408 220108
rect 557540 220056 557592 220108
rect 625436 220056 625488 220108
rect 647240 220056 647292 220108
rect 652760 220056 652812 220108
rect 676036 219988 676088 220040
rect 677048 219988 677100 220040
rect 542268 219852 542320 219904
rect 562692 219920 562744 219972
rect 582380 219920 582432 219972
rect 547604 219852 547656 219904
rect 553676 219852 553728 219904
rect 562876 219852 562928 219904
rect 572076 219852 572128 219904
rect 573180 219852 573232 219904
rect 582196 219852 582248 219904
rect 626816 219852 626868 219904
rect 124404 219784 124456 219836
rect 193496 219784 193548 219836
rect 197268 219784 197320 219836
rect 249892 219784 249944 219836
rect 293592 219784 293644 219836
rect 299756 219784 299808 219836
rect 522028 219716 522080 219768
rect 522580 219716 522632 219768
rect 531320 219716 531372 219768
rect 532516 219716 532568 219768
rect 621020 219716 621072 219768
rect 676036 219716 676088 219768
rect 677416 219716 677468 219768
rect 131028 219648 131080 219700
rect 137284 219648 137336 219700
rect 147496 219648 147548 219700
rect 148048 219648 148100 219700
rect 205824 219648 205876 219700
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 668400 219648 668452 219700
rect 669320 219648 669372 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 520188 219580 520240 219632
rect 105820 219444 105872 219496
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 72240 219376 72292 219428
rect 73160 219376 73212 219428
rect 80520 219376 80572 219428
rect 90272 219376 90324 219428
rect 90456 219376 90508 219428
rect 106924 219240 106976 219292
rect 117964 219376 118016 219428
rect 119252 219376 119304 219428
rect 119436 219376 119488 219428
rect 119988 219376 120040 219428
rect 126060 219376 126112 219428
rect 126888 219376 126940 219428
rect 127716 219376 127768 219428
rect 128268 219376 128320 219428
rect 130200 219376 130252 219428
rect 132684 219376 132736 219428
rect 133788 219376 133840 219428
rect 137468 219512 137520 219564
rect 137652 219512 137704 219564
rect 203432 219512 203484 219564
rect 210240 219512 210292 219564
rect 218612 219512 218664 219564
rect 270776 219512 270828 219564
rect 279240 219512 279292 219564
rect 515956 219512 516008 219564
rect 618260 219580 618312 219632
rect 221648 219444 221700 219496
rect 142436 219376 142488 219428
rect 142620 219376 142672 219428
rect 143172 219376 143224 219428
rect 143632 219376 143684 219428
rect 197912 219376 197964 219428
rect 199752 219376 199804 219428
rect 204720 219376 204772 219428
rect 208860 219376 208912 219428
rect 209780 219376 209832 219428
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 232504 219376 232556 219428
rect 233700 219376 233752 219428
rect 234620 219376 234672 219428
rect 152372 219240 152424 219292
rect 152556 219240 152608 219292
rect 153108 219240 153160 219292
rect 153384 219240 153436 219292
rect 158996 219240 159048 219292
rect 159180 219240 159232 219292
rect 160008 219240 160060 219292
rect 160192 219240 160244 219292
rect 163964 219240 164016 219292
rect 164976 219240 165028 219292
rect 165436 219240 165488 219292
rect 165804 219240 165856 219292
rect 166540 219240 166592 219292
rect 85304 219104 85356 219156
rect 117964 219104 118016 219156
rect 119252 219104 119304 219156
rect 123392 219104 123444 219156
rect 123576 219104 123628 219156
rect 128728 219104 128780 219156
rect 131856 219104 131908 219156
rect 132408 219104 132460 219156
rect 70584 218968 70636 219020
rect 134432 218968 134484 219020
rect 135076 218968 135128 219020
rect 135996 218968 136048 219020
rect 136548 218968 136600 219020
rect 136824 218968 136876 219020
rect 137836 218968 137888 219020
rect 138112 219104 138164 219156
rect 143632 219104 143684 219156
rect 143816 219104 143868 219156
rect 152280 219104 152332 219156
rect 168932 219240 168984 219292
rect 169300 219240 169352 219292
rect 139952 218968 140004 219020
rect 140136 218968 140188 219020
rect 142252 218968 142304 219020
rect 142436 218968 142488 219020
rect 167000 219104 167052 219156
rect 190092 219104 190144 219156
rect 193128 219240 193180 219292
rect 195428 219240 195480 219292
rect 196072 219240 196124 219292
rect 199384 219240 199436 219292
rect 195060 219104 195112 219156
rect 195244 219104 195296 219156
rect 226892 219240 226944 219292
rect 232872 219240 232924 219292
rect 237840 219240 237892 219292
rect 239404 219240 239456 219292
rect 246120 219376 246172 219428
rect 285956 219376 286008 219428
rect 287520 219376 287572 219428
rect 288440 219376 288492 219428
rect 291660 219376 291712 219428
rect 324688 219376 324740 219428
rect 325608 219376 325660 219428
rect 326344 219376 326396 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 352104 219376 352156 219428
rect 366364 219376 366416 219428
rect 374460 219376 374512 219428
rect 375380 219376 375432 219428
rect 380256 219376 380308 219428
rect 384304 219376 384356 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 403440 219376 403492 219428
rect 404360 219376 404412 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 557724 219444 557776 219496
rect 558736 219444 558788 219496
rect 438216 219376 438268 219428
rect 438860 219376 438912 219428
rect 439872 219376 439924 219428
rect 440332 219376 440384 219428
rect 488724 219376 488776 219428
rect 489184 219376 489236 219428
rect 518808 219376 518860 219428
rect 519820 219376 519872 219428
rect 504640 219308 504692 219360
rect 505284 219308 505336 219360
rect 540244 219308 540296 219360
rect 540796 219308 540848 219360
rect 542268 219308 542320 219360
rect 542452 219308 542504 219360
rect 555608 219308 555660 219360
rect 555792 219308 555844 219360
rect 571984 219308 572036 219360
rect 573824 219308 573876 219360
rect 575296 219308 575348 219360
rect 582196 219308 582248 219360
rect 599032 219308 599084 219360
rect 601792 219444 601844 219496
rect 628196 219444 628248 219496
rect 676220 219376 676272 219428
rect 677600 219376 677652 219428
rect 601976 219308 602028 219360
rect 270776 219240 270828 219292
rect 327264 219240 327316 219292
rect 152740 218968 152792 219020
rect 166264 218968 166316 219020
rect 167184 218968 167236 219020
rect 200580 218968 200632 219020
rect 201500 218968 201552 219020
rect 204720 219104 204772 219156
rect 246304 219104 246356 219156
rect 258540 219104 258592 219156
rect 259276 219104 259328 219156
rect 259460 219104 259512 219156
rect 291844 219104 291896 219156
rect 294144 219104 294196 219156
rect 311808 219104 311860 219156
rect 315672 219104 315724 219156
rect 317972 219104 318024 219156
rect 320640 219104 320692 219156
rect 340144 219104 340196 219156
rect 383568 219240 383620 219292
rect 387064 219240 387116 219292
rect 450728 219240 450780 219292
rect 453856 219240 453908 219292
rect 479708 219240 479760 219292
rect 480352 219240 480404 219292
rect 534172 219240 534224 219292
rect 534632 219240 534684 219292
rect 544936 219172 544988 219224
rect 553492 219172 553544 219224
rect 345664 219104 345716 219156
rect 204904 218968 204956 219020
rect 206376 218968 206428 219020
rect 255872 218968 255924 219020
rect 259276 218968 259328 219020
rect 293592 218968 293644 219020
rect 300768 218968 300820 219020
rect 329288 218968 329340 219020
rect 333704 218968 333756 219020
rect 352564 219104 352616 219156
rect 354404 219104 354456 219156
rect 355508 219104 355560 219156
rect 358728 219104 358780 219156
rect 364984 219104 365036 219156
rect 419172 219104 419224 219156
rect 422668 219104 422720 219156
rect 483572 219104 483624 219156
rect 490288 219104 490340 219156
rect 503076 219104 503128 219156
rect 503536 219104 503588 219156
rect 507124 219104 507176 219156
rect 514944 219104 514996 219156
rect 535184 219104 535236 219156
rect 544016 219104 544068 219156
rect 544476 219036 544528 219088
rect 351368 218968 351420 219020
rect 355232 218968 355284 219020
rect 355416 218968 355468 219020
rect 369124 218968 369176 219020
rect 373632 218968 373684 219020
rect 380072 218968 380124 219020
rect 384396 218968 384448 219020
rect 393964 218968 394016 219020
rect 401784 218968 401836 219020
rect 407764 218968 407816 219020
rect 514760 218968 514812 219020
rect 519820 218968 519872 219020
rect 524420 218968 524472 219020
rect 544200 218968 544252 219020
rect 558276 219104 558328 219156
rect 558736 219104 558788 219156
rect 566556 219172 566608 219224
rect 567844 219172 567896 219224
rect 573272 219172 573324 219224
rect 573456 219172 573508 219224
rect 582288 219172 582340 219224
rect 567016 219104 567068 219156
rect 553860 218968 553912 219020
rect 555240 218968 555292 219020
rect 555608 218968 555660 219020
rect 62304 218832 62356 218884
rect 76564 218832 76616 218884
rect 83832 218832 83884 218884
rect 152096 218832 152148 218884
rect 152280 218832 152332 218884
rect 166448 218832 166500 218884
rect 167184 218832 167236 218884
rect 215944 218832 215996 218884
rect 217968 218832 218020 218884
rect 220084 218832 220136 218884
rect 77208 218696 77260 218748
rect 147496 218696 147548 218748
rect 59820 218560 59872 218612
rect 69572 218560 69624 218612
rect 92940 218560 92992 218612
rect 93768 218560 93820 218612
rect 93768 218424 93820 218476
rect 139952 218560 140004 218612
rect 140136 218560 140188 218612
rect 143816 218560 143868 218612
rect 144276 218560 144328 218612
rect 144828 218560 144880 218612
rect 146760 218560 146812 218612
rect 152740 218696 152792 218748
rect 152924 218696 152976 218748
rect 156328 218696 156380 218748
rect 156696 218696 156748 218748
rect 162124 218696 162176 218748
rect 149060 218560 149112 218612
rect 157984 218560 158036 218612
rect 158996 218560 159048 218612
rect 166264 218696 166316 218748
rect 167368 218696 167420 218748
rect 213184 218696 213236 218748
rect 213552 218696 213604 218748
rect 217324 218696 217376 218748
rect 218796 218696 218848 218748
rect 219348 218696 219400 218748
rect 219624 218696 219676 218748
rect 221096 218696 221148 218748
rect 224224 218696 224276 218748
rect 225972 218832 226024 218884
rect 264152 218696 264204 218748
rect 162676 218560 162728 218612
rect 166540 218560 166592 218612
rect 169944 218560 169996 218612
rect 181076 218560 181128 218612
rect 182364 218560 182416 218612
rect 183284 218560 183336 218612
rect 113640 218424 113692 218476
rect 119988 218424 120040 218476
rect 128728 218424 128780 218476
rect 174544 218424 174596 218476
rect 174728 218424 174780 218476
rect 195244 218560 195296 218612
rect 195428 218560 195480 218612
rect 243452 218560 243504 218612
rect 252744 218560 252796 218612
rect 259460 218560 259512 218612
rect 274272 218832 274324 218884
rect 280712 218832 280764 218884
rect 281080 218832 281132 218884
rect 312544 218832 312596 218884
rect 314016 218832 314068 218884
rect 329104 218832 329156 218884
rect 337200 218832 337252 218884
rect 357716 218832 357768 218884
rect 366732 218832 366784 218884
rect 378784 218832 378836 218884
rect 386052 218832 386104 218884
rect 396632 218832 396684 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412456 218832 412508 218884
rect 505836 218832 505888 218884
rect 265992 218696 266044 218748
rect 302884 218696 302936 218748
rect 307392 218696 307444 218748
rect 337016 218696 337068 218748
rect 340512 218696 340564 218748
rect 360844 218696 360896 218748
rect 379152 218696 379204 218748
rect 392124 218696 392176 218748
rect 395804 218696 395856 218748
rect 404544 218696 404596 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 460204 218696 460256 218748
rect 461308 218696 461360 218748
rect 502524 218628 502576 218680
rect 505008 218628 505060 218680
rect 267832 218560 267884 218612
rect 272616 218560 272668 218612
rect 296996 218560 297048 218612
rect 429936 218560 429988 218612
rect 432696 218560 432748 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 518808 218696 518860 218748
rect 519544 218832 519596 218884
rect 526444 218832 526496 218884
rect 533436 218832 533488 218884
rect 533896 218832 533948 218884
rect 537576 218832 537628 218884
rect 524604 218696 524656 218748
rect 525064 218696 525116 218748
rect 529388 218696 529440 218748
rect 533620 218696 533672 218748
rect 534356 218696 534408 218748
rect 535000 218696 535052 218748
rect 547972 218696 548024 218748
rect 549076 218832 549128 218884
rect 556160 218832 556212 218884
rect 567200 218968 567252 219020
rect 572260 219036 572312 219088
rect 574560 219036 574612 219088
rect 571800 218968 571852 219020
rect 574744 218968 574796 219020
rect 586520 218968 586572 219020
rect 559748 218832 559800 218884
rect 567844 218832 567896 218884
rect 568028 218832 568080 218884
rect 572904 218900 572956 218952
rect 573088 218832 573140 218884
rect 591672 218832 591724 218884
rect 186504 218424 186556 218476
rect 235172 218424 235224 218476
rect 239496 218424 239548 218476
rect 272432 218424 272484 218476
rect 279240 218424 279292 218476
rect 281080 218424 281132 218476
rect 285864 218424 285916 218476
rect 306748 218424 306800 218476
rect 482928 218424 482980 218476
rect 485320 218424 485372 218476
rect 501052 218424 501104 218476
rect 510344 218424 510396 218476
rect 544476 218560 544528 218612
rect 548708 218696 548760 218748
rect 555792 218696 555844 218748
rect 556160 218560 556212 218612
rect 558552 218560 558604 218612
rect 559104 218696 559156 218748
rect 562876 218696 562928 218748
rect 563060 218696 563112 218748
rect 572076 218696 572128 218748
rect 572444 218696 572496 218748
rect 575112 218696 575164 218748
rect 582196 218696 582248 218748
rect 586336 218696 586388 218748
rect 562876 218560 562928 218612
rect 527548 218424 527600 218476
rect 567016 218560 567068 218612
rect 567200 218560 567252 218612
rect 563520 218424 563572 218476
rect 597468 218560 597520 218612
rect 75552 218288 75604 218340
rect 83464 218288 83516 218340
rect 100392 218288 100444 218340
rect 105820 218288 105872 218340
rect 107016 218288 107068 218340
rect 149060 218288 149112 218340
rect 149244 218288 149296 218340
rect 150348 218288 150400 218340
rect 150532 218288 150584 218340
rect 157248 218288 157300 218340
rect 56324 218152 56376 218204
rect 62764 218152 62816 218204
rect 79692 218152 79744 218204
rect 82084 218152 82136 218204
rect 119988 218152 120040 218204
rect 159824 218288 159876 218340
rect 160008 218288 160060 218340
rect 162676 218288 162728 218340
rect 162860 218288 162912 218340
rect 166448 218288 166500 218340
rect 166632 218288 166684 218340
rect 213552 218288 213604 218340
rect 216312 218288 216364 218340
rect 221648 218288 221700 218340
rect 224592 218288 224644 218340
rect 225604 218288 225656 218340
rect 227904 218288 227956 218340
rect 229192 218288 229244 218340
rect 244464 218288 244516 218340
rect 247684 218288 247736 218340
rect 365352 218288 365404 218340
rect 373264 218288 373316 218340
rect 426624 218288 426676 218340
rect 429568 218288 429620 218340
rect 475568 218288 475620 218340
rect 482836 218288 482888 218340
rect 500040 218288 500092 218340
rect 507124 218288 507176 218340
rect 507676 218288 507728 218340
rect 157708 218152 157760 218204
rect 161296 218152 161348 218204
rect 162124 218152 162176 218204
rect 167644 218152 167696 218204
rect 168104 218152 168156 218204
rect 171048 218152 171100 218204
rect 171600 218152 171652 218204
rect 55680 218016 55732 218068
rect 56508 218016 56560 218068
rect 57336 218016 57388 218068
rect 57888 218016 57940 218068
rect 58164 218016 58216 218068
rect 61292 218016 61344 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 73896 218016 73948 218068
rect 74448 218016 74500 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 82728 218016 82780 218068
rect 84660 218016 84712 218068
rect 85488 218016 85540 218068
rect 86316 218016 86368 218068
rect 86868 218016 86920 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 94596 218016 94648 218068
rect 95148 218016 95200 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 101220 218016 101272 218068
rect 102140 218016 102192 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 103704 218016 103756 218068
rect 104808 218016 104860 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 110328 218016 110380 218068
rect 110972 218016 111024 218068
rect 111984 218016 112036 218068
rect 112812 218016 112864 218068
rect 115296 218016 115348 218068
rect 115756 218016 115808 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 120264 218016 120316 218068
rect 162860 218016 162912 218068
rect 163320 218016 163372 218068
rect 167460 218016 167512 218068
rect 168288 218016 168340 218068
rect 169116 218016 169168 218068
rect 169576 218016 169628 218068
rect 173256 218016 173308 218068
rect 169300 217880 169352 217932
rect 174084 218016 174136 218068
rect 175188 218016 175240 218068
rect 175740 218152 175792 218204
rect 176476 218152 176528 218204
rect 179880 218152 179932 218204
rect 221096 218152 221148 218204
rect 221280 218152 221332 218204
rect 221832 218152 221884 218204
rect 222936 218152 222988 218204
rect 223396 218152 223448 218204
rect 223764 218152 223816 218204
rect 224868 218152 224920 218204
rect 225420 218152 225472 218204
rect 226156 218152 226208 218204
rect 229560 218152 229612 218204
rect 231032 218152 231084 218204
rect 231216 218152 231268 218204
rect 231676 218152 231728 218204
rect 232044 218152 232096 218204
rect 233148 218152 233200 218204
rect 235356 218152 235408 218204
rect 235908 218152 235960 218204
rect 236184 218152 236236 218204
rect 236920 218152 236972 218204
rect 176292 218016 176344 218068
rect 176568 218016 176620 218068
rect 177580 218016 177632 218068
rect 189816 218016 189868 218068
rect 190276 218016 190328 218068
rect 174728 217880 174780 217932
rect 190092 217880 190144 217932
rect 192116 218016 192168 218068
rect 192300 218016 192352 218068
rect 192944 218016 192996 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 196440 218016 196492 218068
rect 197084 218016 197136 218068
rect 198924 218016 198976 218068
rect 200028 218016 200080 218068
rect 202236 218016 202288 218068
rect 202696 218016 202748 218068
rect 203064 218016 203116 218068
rect 203708 218016 203760 218068
rect 204720 218016 204772 218068
rect 206008 218016 206060 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 213000 218016 213052 218068
rect 215484 218016 215536 218068
rect 216496 218016 216548 218068
rect 249064 218152 249116 218204
rect 249432 218152 249484 218204
rect 251732 218152 251784 218204
rect 269304 218152 269356 218204
rect 273904 218152 273956 218204
rect 299112 218152 299164 218204
rect 300308 218152 300360 218204
rect 302424 218152 302476 218204
rect 304632 218152 304684 218204
rect 310704 218152 310756 218204
rect 315304 218152 315356 218204
rect 330668 218152 330720 218204
rect 333244 218152 333296 218204
rect 348792 218152 348844 218204
rect 351184 218152 351236 218204
rect 364524 218152 364576 218204
rect 367652 218152 367704 218204
rect 369492 218152 369544 218204
rect 370504 218152 370556 218204
rect 376944 218152 376996 218204
rect 382924 218152 382976 218204
rect 386880 218152 386932 218204
rect 388444 218152 388496 218204
rect 394332 218152 394384 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 427912 218152 427964 218204
rect 428464 218152 428516 218204
rect 430120 218152 430172 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 435732 218152 435784 218204
rect 436652 218152 436704 218204
rect 455052 218152 455104 218204
rect 460480 218152 460532 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 494612 218152 494664 218204
rect 495256 218152 495308 218204
rect 519544 218152 519596 218204
rect 519820 218152 519872 218204
rect 524420 218152 524472 218204
rect 529388 218288 529440 218340
rect 571892 218288 571944 218340
rect 573456 218424 573508 218476
rect 573640 218424 573692 218476
rect 606484 218424 606536 218476
rect 573272 218288 573324 218340
rect 574376 218288 574428 218340
rect 574560 218288 574612 218340
rect 605288 218288 605340 218340
rect 548708 218152 548760 218204
rect 548892 218152 548944 218204
rect 553492 218152 553544 218204
rect 553676 218152 553728 218204
rect 563336 218152 563388 218204
rect 571984 218152 572036 218204
rect 572168 218152 572220 218204
rect 574928 218152 574980 218204
rect 586336 218152 586388 218204
rect 594984 218152 595036 218204
rect 596916 218152 596968 218204
rect 601332 218152 601384 218204
rect 563014 218084 563066 218136
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249708 218016 249760 218068
rect 250260 218016 250312 218068
rect 251180 218016 251232 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 262680 218016 262732 218068
rect 263600 218016 263652 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 266820 218016 266872 218068
rect 267694 218016 267746 218068
rect 268476 218016 268528 218068
rect 269028 218016 269080 218068
rect 270960 218016 271012 218068
rect 271604 218016 271656 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278504 218016 278556 218068
rect 281724 218016 281776 218068
rect 282552 218016 282604 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 289176 218016 289228 218068
rect 289636 218016 289688 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 295800 218016 295852 218068
rect 296444 218016 296496 218068
rect 297456 218016 297508 218068
rect 298008 218016 298060 218068
rect 298284 218016 298336 218068
rect 299296 218016 299348 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 304080 218016 304132 218068
rect 305552 218016 305604 218068
rect 305736 218016 305788 218068
rect 306288 218016 306340 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 308220 218016 308272 218068
rect 308772 218016 308824 218068
rect 312360 218016 312412 218068
rect 314568 218016 314620 218068
rect 314844 218016 314896 218068
rect 315856 218016 315908 218068
rect 316500 218016 316552 218068
rect 317144 218016 317196 218068
rect 318984 218016 319036 218068
rect 319996 218016 320048 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 328920 218016 328972 218068
rect 330484 218016 330536 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335268 218016 335320 218068
rect 335544 218016 335596 218068
rect 336372 218016 336424 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 342996 218016 343048 218068
rect 343548 218016 343600 218068
rect 347136 218016 347188 218068
rect 347596 218016 347648 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 353760 218016 353812 218068
rect 354588 218016 354640 218068
rect 356244 218016 356296 218068
rect 357348 218016 357400 218068
rect 357900 218016 357952 218068
rect 359372 218016 359424 218068
rect 363696 218016 363748 218068
rect 364156 218016 364208 218068
rect 366180 218016 366232 218068
rect 366916 218016 366968 218068
rect 368664 218016 368716 218068
rect 369768 218016 369820 218068
rect 370320 218016 370372 218068
rect 370964 218016 371016 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373816 218016 373868 218068
rect 376116 218016 376168 218068
rect 376576 218016 376628 218068
rect 378600 218016 378652 218068
rect 379336 218016 379388 218068
rect 381084 218016 381136 218068
rect 381728 218016 381780 218068
rect 385224 218016 385276 218068
rect 386328 218016 386380 218068
rect 388536 218016 388588 218068
rect 389088 218016 389140 218068
rect 389364 218016 389416 218068
rect 390284 218016 390336 218068
rect 392676 218016 392728 218068
rect 393228 218016 393280 218068
rect 393504 218016 393556 218068
rect 394608 218016 394660 218068
rect 395160 218016 395212 218068
rect 395988 218016 396040 218068
rect 396816 218016 396868 218068
rect 397368 218016 397420 218068
rect 400956 218016 401008 218068
rect 401416 218016 401468 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 418344 218016 418396 218068
rect 419448 218016 419500 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 428280 218016 428332 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 434904 218016 434956 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437756 218016 437808 218068
rect 453304 218016 453356 218068
rect 455512 218016 455564 218068
rect 456708 218016 456760 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 471704 218016 471756 218068
rect 472900 218016 472952 218068
rect 488724 218016 488776 218068
rect 497556 218016 497608 218068
rect 505284 218016 505336 218068
rect 505652 218016 505704 218068
rect 613844 218016 613896 218068
rect 528376 217812 528428 217864
rect 602896 217812 602948 217864
rect 604092 217812 604144 217864
rect 612280 217812 612332 217864
rect 524604 217676 524656 217728
rect 523408 217472 523460 217524
rect 533620 217540 533672 217592
rect 534356 217676 534408 217728
rect 542084 217676 542136 217728
rect 542268 217676 542320 217728
rect 548432 217676 548484 217728
rect 535184 217540 535236 217592
rect 535920 217540 535972 217592
rect 538864 217540 538916 217592
rect 543004 217540 543056 217592
rect 596916 217676 596968 217728
rect 597100 217676 597152 217728
rect 604460 217676 604512 217728
rect 605288 217676 605340 217728
rect 615684 217676 615736 217728
rect 549444 217540 549496 217592
rect 562048 217540 562100 217592
rect 562508 217540 562560 217592
rect 609060 217540 609112 217592
rect 542268 217404 542320 217456
rect 543280 217404 543332 217456
rect 548800 217404 548852 217456
rect 566188 217404 566240 217456
rect 567016 217404 567068 217456
rect 597100 217404 597152 217456
rect 544016 217336 544068 217388
rect 533436 217268 533488 217320
rect 543188 217268 543240 217320
rect 565268 217268 565320 217320
rect 565820 217268 565872 217320
rect 597100 217268 597152 217320
rect 145058 217200 145110 217252
rect 147772 217200 147824 217252
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 543832 217200 543884 217252
rect 530906 217132 530958 217184
rect 541900 217132 541952 217184
rect 147542 217064 147594 217116
rect 150716 217064 150768 217116
rect 520970 217064 521022 217116
rect 543464 217132 543516 217184
rect 544660 217132 544712 217184
rect 564624 217132 564676 217184
rect 566004 217132 566056 217184
rect 567200 217132 567252 217184
rect 569316 217132 569368 217184
rect 603448 217404 603500 217456
rect 597468 217268 597520 217320
rect 601148 217268 601200 217320
rect 601332 217268 601384 217320
rect 605104 217268 605156 217320
rect 606484 217268 606536 217320
rect 616144 217268 616196 217320
rect 598848 217132 598900 217184
rect 614120 217132 614172 217184
rect 566188 217064 566240 217116
rect 567016 217064 567068 217116
rect 574284 216860 574336 216912
rect 574928 216860 574980 216912
rect 590844 216860 590896 216912
rect 594800 216860 594852 216912
rect 594984 216860 595036 216912
rect 598848 216860 598900 216912
rect 601148 216996 601200 217048
rect 623320 216996 623372 217048
rect 605840 216860 605892 216912
rect 574560 216724 574612 216776
rect 575664 216724 575716 216776
rect 590844 216724 590896 216776
rect 592040 216724 592092 216776
rect 595628 216724 595680 216776
rect 596272 216724 596324 216776
rect 597100 216724 597152 216776
rect 604000 216724 604052 216776
rect 574192 216588 574244 216640
rect 576124 216588 576176 216640
rect 576860 216452 576912 216504
rect 586704 216452 586756 216504
rect 595996 216384 596048 216436
rect 596824 216384 596876 216436
rect 599768 215908 599820 215960
rect 613384 215908 613436 215960
rect 582104 215840 582156 215892
rect 595996 215840 596048 215892
rect 613844 215364 613896 215416
rect 615040 215364 615092 215416
rect 636660 215296 636712 215348
rect 639604 215296 639656 215348
rect 574744 215228 574796 215280
rect 621664 215228 621716 215280
rect 574284 215092 574336 215144
rect 619640 215092 619692 215144
rect 675852 215092 675904 215144
rect 677232 215092 677284 215144
rect 577688 214956 577740 215008
rect 626080 214956 626132 215008
rect 663524 214888 663576 214940
rect 664444 214888 664496 214940
rect 575112 214820 575164 214872
rect 622400 214820 622452 214872
rect 575664 214684 575716 214736
rect 616696 214684 616748 214736
rect 616880 214684 616932 214736
rect 617800 214684 617852 214736
rect 624424 214684 624476 214736
rect 633808 214684 633860 214736
rect 575940 214548 575992 214600
rect 576124 214412 576176 214464
rect 620008 214412 620060 214464
rect 626632 214548 626684 214600
rect 627184 214548 627236 214600
rect 630772 214548 630824 214600
rect 631600 214548 631652 214600
rect 662052 214548 662104 214600
rect 663248 214548 663300 214600
rect 628288 214412 628340 214464
rect 658740 214344 658792 214396
rect 661684 214344 661736 214396
rect 600412 214276 600464 214328
rect 600780 214276 600832 214328
rect 608692 214276 608744 214328
rect 609520 214276 609572 214328
rect 616696 214276 616748 214328
rect 624424 214276 624476 214328
rect 35808 213936 35860 213988
rect 40684 213936 40736 213988
rect 626448 213868 626500 213920
rect 629392 213868 629444 213920
rect 638316 213868 638368 213920
rect 640064 213868 640116 213920
rect 648528 213868 648580 213920
rect 650644 213868 650696 213920
rect 655704 213868 655756 213920
rect 656808 213868 656860 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 645492 213732 645544 213784
rect 651196 213732 651248 213784
rect 660948 213732 661000 213784
rect 662972 213732 663024 213784
rect 575296 213596 575348 213648
rect 601792 213596 601844 213648
rect 652024 213596 652076 213648
rect 658004 213596 658056 213648
rect 659568 213596 659620 213648
rect 664628 213596 664680 213648
rect 575480 213460 575532 213512
rect 601240 213460 601292 213512
rect 639972 213460 640024 213512
rect 642088 213460 642140 213512
rect 650460 213460 650512 213512
rect 658924 213460 658976 213512
rect 576308 213324 576360 213376
rect 612832 213324 612884 213376
rect 641628 213324 641680 213376
rect 654784 213324 654836 213376
rect 574928 213188 574980 213240
rect 623872 213188 623924 213240
rect 635556 213188 635608 213240
rect 651840 213188 651892 213240
rect 652852 213188 652904 213240
rect 660212 213188 660264 213240
rect 675852 213188 675904 213240
rect 676680 213188 676732 213240
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 632704 212848 632756 212900
rect 634360 212848 634412 212900
rect 628656 212712 628708 212764
rect 632704 212712 632756 212764
rect 637212 212712 637264 212764
rect 641444 212712 641496 212764
rect 35808 211148 35860 211200
rect 41696 211148 41748 211200
rect 610072 210264 610124 210316
rect 610624 210264 610676 210316
rect 578792 209856 578844 209908
rect 581000 209856 581052 209908
rect 591304 208632 591356 208684
rect 632152 209516 632204 209568
rect 652208 209516 652260 209568
rect 667020 209040 667072 209092
rect 35808 208360 35860 208412
rect 40040 208360 40092 208412
rect 578608 208292 578660 208344
rect 589464 208292 589516 208344
rect 579620 207612 579672 207664
rect 589464 207612 589516 207664
rect 581000 206252 581052 206304
rect 589648 206252 589700 206304
rect 578240 205776 578292 205828
rect 581000 205776 581052 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 669320 199044 669372 199096
rect 670792 199044 670844 199096
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 45468 196596 45520 196648
rect 48780 196596 48832 196648
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 669412 194148 669464 194200
rect 670792 194148 670844 194200
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 667940 189252 667992 189304
rect 670792 189252 670844 189304
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 583024 175244 583076 175296
rect 589464 175312 589516 175364
rect 667940 174564 667992 174616
rect 669780 174564 669832 174616
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 581644 171096 581696 171148
rect 589464 171096 589516 171148
rect 579528 170960 579580 171012
rect 583024 170960 583076 171012
rect 582380 169736 582432 169788
rect 589464 169736 589516 169788
rect 578332 169668 578384 169720
rect 580908 169668 580960 169720
rect 668032 169668 668084 169720
rect 670332 169668 670384 169720
rect 579620 168376 579672 168428
rect 589464 168376 589516 168428
rect 578976 167152 579028 167204
rect 581644 167152 581696 167204
rect 581644 167016 581696 167068
rect 589464 167016 589516 167068
rect 578884 165520 578936 165572
rect 582380 165520 582432 165572
rect 667940 164772 667992 164824
rect 670148 164772 670200 164824
rect 585968 164228 586020 164280
rect 589464 164228 589516 164280
rect 584404 162868 584456 162920
rect 589464 162868 589516 162920
rect 676128 162800 676180 162852
rect 678244 162800 678296 162852
rect 675944 162596 675996 162648
rect 679624 162596 679676 162648
rect 675852 161712 675904 161764
rect 681004 161712 681056 161764
rect 580264 161440 580316 161492
rect 589464 161440 589516 161492
rect 582380 160080 582432 160132
rect 589464 160080 589516 160132
rect 579252 160012 579304 160064
rect 581644 160012 581696 160064
rect 581828 158788 581880 158840
rect 589464 158788 589516 158840
rect 579160 158652 579212 158704
rect 585968 158652 586020 158704
rect 585784 157360 585836 157412
rect 589464 157360 589516 157412
rect 579528 155864 579580 155916
rect 584404 155864 584456 155916
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 578240 154504 578292 154556
rect 580264 154504 580316 154556
rect 580448 153212 580500 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 582380 152736 582432 152788
rect 583024 151784 583076 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 581828 150560 581880 150612
rect 581644 150424 581696 150476
rect 589464 150424 589516 150476
rect 579528 147364 579580 147416
rect 585784 147364 585836 147416
rect 587348 146276 587400 146328
rect 589372 146276 589424 146328
rect 668492 146004 668544 146056
rect 670792 146004 670844 146056
rect 578884 145528 578936 145580
rect 589188 145528 589240 145580
rect 585784 144916 585836 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 578608 143148 578660 143200
rect 580448 143148 580500 143200
rect 580264 142128 580316 142180
rect 589464 142128 589516 142180
rect 579528 140564 579580 140616
rect 583024 140564 583076 140616
rect 584404 139408 584456 139460
rect 589464 139408 589516 139460
rect 578700 139340 578752 139392
rect 581644 139340 581696 139392
rect 581644 136620 581696 136672
rect 589464 136620 589516 136672
rect 668032 136280 668084 136332
rect 669964 136280 670016 136332
rect 578332 135872 578384 135924
rect 587348 135872 587400 135924
rect 587164 135260 587216 135312
rect 589280 135260 589332 135312
rect 578240 134240 578292 134292
rect 585784 134240 585836 134292
rect 585968 133900 586020 133952
rect 589464 133900 589516 133952
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 579252 133152 579304 133204
rect 589096 133152 589148 133204
rect 582380 131724 582432 131776
rect 589924 131724 589976 131776
rect 579528 129684 579580 129736
rect 582380 129684 582432 129736
rect 583024 128324 583076 128376
rect 589464 128324 589516 128376
rect 578332 128256 578384 128308
rect 580264 128256 580316 128308
rect 580448 126964 580500 127016
rect 589464 126964 589516 127016
rect 668216 125128 668268 125180
rect 669780 125128 669832 125180
rect 585784 124176 585836 124228
rect 589464 124176 589516 124228
rect 579252 124108 579304 124160
rect 584404 124108 584456 124160
rect 579252 122816 579304 122868
rect 589464 122816 589516 122868
rect 584404 121456 584456 121508
rect 589464 121456 589516 121508
rect 579068 121116 579120 121168
rect 581644 121116 581696 121168
rect 582012 120708 582064 120760
rect 590108 120708 590160 120760
rect 578516 118600 578568 118652
rect 587164 118600 587216 118652
rect 668032 117648 668084 117700
rect 670332 117648 670384 117700
rect 675852 117240 675904 117292
rect 682384 117240 682436 117292
rect 579528 116900 579580 116952
rect 585968 116900 586020 116952
rect 587808 115948 587860 116000
rect 589464 115948 589516 116000
rect 585140 115336 585192 115388
rect 590292 115336 590344 115388
rect 579068 115200 579120 115252
rect 587808 115200 587860 115252
rect 587164 114520 587216 114572
rect 589648 114520 589700 114572
rect 579528 114384 579580 114436
rect 591304 114384 591356 114436
rect 668216 114248 668268 114300
rect 669596 114248 669648 114300
rect 579528 113092 579580 113144
rect 588544 113092 588596 113144
rect 588544 110440 588596 110492
rect 589648 110440 589700 110492
rect 579436 110236 579488 110288
rect 582012 110236 582064 110288
rect 581828 109692 581880 109744
rect 589464 109692 589516 109744
rect 578332 108332 578384 108384
rect 585140 108332 585192 108384
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 580264 106904 580316 106956
rect 589280 106904 589332 106956
rect 578332 106496 578384 106548
rect 580448 106496 580500 106548
rect 580632 106292 580684 106344
rect 589464 106292 589516 106344
rect 667204 106156 667256 106208
rect 670700 106156 670752 106208
rect 581644 104864 581696 104916
rect 589464 104864 589516 104916
rect 579528 103300 579580 103352
rect 583024 103300 583076 103352
rect 582380 102756 582432 102808
rect 589924 102756 589976 102808
rect 585968 100716 586020 100768
rect 589464 100716 589516 100768
rect 615224 100104 615276 100156
rect 668032 100104 668084 100156
rect 613384 99968 613436 100020
rect 668492 99968 668544 100020
rect 577504 99288 577556 99340
rect 595260 99288 595312 99340
rect 624608 99288 624660 99340
rect 632980 99288 633032 99340
rect 579528 99152 579580 99204
rect 585784 99152 585836 99204
rect 626816 99152 626868 99204
rect 636384 99152 636436 99204
rect 625068 99016 625120 99068
rect 634084 99016 634136 99068
rect 629760 98880 629812 98932
rect 640984 98880 641036 98932
rect 622308 98744 622360 98796
rect 629484 98744 629536 98796
rect 630496 98744 630548 98796
rect 642548 98744 642600 98796
rect 623688 98608 623740 98660
rect 632152 98608 632204 98660
rect 637856 98608 637908 98660
rect 660396 98608 660448 98660
rect 605472 97928 605524 97980
rect 606484 97928 606536 97980
rect 618720 97928 618772 97980
rect 625620 97928 625672 97980
rect 629024 97928 629076 97980
rect 639880 97928 639932 97980
rect 643008 97928 643060 97980
rect 632704 97792 632756 97844
rect 643284 97792 643336 97844
rect 623136 97656 623188 97708
rect 630864 97656 630916 97708
rect 633348 97656 633400 97708
rect 643468 97656 643520 97708
rect 647148 97656 647200 97708
rect 657544 97792 657596 97844
rect 658188 97928 658240 97980
rect 663064 97928 663116 97980
rect 659752 97792 659804 97844
rect 659936 97792 659988 97844
rect 665180 97792 665232 97844
rect 655428 97656 655480 97708
rect 615040 97520 615092 97572
rect 616144 97520 616196 97572
rect 621664 97520 621716 97572
rect 628380 97520 628432 97572
rect 631876 97520 631928 97572
rect 644940 97520 644992 97572
rect 579528 97452 579580 97504
rect 584404 97452 584456 97504
rect 627552 97384 627604 97436
rect 637580 97384 637632 97436
rect 644296 97384 644348 97436
rect 658832 97520 658884 97572
rect 659200 97656 659252 97708
rect 663892 97656 663944 97708
rect 662512 97520 662564 97572
rect 654600 97384 654652 97436
rect 659568 97384 659620 97436
rect 612648 97248 612700 97300
rect 620284 97248 620336 97300
rect 628196 97248 628248 97300
rect 639052 97248 639104 97300
rect 643744 97248 643796 97300
rect 650828 97248 650880 97300
rect 651104 97248 651156 97300
rect 655060 97248 655112 97300
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 620100 97112 620152 97164
rect 626264 97112 626316 97164
rect 634268 97112 634320 97164
rect 644756 97112 644808 97164
rect 650368 97112 650420 97164
rect 658280 97112 658332 97164
rect 634728 96976 634780 97028
rect 643744 96976 643796 97028
rect 651840 96976 651892 97028
rect 654600 96976 654652 97028
rect 597652 96908 597704 96960
rect 598204 96908 598256 96960
rect 615776 96908 615828 96960
rect 618904 96908 618956 96960
rect 645216 96908 645268 96960
rect 649264 96908 649316 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 660672 96908 660724 96960
rect 663432 96908 663484 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 626080 96840 626132 96892
rect 635280 96840 635332 96892
rect 653956 96772 654008 96824
rect 655244 96772 655296 96824
rect 657544 96772 657596 96824
rect 661960 96772 662012 96824
rect 606208 96704 606260 96756
rect 612004 96704 612056 96756
rect 617248 96704 617300 96756
rect 618168 96704 618220 96756
rect 646688 96704 646740 96756
rect 647884 96704 647936 96756
rect 631232 96568 631284 96620
rect 643192 96568 643244 96620
rect 642272 96432 642324 96484
rect 644480 96568 644532 96620
rect 649632 96568 649684 96620
rect 650644 96568 650696 96620
rect 652576 96568 652628 96620
rect 665364 96568 665416 96620
rect 609152 96296 609204 96348
rect 621664 96296 621716 96348
rect 640064 96296 640116 96348
rect 647700 96432 647752 96484
rect 648160 96432 648212 96484
rect 652024 96432 652076 96484
rect 643928 96296 643980 96348
rect 653864 96432 653916 96484
rect 653312 96296 653364 96348
rect 664168 96296 664220 96348
rect 610624 96160 610676 96212
rect 623044 96160 623096 96212
rect 640800 96160 640852 96212
rect 663708 96160 663760 96212
rect 583024 96024 583076 96076
rect 600412 96024 600464 96076
rect 607680 96024 607732 96076
rect 620468 96024 620520 96076
rect 620928 96024 620980 96076
rect 626448 96024 626500 96076
rect 641536 96024 641588 96076
rect 663248 96024 663300 96076
rect 577504 95888 577556 95940
rect 598940 95888 598992 95940
rect 613568 95888 613620 95940
rect 635464 95888 635516 95940
rect 639328 95888 639380 95940
rect 643928 95888 643980 95940
rect 647700 95888 647752 95940
rect 653404 95888 653456 95940
rect 646044 95752 646096 95804
rect 648896 95752 648948 95804
rect 664628 95888 664680 95940
rect 638132 95616 638184 95668
rect 638316 95616 638368 95668
rect 638592 95616 638644 95668
rect 646228 95616 646280 95668
rect 648528 95480 648580 95532
rect 579528 95004 579580 95056
rect 582380 95004 582432 95056
rect 616512 94596 616564 94648
rect 625344 94596 625396 94648
rect 584404 94460 584456 94512
rect 601884 94460 601936 94512
rect 608416 94460 608468 94512
rect 624424 94460 624476 94512
rect 578516 93780 578568 93832
rect 588728 93780 588780 93832
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 644480 93780 644532 93832
rect 654876 93780 654928 93832
rect 580448 93100 580500 93152
rect 590108 93100 590160 93152
rect 664444 92488 664496 92540
rect 668308 92488 668360 92540
rect 617984 92420 618036 92472
rect 625436 92420 625488 92472
rect 648528 92420 648580 92472
rect 655428 92420 655480 92472
rect 611268 90992 611320 91044
rect 617340 90992 617392 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 579068 89700 579120 89752
rect 580632 89700 580684 89752
rect 620468 89632 620520 89684
rect 626448 89632 626500 89684
rect 645768 88748 645820 88800
rect 657452 88748 657504 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 579528 88272 579580 88324
rect 587164 88272 587216 88324
rect 607220 88272 607272 88324
rect 626448 88272 626500 88324
rect 655060 88272 655112 88324
rect 658464 88272 658516 88324
rect 617340 88136 617392 88188
rect 625620 88136 625672 88188
rect 647884 87116 647936 87168
rect 657176 87116 657228 87168
rect 650828 86980 650880 87032
rect 661408 86980 661460 87032
rect 649264 86844 649316 86896
rect 660672 86844 660724 86896
rect 578516 86708 578568 86760
rect 580264 86708 580316 86760
rect 650644 86708 650696 86760
rect 658832 86708 658884 86760
rect 659568 86708 659620 86760
rect 663432 86708 663484 86760
rect 652024 86572 652076 86624
rect 662512 86572 662564 86624
rect 623044 86436 623096 86488
rect 626448 86436 626500 86488
rect 653404 86436 653456 86488
rect 660120 86436 660172 86488
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 621664 84124 621716 84176
rect 625620 84124 625672 84176
rect 579344 83988 579396 84040
rect 581828 83988 581880 84040
rect 579252 82764 579304 82816
rect 588544 82764 588596 82816
rect 628656 80928 628708 80980
rect 642456 80928 642508 80980
rect 614028 80792 614080 80844
rect 647332 80792 647384 80844
rect 595444 80656 595496 80708
rect 636108 80656 636160 80708
rect 579252 80044 579304 80096
rect 585968 80044 586020 80096
rect 629208 79432 629260 79484
rect 638868 79432 638920 79484
rect 616144 79296 616196 79348
rect 648988 79296 649040 79348
rect 638868 78276 638920 78328
rect 645308 78276 645360 78328
rect 631048 78072 631100 78124
rect 639052 78072 639104 78124
rect 612648 77936 612700 77988
rect 647516 77936 647568 77988
rect 628196 77528 628248 77580
rect 633900 77528 633952 77580
rect 578884 77392 578936 77444
rect 631048 77392 631100 77444
rect 589924 77256 589976 77308
rect 628196 77256 628248 77308
rect 628380 77256 628432 77308
rect 631508 77256 631560 77308
rect 620284 76780 620336 76832
rect 649172 76780 649224 76832
rect 612004 76644 612056 76696
rect 647056 76644 647108 76696
rect 606484 76508 606536 76560
rect 662420 76508 662472 76560
rect 579252 75556 579304 75608
rect 581644 75556 581696 75608
rect 618904 75148 618956 75200
rect 646872 75148 646924 75200
rect 588544 74808 588596 74860
rect 628012 74808 628064 74860
rect 578608 73108 578660 73160
rect 580448 73108 580500 73160
rect 579528 67600 579580 67652
rect 624424 67600 624476 67652
rect 579528 66240 579580 66292
rect 605840 66240 605892 66292
rect 581644 65492 581696 65544
rect 603080 65492 603132 65544
rect 579528 64812 579580 64864
rect 613384 64812 613436 64864
rect 580264 62772 580316 62824
rect 601884 62772 601936 62824
rect 578516 62024 578568 62076
rect 664444 62024 664496 62076
rect 579528 60664 579580 60716
rect 614856 60664 614908 60716
rect 579068 58624 579120 58676
rect 600504 58624 600556 58676
rect 605840 58624 605892 58676
rect 663800 58624 663852 58676
rect 579528 57876 579580 57928
rect 666560 57876 666612 57928
rect 579528 56516 579580 56568
rect 588544 56516 588596 56568
rect 574928 56108 574980 56160
rect 596456 56108 596508 56160
rect 574560 55972 574612 56024
rect 596180 55972 596232 56024
rect 574744 55836 574796 55888
rect 599124 55836 599176 55888
rect 624424 55836 624476 55888
rect 663984 55836 664036 55888
rect 459468 53592 459520 53644
rect 577504 55156 577556 55208
rect 465172 53592 465224 53644
rect 465724 53592 465776 53644
rect 465908 53592 465960 53644
rect 585784 55020 585836 55072
rect 583024 54884 583076 54936
rect 589924 54748 589976 54800
rect 597836 54612 597888 54664
rect 597652 54476 597704 54528
rect 578884 54340 578936 54392
rect 469956 53592 470008 53644
rect 470140 53592 470192 53644
rect 470416 53592 470468 53644
rect 461308 53456 461360 53508
rect 579068 54204 579120 54256
rect 477960 53592 478012 53644
rect 574744 54068 574796 54120
rect 574560 53932 574612 53984
rect 481732 53592 481784 53644
rect 482008 53592 482060 53644
rect 574928 53796 574980 53848
rect 50528 53320 50580 53372
rect 129004 53320 129056 53372
rect 463608 53320 463660 53372
rect 470140 53320 470192 53372
rect 47768 53184 47820 53236
rect 130384 53184 130436 53236
rect 463148 53184 463200 53236
rect 477960 53184 478012 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 46204 53048 46256 53100
rect 130568 53048 130620 53100
rect 464896 53048 464948 53100
rect 481732 53048 481784 53100
rect 464068 52912 464120 52964
rect 482008 52912 482060 52964
rect 460066 52776 460118 52828
rect 464206 52776 464258 52828
rect 469956 52776 470008 52828
rect 470416 52640 470468 52692
rect 145380 52436 145432 52488
rect 306012 52436 306064 52488
rect 50712 51960 50764 52012
rect 130752 51960 130804 52012
rect 49148 51824 49200 51876
rect 127164 51824 127216 51876
rect 48964 51688 49016 51740
rect 129464 51688 129516 51740
rect 127164 50736 127216 50788
rect 129280 50736 129332 50788
rect 50344 50464 50396 50516
rect 128636 50464 128688 50516
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 129004 50328 129056 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 51724 49104 51776 49156
rect 128452 49104 128504 49156
rect 47584 48968 47636 49020
rect 129648 48968 129700 49020
rect 128636 47812 128688 47864
rect 132132 47812 132184 47864
rect 129556 45024 129608 45076
rect 129740 44888 129792 44940
rect 128452 44752 128504 44804
rect 129372 44548 129424 44600
rect 129188 44412 129240 44464
rect 132132 44448 132184 44500
rect 132408 44412 132460 44464
rect 130752 44276 130804 44328
rect 129004 44140 129056 44192
rect 132224 44140 132276 44192
rect 130568 44004 130620 44056
rect 130384 43868 130436 43920
rect 43444 42780 43496 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 307300 42712 307352 42764
rect 369400 42712 369452 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 464344 42712 464396 42764
rect 427084 42576 427136 42628
rect 455880 42576 455932 42628
rect 463976 42576 464028 42628
rect 361764 42440 361816 42492
rect 369400 42440 369452 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 308956 42173 309008 42225
rect 427084 42032 427136 42084
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 455880 41896 455932 41948
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 113824 1007412 113876 1007418
rect 113824 1007354 113876 1007360
rect 106832 1007344 106884 1007350
rect 106830 1007312 106832 1007321
rect 106884 1007312 106886 1007321
rect 106830 1007247 106886 1007256
rect 101954 1006632 102010 1006641
rect 94504 1006596 94556 1006602
rect 101954 1006567 101956 1006576
rect 94504 1006538 94556 1006544
rect 102008 1006567 102010 1006576
rect 101956 1006538 102008 1006544
rect 93124 1006324 93176 1006330
rect 93124 1006266 93176 1006272
rect 92296 1003944 92348 1003950
rect 92296 1003886 92348 1003892
rect 92308 998850 92336 1003886
rect 92296 998844 92348 998850
rect 92296 998786 92348 998792
rect 92940 998844 92992 998850
rect 92940 998786 92992 998792
rect 92388 998436 92440 998442
rect 92388 998378 92440 998384
rect 84658 995752 84714 995761
rect 84502 995710 84658 995738
rect 85210 995752 85266 995761
rect 85054 995710 85210 995738
rect 84658 995687 84714 995696
rect 86038 995752 86094 995761
rect 85698 995710 86038 995738
rect 85210 995687 85266 995696
rect 90270 995752 90326 995761
rect 90022 995710 90270 995738
rect 86038 995687 86094 995696
rect 90270 995687 90326 995696
rect 88982 995616 89038 995625
rect 88734 995574 88982 995602
rect 89534 995616 89590 995625
rect 89378 995574 89534 995602
rect 88982 995551 89038 995560
rect 89534 995551 89590 995560
rect 77050 995438 77248 995466
rect 77220 995353 77248 995438
rect 77206 995344 77262 995353
rect 77206 995279 77262 995288
rect 77680 994566 77708 995452
rect 78324 994838 78352 995452
rect 80164 995081 80192 995452
rect 80730 995438 81112 995466
rect 80150 995072 80206 995081
rect 80150 995007 80206 995016
rect 78312 994832 78364 994838
rect 78312 994774 78364 994780
rect 77668 994560 77720 994566
rect 77668 994502 77720 994508
rect 81084 993993 81112 995438
rect 81360 994702 81388 995452
rect 82004 994809 82032 995452
rect 81990 994800 82046 994809
rect 81990 994735 82046 994744
rect 81348 994696 81400 994702
rect 81348 994638 81400 994644
rect 86328 994537 86356 995452
rect 87538 995438 87920 995466
rect 91218 995438 91692 995466
rect 86314 994528 86370 994537
rect 86314 994463 86370 994472
rect 87892 994265 87920 995438
rect 91664 995330 91692 995438
rect 92400 995330 92428 998378
rect 92756 998028 92808 998034
rect 92756 997970 92808 997976
rect 92572 997688 92624 997694
rect 92572 997630 92624 997636
rect 92584 997257 92612 997630
rect 92570 997248 92626 997257
rect 92570 997183 92626 997192
rect 92768 996305 92796 997970
rect 92952 996985 92980 998786
rect 92938 996976 92994 996985
rect 92938 996911 92994 996920
rect 92754 996296 92810 996305
rect 92754 996231 92810 996240
rect 91664 995302 92428 995330
rect 93136 994809 93164 1006266
rect 93308 1006188 93360 1006194
rect 93308 1006130 93360 1006136
rect 93122 994800 93178 994809
rect 93122 994735 93178 994744
rect 93320 994566 93348 1006130
rect 93492 997892 93544 997898
rect 93492 997834 93544 997840
rect 93504 995761 93532 997834
rect 93490 995752 93546 995761
rect 93490 995687 93546 995696
rect 93308 994560 93360 994566
rect 93308 994502 93360 994508
rect 87878 994256 87934 994265
rect 87878 994191 87934 994200
rect 94516 993993 94544 1006538
rect 104806 1006496 104862 1006505
rect 101588 1006460 101640 1006466
rect 104806 1006431 104808 1006440
rect 101588 1006402 101640 1006408
rect 104860 1006431 104862 1006440
rect 104808 1006402 104860 1006408
rect 100298 1006360 100354 1006369
rect 100298 1006295 100300 1006304
rect 100352 1006295 100354 1006304
rect 100300 1006266 100352 1006272
rect 101404 1006188 101456 1006194
rect 101404 1006130 101456 1006136
rect 98274 1006088 98330 1006097
rect 94688 1006052 94740 1006058
rect 98274 1006023 98276 1006032
rect 94688 1005994 94740 1006000
rect 98328 1006023 98330 1006032
rect 98276 1005994 98328 1006000
rect 94700 997898 94728 1005994
rect 98644 1002652 98696 1002658
rect 98644 1002594 98696 1002600
rect 97448 1002516 97500 1002522
rect 97448 1002458 97500 1002464
rect 96068 1002380 96120 1002386
rect 96068 1002322 96120 1002328
rect 95884 1001972 95936 1001978
rect 95884 1001914 95936 1001920
rect 95148 999184 95200 999190
rect 95148 999126 95200 999132
rect 94688 997892 94740 997898
rect 94688 997834 94740 997840
rect 95160 994265 95188 999126
rect 95146 994256 95202 994265
rect 95146 994191 95202 994200
rect 81070 993984 81126 993993
rect 81070 993919 81126 993928
rect 94502 993984 94558 993993
rect 94502 993919 94558 993928
rect 50344 993200 50396 993206
rect 50344 993142 50396 993148
rect 44824 993064 44876 993070
rect 44824 993006 44876 993012
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 969218 42196 969272
rect 42260 969258 42564 969286
rect 42260 969218 42288 969258
rect 42168 969190 42288 969218
rect 42536 968810 42564 969258
rect 42536 968782 42840 968810
rect 42168 967609 42196 968048
rect 42154 967600 42210 967609
rect 42154 967535 42210 967544
rect 42614 967600 42670 967609
rect 42614 967535 42670 967544
rect 41800 967201 41828 967405
rect 41786 967192 41842 967201
rect 41786 967127 41842 967136
rect 42154 967192 42210 967201
rect 42154 967127 42210 967136
rect 42168 966756 42196 967127
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42444 963937 42472 964362
rect 42430 963928 42486 963937
rect 42430 963863 42486 963872
rect 42182 963711 42472 963739
rect 42444 963393 42472 963711
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42430 963112 42486 963121
rect 42182 963070 42430 963098
rect 42430 963047 42486 963056
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 41786 959103 41842 959112
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 41800 957817 41828 958188
rect 41786 957808 41842 957817
rect 41786 957743 41842 957752
rect 42182 956338 42288 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 41800 954689 41828 955060
rect 41786 954680 41842 954689
rect 41786 954615 41842 954624
rect 41786 954408 41842 954417
rect 41786 954343 41842 954352
rect 35162 952912 35218 952921
rect 35162 952847 35218 952856
rect 33784 951516 33836 951522
rect 33784 951458 33836 951464
rect 31758 946656 31814 946665
rect 31758 946591 31814 946600
rect 31772 945334 31800 946591
rect 28724 945328 28776 945334
rect 28724 945270 28776 945276
rect 31760 945328 31812 945334
rect 31760 945270 31812 945276
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28736 942721 28764 945270
rect 28722 942712 28778 942721
rect 28722 942647 28778 942656
rect 33796 938233 33824 951458
rect 33782 938224 33838 938233
rect 33782 938159 33838 938168
rect 35176 937825 35204 952847
rect 41800 952626 41828 954343
rect 41524 952598 41828 952626
rect 37922 952504 37978 952513
rect 37922 952439 37978 952448
rect 36544 952400 36596 952406
rect 36544 952342 36596 952348
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35820 942614 35848 943055
rect 35808 942608 35860 942614
rect 35808 942550 35860 942556
rect 35806 941896 35862 941905
rect 35806 941831 35862 941840
rect 35820 941254 35848 941831
rect 35808 941248 35860 941254
rect 35808 941190 35860 941196
rect 35806 940264 35862 940273
rect 35806 940199 35862 940208
rect 35820 939826 35848 940199
rect 35808 939820 35860 939826
rect 35808 939762 35860 939768
rect 36556 939049 36584 952342
rect 36542 939040 36598 939049
rect 36542 938975 36598 938984
rect 37936 938641 37964 952439
rect 39302 952232 39358 952241
rect 39302 952167 39358 952176
rect 37922 938632 37978 938641
rect 37922 938567 37978 938576
rect 35162 937816 35218 937825
rect 35162 937751 35218 937760
rect 39316 937417 39344 952167
rect 40038 951688 40094 951697
rect 40038 951623 40094 951632
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 40052 934561 40080 951623
rect 41524 951522 41552 952598
rect 42260 952490 42288 956338
rect 41708 952462 42288 952490
rect 41708 952406 41736 952462
rect 41696 952400 41748 952406
rect 41696 952342 41748 952348
rect 41512 951516 41564 951522
rect 41512 951458 41564 951464
rect 42628 949454 42656 967535
rect 42536 949426 42656 949454
rect 41696 942608 41748 942614
rect 41748 942556 41920 942562
rect 41696 942550 41920 942556
rect 41708 942534 41920 942550
rect 41696 941180 41748 941186
rect 41696 941122 41748 941128
rect 41512 939820 41564 939826
rect 41512 939762 41564 939768
rect 40038 934552 40094 934561
rect 40038 934487 40094 934496
rect 41524 911713 41552 939762
rect 41708 911985 41736 941122
rect 41892 937034 41920 942534
rect 42062 940672 42118 940681
rect 42062 940607 42118 940616
rect 42076 939865 42104 940607
rect 42062 939856 42118 939865
rect 42062 939791 42118 939800
rect 42536 939794 42564 949426
rect 42260 939766 42564 939794
rect 41892 937006 42104 937034
rect 42076 935785 42104 937006
rect 42062 935776 42118 935785
rect 42062 935711 42118 935720
rect 42260 932929 42288 939766
rect 42812 937009 42840 968782
rect 43456 967201 43484 975666
rect 43442 967192 43498 967201
rect 43442 967127 43498 967136
rect 43442 964744 43498 964753
rect 43442 964679 43498 964688
rect 43258 963928 43314 963937
rect 43258 963863 43314 963872
rect 43074 963384 43130 963393
rect 43074 963319 43130 963328
rect 42798 937000 42854 937009
rect 42798 936935 42854 936944
rect 43088 934969 43116 963319
rect 43074 934960 43130 934969
rect 43074 934895 43130 934904
rect 43272 933745 43300 963863
rect 43456 935377 43484 964679
rect 44270 963112 44326 963121
rect 44270 963047 44326 963056
rect 43442 935368 43498 935377
rect 43442 935303 43498 935312
rect 44284 934153 44312 963047
rect 44454 958760 44510 958769
rect 44454 958695 44510 958704
rect 44468 936193 44496 958695
rect 44836 941497 44864 993006
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 46204 961920 46256 961926
rect 46204 961862 46256 961868
rect 46216 946665 46244 961862
rect 46202 946656 46258 946665
rect 46202 946591 46258 946600
rect 45560 946008 45612 946014
rect 45560 945950 45612 945956
rect 45572 943537 45600 945950
rect 45558 943528 45614 943537
rect 45558 943463 45614 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44638 941080 44694 941089
rect 44638 941015 44694 941024
rect 44454 936184 44510 936193
rect 44454 936119 44510 936128
rect 44270 934144 44326 934153
rect 44270 934079 44326 934088
rect 43258 933736 43314 933745
rect 43258 933671 43314 933680
rect 43350 933328 43406 933337
rect 43350 933263 43406 933272
rect 42246 932920 42302 932929
rect 42246 932855 42302 932864
rect 41694 911976 41750 911985
rect 41694 911911 41750 911920
rect 41510 911704 41566 911713
rect 41510 911639 41566 911648
rect 42936 892528 42992 892537
rect 42936 892463 42992 892472
rect 42950 892328 42978 892463
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43074 892256 43130 892265
rect 43074 892191 43130 892200
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817086 35848 817255
rect 35808 817080 35860 817086
rect 35808 817022 35860 817028
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 815658 35848 816439
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814298 35848 814807
rect 41432 814298 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815674 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815658 41644 815674
rect 41524 815652 41656 815658
rect 41524 815646 41604 815652
rect 41604 815594 41656 815600
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41420 814292 41472 814298
rect 41420 814234 41472 814240
rect 41326 812832 41382 812841
rect 41326 812767 41382 812776
rect 40958 812424 41014 812433
rect 40958 812359 41014 812368
rect 35162 811608 35218 811617
rect 35162 811543 35218 811552
rect 35176 802466 35204 811543
rect 35898 811200 35954 811209
rect 35898 811135 35954 811144
rect 35164 802460 35216 802466
rect 35164 802402 35216 802408
rect 35912 802330 35940 811135
rect 40776 808988 40828 808994
rect 40776 808930 40828 808936
rect 40590 808344 40646 808353
rect 40590 808279 40646 808288
rect 40604 805089 40632 808279
rect 40788 805497 40816 808930
rect 40774 805488 40830 805497
rect 40774 805423 40830 805432
rect 40972 805361 41000 812359
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 41156 805633 41184 811951
rect 41340 811646 41368 812767
rect 41328 811640 41380 811646
rect 41328 811582 41380 811588
rect 41696 811640 41748 811646
rect 41696 811582 41748 811588
rect 41708 811458 41736 811582
rect 41708 811430 42472 811458
rect 41786 809160 41842 809169
rect 41616 809118 41786 809146
rect 41616 808994 41644 809118
rect 41786 809095 41842 809104
rect 41604 808988 41656 808994
rect 41604 808930 41656 808936
rect 42246 806712 42302 806721
rect 42246 806647 42302 806656
rect 41142 805624 41198 805633
rect 41142 805559 41198 805568
rect 40958 805352 41014 805361
rect 40958 805287 41014 805296
rect 40590 805080 40646 805089
rect 40590 805015 40646 805024
rect 41694 802496 41750 802505
rect 41694 802431 41696 802440
rect 41748 802431 41750 802440
rect 41696 802402 41748 802408
rect 35900 802324 35952 802330
rect 35900 802266 35952 802272
rect 41696 802324 41748 802330
rect 41696 802266 41748 802272
rect 41708 802210 41736 802266
rect 41708 802182 41828 802210
rect 41800 800329 41828 802182
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 806647
rect 42444 804554 42472 811430
rect 43166 810792 43222 810801
rect 43166 810727 43222 810736
rect 42798 809976 42854 809985
rect 42798 809911 42854 809920
rect 42182 798238 42288 798266
rect 42352 804526 42472 804554
rect 42352 797619 42380 804526
rect 42522 802496 42578 802505
rect 42578 802454 42748 802482
rect 42522 802431 42578 802440
rect 42522 798960 42578 798969
rect 42522 798895 42578 798904
rect 42182 797591 42380 797619
rect 42536 796974 42564 798895
rect 42182 796946 42564 796974
rect 42154 796240 42210 796249
rect 42154 796175 42210 796184
rect 42168 795765 42196 796175
rect 42522 795424 42578 795433
rect 42522 795359 42578 795368
rect 42536 795274 42564 795359
rect 42444 795246 42564 795274
rect 42062 795016 42118 795025
rect 42062 794951 42118 794960
rect 42076 794580 42104 794951
rect 41786 794200 41842 794209
rect 41786 794135 41842 794144
rect 41800 793900 41828 794135
rect 42444 793302 42472 795246
rect 42720 794894 42748 802454
rect 42182 793274 42472 793302
rect 42536 794866 42748 794894
rect 42536 792758 42564 794866
rect 42182 792730 42564 792758
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42812 792146 42840 809911
rect 42982 807528 43038 807537
rect 42982 807463 43038 807472
rect 42720 792134 42840 792146
rect 42168 790622 42288 790650
rect 42352 792118 42840 792134
rect 42352 792106 42748 792118
rect 42168 790228 42196 790622
rect 42352 789630 42380 792106
rect 42182 789602 42380 789630
rect 42154 789304 42210 789313
rect 42154 789239 42210 789248
rect 42168 788936 42196 789239
rect 42706 789032 42762 789041
rect 42536 788990 42706 789018
rect 41786 788624 41842 788633
rect 41786 788559 41842 788568
rect 41800 788392 41828 788559
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 41786 786856 41842 786865
rect 41786 786791 41842 786800
rect 41800 786556 41828 786791
rect 42260 786162 42288 788151
rect 42076 786134 42288 786162
rect 42076 785944 42104 786134
rect 42536 785278 42564 788990
rect 42706 788967 42762 788976
rect 42706 788624 42762 788633
rect 42706 788559 42762 788568
rect 42182 785250 42564 785278
rect 42720 779714 42748 788559
rect 41708 779686 42748 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 772886 35848 773463
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 35622 769448 35678 769457
rect 35622 769383 35678 769392
rect 35438 769040 35494 769049
rect 35438 768975 35494 768984
rect 35452 768738 35480 768975
rect 35636 768874 35664 769383
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35860 768975 35862 768984
rect 41328 769004 41380 769010
rect 35808 768946 35860 768952
rect 41328 768946 41380 768952
rect 35624 768868 35676 768874
rect 35624 768810 35676 768816
rect 35440 768732 35492 768738
rect 35440 768674 35492 768680
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 31022 768224 31078 768233
rect 31022 768159 31078 768168
rect 31036 758266 31064 768159
rect 35530 767816 35586 767825
rect 35530 767751 35586 767760
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35544 767378 35572 767751
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35532 767372 35584 767378
rect 35532 767314 35584 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 35176 758470 35204 766935
rect 35164 758464 35216 758470
rect 35164 758406 35216 758412
rect 31024 758260 31076 758266
rect 31024 758202 31076 758208
rect 36556 757761 36584 767450
rect 37924 767372 37976 767378
rect 37924 767314 37976 767320
rect 37094 763328 37150 763337
rect 37094 763263 37096 763272
rect 37148 763263 37150 763272
rect 37096 763234 37148 763240
rect 37936 759082 37964 767314
rect 40052 764561 40080 768674
rect 41340 765785 41368 768946
rect 41696 768868 41748 768874
rect 41696 768810 41748 768816
rect 41708 765914 41736 768810
rect 41524 765886 41736 765914
rect 41326 765776 41382 765785
rect 41326 765711 41382 765720
rect 40038 764552 40094 764561
rect 40038 764487 40094 764496
rect 39304 763292 39356 763298
rect 39304 763234 39356 763240
rect 37924 759076 37976 759082
rect 37924 759018 37976 759024
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 39316 757654 39344 763234
rect 39488 759076 39540 759082
rect 39488 759018 39540 759024
rect 39304 757648 39356 757654
rect 39304 757590 39356 757596
rect 39500 757353 39528 759018
rect 40684 758192 40736 758198
rect 40682 758160 40684 758169
rect 40736 758160 40738 758169
rect 40682 758095 40738 758104
rect 41524 757874 41552 765886
rect 42706 765776 42762 765785
rect 42706 765711 42762 765720
rect 42720 763154 42748 765711
rect 42628 763126 42748 763154
rect 41696 758464 41748 758470
rect 41748 758412 42104 758418
rect 41696 758406 42104 758412
rect 41708 758402 42104 758406
rect 41708 758396 42116 758402
rect 41708 758390 42064 758396
rect 42064 758338 42116 758344
rect 42064 758056 42116 758062
rect 42116 758004 42564 758010
rect 42064 757998 42564 758004
rect 42076 757982 42564 757998
rect 41524 757846 42472 757874
rect 41696 757648 41748 757654
rect 41748 757596 42288 757602
rect 41696 757590 42288 757596
rect 41708 757574 42288 757590
rect 39486 757344 39542 757353
rect 39486 757279 39542 757288
rect 41786 756664 41842 756673
rect 42260 756650 42288 757574
rect 42260 756622 42380 756650
rect 41786 756599 41842 756608
rect 41800 756228 41828 756599
rect 42168 755018 42196 755072
rect 42352 755018 42380 756622
rect 42168 754990 42380 755018
rect 42444 754610 42472 757846
rect 42168 754582 42472 754610
rect 42168 754392 42196 754582
rect 42338 754216 42394 754225
rect 42338 754151 42394 754160
rect 41970 754080 42026 754089
rect 41970 754015 42026 754024
rect 41984 753780 42012 754015
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42154 751768 42210 751777
rect 42154 751703 42210 751712
rect 42168 751369 42196 751703
rect 42352 750734 42380 754151
rect 42536 753494 42564 757982
rect 42182 750706 42380 750734
rect 42444 753466 42564 753494
rect 42246 750544 42302 750553
rect 42246 750479 42302 750488
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42260 749543 42288 750479
rect 42182 749515 42288 749543
rect 41786 747416 41842 747425
rect 41786 747351 41842 747360
rect 41800 747048 41828 747351
rect 42154 746736 42210 746745
rect 42154 746671 42210 746680
rect 42168 746401 42196 746671
rect 42444 745770 42472 753466
rect 42628 750258 42656 763126
rect 42798 757888 42854 757897
rect 42798 757823 42854 757832
rect 42812 750553 42840 757823
rect 42798 750544 42854 750553
rect 42798 750479 42854 750488
rect 42628 750230 42748 750258
rect 42182 745742 42472 745770
rect 42720 745362 42748 750230
rect 42536 745334 42748 745362
rect 42536 745226 42564 745334
rect 42182 745198 42564 745226
rect 42430 745104 42486 745113
rect 42430 745039 42486 745048
rect 42246 744832 42302 744841
rect 42246 744767 42302 744776
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743050 42288 744767
rect 42168 743022 42288 743050
rect 42168 742696 42196 743022
rect 42444 742098 42472 745039
rect 42614 743064 42670 743073
rect 42614 742999 42670 743008
rect 42182 742070 42472 742098
rect 42628 741962 42656 742999
rect 42260 741934 42656 741962
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42260 731414 42288 741934
rect 42430 741704 42486 741713
rect 42430 741639 42486 741648
rect 42444 731414 42472 741639
rect 41708 731386 42288 731414
rect 42352 731386 42472 731414
rect 35622 731368 35678 731377
rect 35622 731303 35678 731312
rect 35636 730114 35664 731303
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35820 730250 35848 730895
rect 41708 730250 41736 731386
rect 35808 730244 35860 730250
rect 35808 730186 35860 730192
rect 41696 730244 41748 730250
rect 41696 730186 41748 730192
rect 42352 730130 42380 731386
rect 41708 730114 42380 730130
rect 35624 730108 35676 730114
rect 35624 730050 35676 730056
rect 41696 730108 42380 730114
rect 41748 730102 42380 730108
rect 41696 730050 41748 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41142 726064 41198 726073
rect 41142 725999 41198 726008
rect 31022 725248 31078 725257
rect 31022 725183 31078 725192
rect 31036 716854 31064 725183
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 33046 724024 33102 724033
rect 33046 723959 33102 723968
rect 31024 716848 31076 716854
rect 31024 716790 31076 716796
rect 33060 715562 33088 723959
rect 33782 723208 33838 723217
rect 33782 723143 33838 723152
rect 33796 715698 33824 723143
rect 33784 715692 33836 715698
rect 33784 715634 33836 715640
rect 33048 715556 33100 715562
rect 33048 715498 33100 715504
rect 36556 715426 36584 724775
rect 40682 724432 40738 724441
rect 40682 724367 40738 724376
rect 36544 715420 36596 715426
rect 36544 715362 36596 715368
rect 40696 714785 40724 724367
rect 41156 721777 41184 725999
rect 41340 725966 41368 726407
rect 41328 725960 41380 725966
rect 41328 725902 41380 725908
rect 41696 725960 41748 725966
rect 41748 725908 41920 725914
rect 41696 725902 41920 725908
rect 41708 725886 41920 725902
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724538 41368 725591
rect 41328 724532 41380 724538
rect 41328 724474 41380 724480
rect 41696 724532 41748 724538
rect 41696 724474 41748 724480
rect 41142 721768 41198 721777
rect 41708 721754 41736 724474
rect 41892 721754 41920 725886
rect 41708 721726 41828 721754
rect 41892 721726 42472 721754
rect 41142 721703 41198 721712
rect 41326 720352 41382 720361
rect 41326 720287 41382 720296
rect 40682 714776 40738 714785
rect 40682 714711 40738 714720
rect 41340 714241 41368 720287
rect 41800 717614 41828 721726
rect 42444 717614 42472 721726
rect 41800 717586 41920 717614
rect 41604 716848 41656 716854
rect 41604 716790 41656 716796
rect 41616 715873 41644 716790
rect 41602 715864 41658 715873
rect 41602 715799 41658 715808
rect 41512 715692 41564 715698
rect 41512 715634 41564 715640
rect 41524 715170 41552 715634
rect 41892 715601 41920 717586
rect 42352 717586 42472 717614
rect 41878 715592 41934 715601
rect 41696 715556 41748 715562
rect 41878 715527 41934 715536
rect 41696 715498 41748 715504
rect 41708 715306 41736 715498
rect 42352 715442 42380 717586
rect 42706 715864 42762 715873
rect 42762 715822 42932 715850
rect 42706 715799 42762 715808
rect 42614 715592 42670 715601
rect 42614 715527 42670 715536
rect 42352 715414 42564 715442
rect 41708 715278 42472 715306
rect 41524 715142 42380 715170
rect 41604 715080 41656 715086
rect 41656 715028 41828 715034
rect 41604 715022 41828 715028
rect 41616 715006 41828 715022
rect 41326 714232 41382 714241
rect 41326 714167 41382 714176
rect 41800 713969 41828 715006
rect 42352 714762 42380 715142
rect 42076 714734 42380 714762
rect 42076 714513 42104 714734
rect 42062 714504 42118 714513
rect 42062 714439 42118 714448
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 41786 713552 41842 713561
rect 41786 713487 41842 713496
rect 41800 713048 41828 713487
rect 42062 713280 42118 713289
rect 42444 713266 42472 715278
rect 42118 713238 42472 713266
rect 42062 713215 42118 713224
rect 42536 712586 42564 715414
rect 42352 712558 42564 712586
rect 41786 712192 41842 712201
rect 41786 712127 41842 712136
rect 41800 711824 41828 712127
rect 42352 711362 42380 712558
rect 42260 711334 42380 711362
rect 42260 711226 42288 711334
rect 42628 711226 42656 715527
rect 42182 711198 42288 711226
rect 42536 711198 42656 711226
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 42536 710002 42564 711198
rect 42706 711104 42762 711113
rect 42706 711039 42762 711048
rect 42352 709974 42564 710002
rect 41878 709880 41934 709889
rect 41878 709815 41934 709824
rect 41892 709376 41920 709815
rect 42154 708520 42210 708529
rect 42154 708455 42210 708464
rect 42168 708152 42196 708455
rect 42062 707704 42118 707713
rect 42062 707639 42118 707648
rect 42076 707540 42104 707639
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42062 706752 42118 706761
rect 42062 706687 42118 706696
rect 42076 706316 42104 706687
rect 42352 706602 42380 709974
rect 42720 708665 42748 711039
rect 42706 708656 42762 708665
rect 42706 708591 42762 708600
rect 42904 707554 42932 715822
rect 42536 707526 42932 707554
rect 42536 706761 42564 707526
rect 42706 707432 42762 707441
rect 42706 707367 42762 707376
rect 42522 706752 42578 706761
rect 42522 706687 42578 706696
rect 42352 706574 42472 706602
rect 42246 706480 42302 706489
rect 42246 706415 42302 706424
rect 42260 704290 42288 706415
rect 42076 704262 42288 704290
rect 42076 703868 42104 704262
rect 42062 703488 42118 703497
rect 42062 703423 42118 703432
rect 42076 703188 42104 703423
rect 42062 702808 42118 702817
rect 42062 702743 42118 702752
rect 42076 702576 42104 702743
rect 42444 702046 42472 706574
rect 42720 702817 42748 707367
rect 42706 702808 42762 702817
rect 42706 702743 42762 702752
rect 42614 702400 42670 702409
rect 42614 702335 42670 702344
rect 42168 701978 42196 702032
rect 42260 702018 42472 702046
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42154 699952 42210 699961
rect 42154 699887 42210 699896
rect 42168 699516 42196 699887
rect 42628 698918 42656 702335
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 41694 697912 41750 697921
rect 41694 697847 41750 697856
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35622 687304 35678 687313
rect 35820 687274 35848 687647
rect 41708 687274 41736 697847
rect 35622 687239 35678 687248
rect 35808 687268 35860 687274
rect 35808 687210 35860 687216
rect 41696 687268 41748 687274
rect 41696 687210 41748 687216
rect 35806 683224 35862 683233
rect 35806 683159 35808 683168
rect 35860 683159 35862 683168
rect 41512 683188 41564 683194
rect 35808 683130 35860 683136
rect 41512 683130 41564 683136
rect 35438 682816 35494 682825
rect 35438 682751 35494 682760
rect 35452 681086 35480 682751
rect 35622 682408 35678 682417
rect 35622 682343 35678 682352
rect 35636 681902 35664 682343
rect 35806 682000 35862 682009
rect 35806 681935 35862 681944
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35820 681766 35848 681935
rect 35808 681760 35860 681766
rect 35808 681702 35860 681708
rect 41328 681760 41380 681766
rect 41524 681748 41552 683130
rect 41696 681896 41748 681902
rect 41748 681844 42196 681850
rect 41696 681838 42196 681844
rect 41708 681822 42196 681838
rect 41524 681720 42104 681748
rect 41328 681702 41380 681708
rect 35622 681592 35678 681601
rect 35622 681527 35678 681536
rect 35440 681080 35492 681086
rect 35440 681022 35492 681028
rect 35162 680776 35218 680785
rect 35162 680711 35218 680720
rect 35176 672790 35204 680711
rect 35636 680406 35664 681527
rect 35806 681184 35862 681193
rect 35806 681119 35862 681128
rect 35820 680678 35848 681119
rect 35808 680672 35860 680678
rect 35808 680614 35860 680620
rect 37924 680672 37976 680678
rect 37924 680614 37976 680620
rect 35624 680400 35676 680406
rect 35624 680342 35676 680348
rect 36544 680400 36596 680406
rect 36544 680342 36596 680348
rect 35164 672784 35216 672790
rect 35164 672726 35216 672732
rect 36556 672110 36584 680342
rect 36544 672104 36596 672110
rect 36544 672046 36596 672052
rect 37936 671265 37964 680614
rect 41340 678858 41368 681702
rect 41604 681080 41656 681086
rect 41786 681048 41842 681057
rect 41656 681028 41786 681034
rect 41604 681022 41786 681028
rect 41616 681006 41786 681022
rect 41786 680983 41842 680992
rect 41340 678830 41552 678858
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 39960 671498 39988 677039
rect 40500 672784 40552 672790
rect 40500 672726 40552 672732
rect 40512 672625 40540 672726
rect 40498 672616 40554 672625
rect 40498 672551 40554 672560
rect 41524 672353 41552 678830
rect 42076 673169 42104 681720
rect 42168 678974 42196 681822
rect 42798 679960 42854 679969
rect 42798 679895 42854 679904
rect 42168 678946 42472 678974
rect 42062 673160 42118 673169
rect 42062 673095 42118 673104
rect 42444 672466 42472 678946
rect 42812 672897 42840 679895
rect 42798 672888 42854 672897
rect 42798 672823 42854 672832
rect 42798 672616 42854 672625
rect 42798 672551 42854 672560
rect 42444 672438 42564 672466
rect 41510 672344 41566 672353
rect 41510 672279 41566 672288
rect 42246 672344 42302 672353
rect 42302 672302 42472 672330
rect 42246 672279 42302 672288
rect 41604 672104 41656 672110
rect 41524 672052 41604 672058
rect 41524 672046 41656 672052
rect 41524 672030 41644 672046
rect 39948 671492 40000 671498
rect 39948 671434 40000 671440
rect 41524 671378 41552 672030
rect 41708 671498 42380 671514
rect 41696 671492 42380 671498
rect 41748 671486 42380 671492
rect 41696 671434 41748 671440
rect 41524 671350 41920 671378
rect 37922 671256 37978 671265
rect 37922 671191 37978 671200
rect 41892 671106 41920 671350
rect 41892 671078 42288 671106
rect 42168 669746 42196 669868
rect 42260 669746 42288 671078
rect 42168 669718 42288 669746
rect 42352 669610 42380 671486
rect 42260 669582 42380 669610
rect 42260 668658 42288 669582
rect 42182 668630 42288 668658
rect 42062 668536 42118 668545
rect 42062 668471 42118 668480
rect 42076 668032 42104 668471
rect 42246 668264 42302 668273
rect 42246 668199 42302 668208
rect 42260 668046 42288 668199
rect 42260 668018 42380 668046
rect 41970 667720 42026 667729
rect 41970 667655 42026 667664
rect 41984 667352 42012 667655
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42352 666554 42380 668018
rect 42260 666526 42380 666554
rect 42260 664986 42288 666526
rect 42182 664958 42288 664986
rect 42246 664864 42302 664873
rect 42246 664799 42302 664808
rect 42260 664714 42288 664799
rect 42168 664686 42288 664714
rect 42168 664325 42196 664686
rect 41786 664048 41842 664057
rect 41786 663983 41842 663992
rect 41800 663680 41828 663983
rect 42444 663898 42472 672302
rect 42536 666554 42564 672438
rect 42536 666526 42656 666554
rect 42260 663870 42472 663898
rect 42260 663150 42288 663870
rect 42430 663504 42486 663513
rect 42430 663439 42486 663448
rect 42182 663122 42288 663150
rect 42246 662688 42302 662697
rect 42246 662623 42302 662632
rect 42260 660770 42288 662623
rect 42168 660742 42288 660770
rect 42168 660620 42196 660742
rect 42444 660362 42472 663439
rect 42168 660334 42472 660362
rect 42168 660008 42196 660334
rect 42628 660022 42656 666526
rect 42444 659994 42656 660022
rect 42076 659161 42104 659357
rect 42062 659152 42118 659161
rect 42062 659087 42118 659096
rect 42168 658838 42288 658866
rect 42168 658784 42196 658838
rect 42260 658798 42288 658838
rect 42444 658798 42472 659994
rect 42614 659696 42670 659705
rect 42614 659631 42670 659640
rect 42260 658770 42472 658798
rect 42430 658608 42486 658617
rect 42430 658543 42486 658552
rect 42246 658336 42302 658345
rect 42246 658271 42302 658280
rect 42062 657384 42118 657393
rect 42062 657319 42118 657328
rect 42076 656948 42104 657319
rect 42260 656350 42288 658271
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42444 655670 42472 658543
rect 42628 657393 42656 659631
rect 42812 659161 42840 672551
rect 42798 659152 42854 659161
rect 42798 659087 42854 659096
rect 42614 657384 42670 657393
rect 42614 657319 42670 657328
rect 42260 655642 42472 655670
rect 35806 646776 35862 646785
rect 35806 646711 35862 646720
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35820 644745 35848 646711
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35806 639840 35862 639849
rect 35806 639775 35862 639784
rect 35820 639198 35848 639775
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 41696 639124 41748 639130
rect 41696 639066 41748 639072
rect 35806 639024 35862 639033
rect 41708 639010 41736 639066
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 40040 638988 40092 638994
rect 35808 638930 35860 638936
rect 41708 638982 42472 639010
rect 40040 638930 40092 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 35820 637634 35848 638551
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 40052 637401 40080 638930
rect 41786 638208 41842 638217
rect 41786 638143 41842 638152
rect 41328 637628 41380 637634
rect 41800 637605 41828 638143
rect 41328 637570 41380 637576
rect 41786 637596 41842 637605
rect 40038 637392 40094 637401
rect 40038 637327 40094 637336
rect 41340 634814 41368 637570
rect 41786 637531 41842 637540
rect 42444 634814 42472 638982
rect 41340 634786 41460 634814
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41432 627745 41460 634786
rect 42352 634786 42472 634814
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 41418 627736 41474 627745
rect 41418 627671 41474 627680
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42062 625832 42118 625841
rect 42062 625767 42118 625776
rect 42076 625464 42104 625767
rect 42352 625682 42380 634786
rect 42522 633856 42578 633865
rect 42522 633791 42578 633800
rect 42536 625841 42564 633791
rect 42706 627736 42762 627745
rect 42706 627671 42762 627680
rect 42522 625832 42578 625841
rect 42522 625767 42578 625776
rect 42352 625654 42564 625682
rect 42536 625410 42564 625654
rect 42352 625382 42564 625410
rect 42352 625002 42380 625382
rect 42168 624974 42380 625002
rect 42522 625016 42578 625025
rect 42168 624784 42196 624974
rect 42522 624951 42578 624960
rect 42536 624186 42564 624951
rect 42182 624158 42564 624186
rect 42246 624064 42302 624073
rect 42246 623999 42302 624008
rect 41970 623384 42026 623393
rect 41970 623319 42026 623328
rect 41984 622948 42012 623319
rect 41786 622160 41842 622169
rect 41786 622095 41842 622104
rect 41800 621792 41828 622095
rect 42260 621602 42288 623999
rect 42430 623384 42486 623393
rect 42430 623319 42486 623328
rect 42168 621574 42288 621602
rect 42168 621112 42196 621574
rect 42444 621330 42472 623319
rect 42260 621302 42472 621330
rect 42168 620378 42196 620500
rect 42260 620378 42288 621302
rect 42720 621058 42748 627671
rect 42168 620350 42288 620378
rect 42352 621030 42748 621058
rect 42352 619970 42380 621030
rect 42522 620120 42578 620129
rect 42522 620055 42578 620064
rect 42168 619834 42196 619956
rect 42260 619942 42380 619970
rect 42260 619834 42288 619942
rect 42168 619806 42288 619834
rect 42536 619290 42564 620055
rect 42706 619848 42762 619857
rect 42706 619783 42762 619792
rect 42352 619262 42564 619290
rect 42352 619018 42380 619262
rect 42260 618990 42380 619018
rect 42260 617454 42288 618990
rect 42430 618896 42486 618905
rect 42430 618831 42486 618840
rect 42444 618610 42472 618831
rect 42444 618582 42656 618610
rect 42430 618488 42486 618497
rect 42430 618423 42486 618432
rect 42182 617426 42288 617454
rect 42444 616842 42472 618423
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42628 616434 42656 618582
rect 42168 616406 42656 616434
rect 42168 616148 42196 616406
rect 42062 615904 42118 615913
rect 42062 615839 42118 615848
rect 42076 615604 42104 615839
rect 42430 615496 42486 615505
rect 42430 615431 42486 615440
rect 42062 615224 42118 615233
rect 42118 615182 42380 615210
rect 42062 615159 42118 615168
rect 41878 614136 41934 614145
rect 41878 614071 41934 614080
rect 41892 613768 41920 614071
rect 42352 613135 42380 615182
rect 42182 613107 42380 613135
rect 42444 612490 42472 615431
rect 42182 612462 42472 612490
rect 42720 611017 42748 619783
rect 42996 612377 43024 807463
rect 43180 788225 43208 810727
rect 43166 788216 43222 788225
rect 43166 788151 43222 788160
rect 43166 766320 43222 766329
rect 43166 766255 43222 766264
rect 43180 753001 43208 766255
rect 43166 752992 43222 753001
rect 43166 752927 43222 752936
rect 43166 723616 43222 723625
rect 43166 723551 43222 723560
rect 43180 703497 43208 723551
rect 43166 703488 43222 703497
rect 43166 703423 43222 703432
rect 43166 679144 43222 679153
rect 43166 679079 43222 679088
rect 43180 662697 43208 679079
rect 43166 662688 43222 662697
rect 43166 662623 43222 662632
rect 43166 636304 43222 636313
rect 43166 636239 43222 636248
rect 43180 624073 43208 636239
rect 43166 624064 43222 624073
rect 43166 623999 43222 624008
rect 43364 613034 43392 933263
rect 43534 932104 43590 932113
rect 43534 932039 43590 932048
rect 43364 613006 43411 613034
rect 43383 612746 43411 613006
rect 43548 612950 43576 932039
rect 44086 892800 44142 892809
rect 44086 892735 44088 892744
rect 44140 892735 44142 892744
rect 44088 892706 44140 892712
rect 44086 891984 44142 891993
rect 44086 891919 44088 891928
rect 44140 891919 44142 891928
rect 44088 891890 44140 891896
rect 44454 816096 44510 816105
rect 44454 816031 44510 816040
rect 44270 814464 44326 814473
rect 44270 814399 44326 814408
rect 43902 809568 43958 809577
rect 43902 809503 43958 809512
rect 43718 806304 43774 806313
rect 43718 806239 43774 806248
rect 43536 612944 43588 612950
rect 43536 612886 43588 612892
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43732 612542 43760 806239
rect 43916 796249 43944 809503
rect 43902 796240 43958 796249
rect 43902 796175 43958 796184
rect 44284 771633 44312 814399
rect 44468 773265 44496 816031
rect 44652 815697 44680 941015
rect 47596 891993 47624 991714
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 48976 940137 49004 990082
rect 48962 940128 49018 940137
rect 48962 940063 49018 940072
rect 50356 939865 50384 993142
rect 54484 992928 54536 992934
rect 54484 992870 54536 992876
rect 51724 991636 51776 991642
rect 51724 991578 51776 991584
rect 51736 942313 51764 991578
rect 53288 990276 53340 990282
rect 53288 990218 53340 990224
rect 51722 942304 51778 942313
rect 51722 942239 51778 942248
rect 50342 939856 50398 939865
rect 50342 939791 50398 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44638 815688 44694 815697
rect 44638 815623 44694 815632
rect 44822 815280 44878 815289
rect 44822 815215 44878 815224
rect 44638 813648 44694 813657
rect 44638 813583 44694 813592
rect 44454 773256 44510 773265
rect 44454 773191 44510 773200
rect 44454 772032 44510 772041
rect 44454 771967 44510 771976
rect 44270 771624 44326 771633
rect 44270 771559 44326 771568
rect 44270 766728 44326 766737
rect 44270 766663 44326 766672
rect 44284 746745 44312 766663
rect 44270 746736 44326 746745
rect 44270 746671 44326 746680
rect 44270 729736 44326 729745
rect 44270 729671 44326 729680
rect 44284 729178 44312 729671
rect 44468 729337 44496 771967
rect 44652 771338 44680 813583
rect 44836 772449 44864 815215
rect 45006 810384 45062 810393
rect 45006 810319 45062 810328
rect 45020 789313 45048 810319
rect 45190 807936 45246 807945
rect 45190 807871 45246 807880
rect 45204 795025 45232 807871
rect 45190 795016 45246 795025
rect 45190 794951 45246 794960
rect 45006 789304 45062 789313
rect 45006 789239 45062 789248
rect 45098 772848 45154 772857
rect 45098 772783 45154 772792
rect 44822 772440 44878 772449
rect 44822 772375 44878 772384
rect 44652 771310 44956 771338
rect 44730 771216 44786 771225
rect 44730 771151 44786 771160
rect 44454 729328 44510 729337
rect 44454 729263 44510 729272
rect 44284 729150 44404 729178
rect 44178 722800 44234 722809
rect 44178 722735 44234 722744
rect 43902 721576 43958 721585
rect 43902 721511 43958 721520
rect 43916 711113 43944 721511
rect 43902 711104 43958 711113
rect 43902 711039 43958 711048
rect 44192 707713 44220 722735
rect 44178 707704 44234 707713
rect 44178 707639 44234 707648
rect 44376 686905 44404 729150
rect 44546 728920 44602 728929
rect 44546 728855 44602 728864
rect 44362 686896 44418 686905
rect 44362 686831 44418 686840
rect 44362 686488 44418 686497
rect 44362 686423 44418 686432
rect 44376 685930 44404 686423
rect 44560 686089 44588 728855
rect 44744 728521 44772 771151
rect 44928 770817 44956 771310
rect 44914 770808 44970 770817
rect 44914 770743 44970 770752
rect 44914 770400 44970 770409
rect 44914 770335 44970 770344
rect 44730 728512 44786 728521
rect 44730 728447 44786 728456
rect 44730 728104 44786 728113
rect 44730 728039 44786 728048
rect 44744 721754 44772 728039
rect 44928 727705 44956 770335
rect 45112 730153 45140 772783
rect 45282 764824 45338 764833
rect 45282 764759 45338 764768
rect 45296 753545 45324 764759
rect 45558 764280 45614 764289
rect 45558 764215 45614 764224
rect 45282 753536 45338 753545
rect 45282 753471 45338 753480
rect 45098 730144 45154 730153
rect 45098 730079 45154 730088
rect 44914 727696 44970 727705
rect 44914 727631 44970 727640
rect 45098 727288 45154 727297
rect 45098 727223 45154 727232
rect 44744 721726 44956 721754
rect 44730 721168 44786 721177
rect 44730 721103 44786 721112
rect 44546 686080 44602 686089
rect 44546 686015 44602 686024
rect 44376 685902 44588 685930
rect 44178 680368 44234 680377
rect 44178 680303 44234 680312
rect 44192 663513 44220 680303
rect 44362 679552 44418 679561
rect 44362 679487 44418 679496
rect 44376 664873 44404 679487
rect 44362 664864 44418 664873
rect 44362 664799 44418 664808
rect 44178 663504 44234 663513
rect 44178 663439 44234 663448
rect 44560 643657 44588 685902
rect 44744 653177 44772 721103
rect 44928 685273 44956 721726
rect 44914 685264 44970 685273
rect 44914 685199 44970 685208
rect 45112 684457 45140 727223
rect 45374 685672 45430 685681
rect 45374 685607 45430 685616
rect 45388 685522 45416 685607
rect 45388 685494 45508 685522
rect 45282 684856 45338 684865
rect 45282 684791 45338 684800
rect 45098 684448 45154 684457
rect 45098 684383 45154 684392
rect 44914 684040 44970 684049
rect 44914 683975 44970 683984
rect 44730 653168 44786 653177
rect 44730 653103 44786 653112
rect 44546 643648 44602 643657
rect 44546 643583 44602 643592
rect 44730 643376 44786 643385
rect 44730 643311 44786 643320
rect 44454 642560 44510 642569
rect 44454 642495 44510 642504
rect 43902 635352 43958 635361
rect 43902 635287 43958 635296
rect 43916 623393 43944 635287
rect 44270 633448 44326 633457
rect 44270 633383 44326 633392
rect 43902 623384 43958 623393
rect 43902 623319 43958 623328
rect 43994 614136 44050 614145
rect 43994 614071 44050 614080
rect 43720 612536 43772 612542
rect 43720 612478 43772 612484
rect 42982 612368 43038 612377
rect 42982 612303 43038 612312
rect 43580 612368 43636 612377
rect 43580 612303 43582 612312
rect 43634 612303 43636 612312
rect 43582 612274 43634 612280
rect 44008 611538 44036 614071
rect 44008 611522 44082 611538
rect 44008 611516 44094 611522
rect 44008 611510 44042 611516
rect 44042 611458 44094 611464
rect 44284 611266 44312 633383
rect 44468 630674 44496 642495
rect 44468 630646 44588 630674
rect 44284 611238 44419 611266
rect 42706 611008 42762 611017
rect 42706 610943 42762 610952
rect 44391 610910 44419 611238
rect 44379 610904 44431 610910
rect 44379 610846 44431 610852
rect 44560 605834 44588 630646
rect 44744 611354 44772 643311
rect 44928 641481 44956 683975
rect 45296 644474 45324 684791
rect 45480 659654 45508 685494
rect 45204 644446 45324 644474
rect 45388 659626 45508 659654
rect 45204 642297 45232 644446
rect 45388 643113 45416 659626
rect 45374 643104 45430 643113
rect 45374 643039 45430 643048
rect 45190 642288 45246 642297
rect 45190 642223 45246 642232
rect 44914 641472 44970 641481
rect 44914 641407 44970 641416
rect 45006 641200 45062 641209
rect 45006 641135 45062 641144
rect 45020 636426 45048 641135
rect 45374 640928 45430 640937
rect 45374 640863 45430 640872
rect 45190 636576 45246 636585
rect 45190 636511 45246 636520
rect 45020 636398 45140 636426
rect 44914 635760 44970 635769
rect 44914 635695 44970 635704
rect 44928 620129 44956 635695
rect 44914 620120 44970 620129
rect 44914 620055 44970 620064
rect 44468 605806 44588 605834
rect 44652 611326 44772 611354
rect 44652 605834 44680 611326
rect 44822 611008 44878 611017
rect 44822 610943 44824 610952
rect 44876 610943 44878 610952
rect 44824 610914 44876 610920
rect 44652 605806 44772 605834
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 44468 599729 44496 605806
rect 44744 600545 44772 605806
rect 44730 600536 44786 600545
rect 44730 600471 44786 600480
rect 44914 600128 44970 600137
rect 44914 600063 44970 600072
rect 44454 599720 44510 599729
rect 44454 599655 44510 599664
rect 44730 599312 44786 599321
rect 44730 599247 44786 599256
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 41050 596864 41106 596873
rect 41050 596799 41106 596808
rect 32402 595640 32458 595649
rect 32402 595575 32458 595584
rect 32416 585818 32444 595575
rect 36542 595232 36598 595241
rect 36542 595167 36598 595176
rect 35162 594416 35218 594425
rect 35162 594351 35218 594360
rect 35176 585954 35204 594351
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 32404 585812 32456 585818
rect 32404 585754 32456 585760
rect 36556 585206 36584 595167
rect 37922 594824 37978 594833
rect 37922 594759 37978 594768
rect 36544 585200 36596 585206
rect 37936 585177 37964 594759
rect 40682 593600 40738 593609
rect 40682 593535 40738 593544
rect 40500 592408 40552 592414
rect 40500 592350 40552 592356
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 36544 585142 36596 585148
rect 37922 585168 37978 585177
rect 37922 585103 37978 585112
rect 39960 584905 39988 590679
rect 40512 589665 40540 592350
rect 40498 589656 40554 589665
rect 40498 589591 40554 589600
rect 39946 584896 40002 584905
rect 39946 584831 40002 584840
rect 40696 584633 40724 593535
rect 41064 592074 41092 596799
rect 41234 596048 41290 596057
rect 41234 595983 41290 595992
rect 41248 594726 41276 595983
rect 41236 594720 41288 594726
rect 41236 594662 41288 594668
rect 41512 594720 41564 594726
rect 41512 594662 41564 594668
rect 41326 594008 41382 594017
rect 41326 593943 41382 593952
rect 41340 593434 41368 593943
rect 41328 593428 41380 593434
rect 41328 593370 41380 593376
rect 41052 592068 41104 592074
rect 41052 592010 41104 592016
rect 41524 585449 41552 594662
rect 41696 593428 41748 593434
rect 41748 593388 42840 593416
rect 41696 593370 41748 593376
rect 41878 592784 41934 592793
rect 41878 592719 41934 592728
rect 41892 592498 41920 592719
rect 41708 592470 41920 592498
rect 41708 592414 41736 592470
rect 41696 592408 41748 592414
rect 41696 592350 41748 592356
rect 41696 592068 41748 592074
rect 41748 592016 42288 592034
rect 41696 592010 42288 592016
rect 41708 592006 42288 592010
rect 41694 586120 41750 586129
rect 41694 586055 41750 586064
rect 41708 585954 41736 586055
rect 41696 585948 41748 585954
rect 41696 585890 41748 585896
rect 41878 585848 41934 585857
rect 41708 585818 41878 585834
rect 41696 585812 41878 585818
rect 41748 585806 41878 585812
rect 41878 585783 41934 585792
rect 41696 585754 41748 585760
rect 41510 585440 41566 585449
rect 41510 585375 41566 585384
rect 41420 585200 41472 585206
rect 41420 585142 41472 585148
rect 40682 584624 40738 584633
rect 40682 584559 40738 584568
rect 41432 584474 41460 585142
rect 42260 585018 42288 592006
rect 42522 586120 42578 586129
rect 42578 586078 42748 586106
rect 42522 586055 42578 586064
rect 42430 585848 42486 585857
rect 42486 585806 42656 585834
rect 42430 585783 42486 585792
rect 42260 584990 42564 585018
rect 42154 584896 42210 584905
rect 42210 584854 42380 584882
rect 42154 584831 42210 584840
rect 41432 584446 42288 584474
rect 42260 583454 42288 584446
rect 42182 583426 42288 583454
rect 42352 582263 42380 584854
rect 42182 582235 42380 582263
rect 42536 581618 42564 584990
rect 42182 581590 42564 581618
rect 42246 581496 42302 581505
rect 42246 581431 42302 581440
rect 42260 580975 42288 581431
rect 42182 580947 42288 580975
rect 42246 580816 42302 580825
rect 42246 580751 42302 580760
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42260 578626 42288 580751
rect 42430 580544 42486 580553
rect 42430 580479 42486 580488
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 41786 578232 41842 578241
rect 41786 578167 41842 578176
rect 41800 577932 41828 578167
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42444 577425 42472 580479
rect 42430 577416 42486 577425
rect 42430 577351 42486 577360
rect 42628 576994 42656 585806
rect 42076 576966 42656 576994
rect 42076 576708 42104 576966
rect 42246 576872 42302 576881
rect 42246 576807 42302 576816
rect 42260 574274 42288 576807
rect 42720 575906 42748 586078
rect 42812 579614 42840 593388
rect 42812 579586 42932 579614
rect 42720 575878 42840 575906
rect 42182 574246 42288 574274
rect 42812 574138 42840 575878
rect 42536 574110 42840 574138
rect 42154 573880 42210 573889
rect 42154 573815 42210 573824
rect 42168 573580 42196 573815
rect 42536 572982 42564 574110
rect 42706 573880 42762 573889
rect 42706 573815 42762 573824
rect 42720 573730 42748 573815
rect 42904 573730 42932 579586
rect 42720 573702 42932 573730
rect 42182 572954 42564 572982
rect 42062 572656 42118 572665
rect 42062 572591 42118 572600
rect 42076 572424 42104 572591
rect 42246 572248 42302 572257
rect 42246 572183 42302 572192
rect 42062 571024 42118 571033
rect 42062 570959 42118 570968
rect 42076 570588 42104 570959
rect 42260 569922 42288 572183
rect 42614 571976 42670 571985
rect 42614 571911 42670 571920
rect 42182 569894 42288 569922
rect 42628 569514 42656 571911
rect 42076 569486 42656 569514
rect 42076 569296 42104 569486
rect 42338 569256 42394 569265
rect 42338 569191 42394 569200
rect 42352 567194 42380 569191
rect 41524 567166 42380 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 41524 557598 41552 567166
rect 42062 558512 42118 558521
rect 42062 558447 42118 558456
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 41512 557592 41564 557598
rect 42076 557569 42104 558447
rect 41512 557534 41564 557540
rect 42062 557560 42118 557569
rect 42996 557534 43024 596935
rect 44454 591968 44510 591977
rect 44454 591903 44510 591912
rect 43442 590336 43498 590345
rect 43442 590271 43498 590280
rect 42062 557495 42118 557504
rect 42812 557506 43024 557534
rect 35806 554840 35862 554849
rect 42812 554826 42840 557506
rect 41708 554810 42840 554826
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 41696 554804 42840 554810
rect 35808 554746 35860 554752
rect 41748 554798 42840 554804
rect 41696 554746 41748 554752
rect 35622 554024 35678 554033
rect 35622 553959 35678 553968
rect 35636 553450 35664 553959
rect 35806 553616 35862 553625
rect 35806 553551 35808 553560
rect 35860 553551 35862 553560
rect 41696 553580 41748 553586
rect 35808 553522 35860 553528
rect 41696 553522 41748 553528
rect 41708 553466 41736 553522
rect 35624 553444 35676 553450
rect 41328 553444 41380 553450
rect 35624 553386 35676 553392
rect 40958 553408 41014 553417
rect 41708 553438 41920 553466
rect 41328 553386 41380 553392
rect 41892 553394 41920 553438
rect 40958 553343 41014 553352
rect 33782 551984 33838 551993
rect 33782 551919 33838 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 33796 543046 33824 551919
rect 40972 549794 41000 553343
rect 41340 553058 41368 553386
rect 41892 553366 42472 553394
rect 41694 553072 41750 553081
rect 41340 553030 41694 553058
rect 41694 553007 41750 553016
rect 41142 552800 41198 552809
rect 41142 552735 41198 552744
rect 41156 551834 41184 552735
rect 41326 552392 41382 552401
rect 41326 552327 41382 552336
rect 41340 552090 41368 552327
rect 41786 552120 41842 552129
rect 41328 552084 41380 552090
rect 41328 552026 41380 552032
rect 41604 552084 41656 552090
rect 41656 552064 41786 552072
rect 41656 552055 41842 552064
rect 41656 552044 41828 552055
rect 41604 552026 41656 552032
rect 41694 551848 41750 551857
rect 41156 551806 41694 551834
rect 41694 551783 41750 551792
rect 41326 551168 41382 551177
rect 41326 551103 41382 551112
rect 41340 550798 41368 551103
rect 41328 550792 41380 550798
rect 41328 550734 41380 550740
rect 41604 550792 41656 550798
rect 41656 550752 41828 550780
rect 41604 550734 41656 550740
rect 41800 550633 41828 550752
rect 41786 550624 41842 550633
rect 41786 550559 41842 550568
rect 42062 550216 42118 550225
rect 42062 550151 42118 550160
rect 41786 549944 41842 549953
rect 41524 549902 41786 549930
rect 40972 549766 41184 549794
rect 37096 547460 37148 547466
rect 37096 547402 37148 547408
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 37108 542366 37136 547402
rect 41156 547346 41184 549766
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41156 547318 41368 547346
rect 41340 546417 41368 547318
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 41524 545465 41552 549902
rect 41786 549879 41842 549888
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 42076 545737 42104 550151
rect 42062 545728 42118 545737
rect 42062 545663 42118 545672
rect 41510 545456 41566 545465
rect 41510 545391 41566 545400
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 37096 542360 37148 542366
rect 37096 542302 37148 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538438 42472 553366
rect 42982 552120 43038 552129
rect 42982 552055 43038 552064
rect 42798 550624 42854 550633
rect 42798 550559 42854 550568
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42168 538370 42196 538424
rect 42260 538410 42472 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42168 537798 42288 537826
rect 42168 537744 42196 537798
rect 42260 537758 42288 537798
rect 42628 537758 42656 540223
rect 42260 537730 42656 537758
rect 42522 537568 42578 537577
rect 42522 537503 42578 537512
rect 41786 537024 41842 537033
rect 41786 536959 41842 536968
rect 42154 537024 42210 537033
rect 42154 536959 42210 536968
rect 41800 536588 41828 536959
rect 42168 536738 42196 536959
rect 42168 536710 42288 536738
rect 42260 535378 42288 536710
rect 42182 535350 42288 535378
rect 41786 535256 41842 535265
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42536 534086 42564 537503
rect 42182 534058 42564 534086
rect 42154 533896 42210 533905
rect 42154 533831 42210 533840
rect 42168 533528 42196 533831
rect 42246 533216 42302 533225
rect 42246 533151 42302 533160
rect 42260 531162 42288 533151
rect 42522 532808 42578 532817
rect 42522 532743 42578 532752
rect 42168 531134 42288 531162
rect 42168 531045 42196 531134
rect 42536 530890 42564 532743
rect 42812 531314 42840 550559
rect 42996 533905 43024 552055
rect 43166 549536 43222 549545
rect 43166 549471 43222 549480
rect 42982 533896 43038 533905
rect 42982 533831 43038 533840
rect 43180 533225 43208 549471
rect 43166 533216 43222 533225
rect 43166 533151 43222 533160
rect 42352 530862 42564 530890
rect 42720 531286 42840 531314
rect 42352 530754 42380 530862
rect 42260 530726 42380 530754
rect 42260 530414 42288 530726
rect 42522 530632 42578 530641
rect 42182 530386 42288 530414
rect 42352 530590 42522 530618
rect 42154 530088 42210 530097
rect 42154 530023 42210 530032
rect 42168 529757 42196 530023
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42352 527626 42380 530590
rect 42522 530567 42578 530576
rect 42720 530097 42748 531286
rect 42706 530088 42762 530097
rect 42706 530023 42762 530032
rect 42614 529680 42670 529689
rect 42614 529615 42670 529624
rect 42168 527598 42380 527626
rect 42168 527340 42196 527598
rect 42628 526742 42656 529615
rect 42890 529136 42946 529145
rect 42182 526714 42656 526742
rect 42720 529094 42890 529122
rect 42720 526091 42748 529094
rect 42890 529071 42946 529080
rect 42182 526063 42748 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40958 425640 41014 425649
rect 40958 425575 41014 425584
rect 36542 424416 36598 424425
rect 36542 424351 36598 424360
rect 36556 415410 36584 424351
rect 40972 422226 41000 425575
rect 41340 424946 41368 425983
rect 41340 424918 41552 424946
rect 41326 424008 41382 424017
rect 41326 423943 41382 423952
rect 41340 423706 41368 423943
rect 41328 423700 41380 423706
rect 41328 423642 41380 423648
rect 40972 422198 41184 422226
rect 41156 418849 41184 422198
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 41524 415562 41552 424918
rect 41696 423700 41748 423706
rect 41748 423660 42840 423688
rect 41696 423642 41748 423648
rect 41970 422784 42026 422793
rect 41970 422719 42026 422728
rect 41786 421968 41842 421977
rect 41786 421903 41842 421912
rect 41800 418305 41828 421903
rect 41984 418577 42012 422719
rect 42430 419928 42486 419937
rect 42430 419863 42486 419872
rect 41970 418568 42026 418577
rect 41970 418503 42026 418512
rect 41786 418296 41842 418305
rect 41786 418231 41842 418240
rect 41524 415534 42380 415562
rect 36544 415404 36596 415410
rect 36544 415346 36596 415352
rect 41696 415404 41748 415410
rect 41696 415346 41748 415352
rect 41708 415290 41736 415346
rect 41708 415262 42288 415290
rect 42260 413114 42288 415262
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 412026 42380 415534
rect 42444 415394 42472 419863
rect 42444 415366 42564 415394
rect 42260 411998 42380 412026
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42260 411074 42288 411998
rect 42536 411913 42564 415366
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42288 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42182 407102 42656 407130
rect 42430 407008 42486 407017
rect 42430 406943 42486 406952
rect 42444 406518 42472 406943
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42628 405657 42656 407102
rect 42614 405648 42670 405657
rect 42614 405583 42670 405592
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42182 402138 42472 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42444 400217 42472 402138
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423660
rect 43074 423192 43130 423201
rect 43074 423127 43130 423136
rect 43088 402937 43116 423127
rect 43258 421152 43314 421161
rect 43258 421087 43314 421096
rect 43272 407833 43300 421087
rect 43258 407824 43314 407833
rect 43258 407759 43314 407768
rect 43074 402928 43130 402937
rect 43074 402863 43130 402872
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41340 387654 41552 387682
rect 41142 387152 41198 387161
rect 41142 387087 41144 387096
rect 41196 387087 41198 387096
rect 41144 387058 41196 387064
rect 41340 386753 41368 387654
rect 41524 386753 41552 387654
rect 41708 387122 41920 387138
rect 41696 387116 41920 387122
rect 41748 387110 41920 387116
rect 41696 387058 41748 387064
rect 41892 387025 41920 387110
rect 41878 387016 41934 387025
rect 41878 386951 41934 386960
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41512 382424 41564 382430
rect 41512 382366 41564 382372
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 37922 381440 37978 381449
rect 37922 381375 37978 381384
rect 33782 380216 33838 380225
rect 33782 380151 33838 380160
rect 28538 376544 28594 376553
rect 28538 376479 28594 376488
rect 28552 373289 28580 376479
rect 28538 373280 28594 373289
rect 28538 373215 28594 373224
rect 33796 371929 33824 380151
rect 35808 379704 35860 379710
rect 35808 379646 35860 379652
rect 35820 379409 35848 379646
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35820 375426 35848 376071
rect 35808 375420 35860 375426
rect 35808 375362 35860 375368
rect 37936 373318 37964 381375
rect 40052 376961 40080 382191
rect 40222 381032 40278 381041
rect 40222 380967 40278 380976
rect 40236 378554 40264 380967
rect 41524 379514 41552 382366
rect 41696 379704 41748 379710
rect 41748 379652 42840 379658
rect 41696 379646 42840 379652
rect 41708 379630 42840 379646
rect 41524 379486 42380 379514
rect 40224 378548 40276 378554
rect 40224 378490 40276 378496
rect 41696 378548 41748 378554
rect 41696 378490 41748 378496
rect 41708 378434 41736 378490
rect 41708 378406 42288 378434
rect 40038 376952 40094 376961
rect 40038 376887 40094 376896
rect 41694 375456 41750 375465
rect 41694 375391 41696 375400
rect 41748 375391 41750 375400
rect 41696 375362 41748 375368
rect 37924 373312 37976 373318
rect 41696 373312 41748 373318
rect 37924 373254 37976 373260
rect 41694 373280 41696 373289
rect 41748 373280 41750 373289
rect 41694 373215 41750 373224
rect 33782 371920 33838 371929
rect 33782 371855 33838 371864
rect 42260 369854 42288 378406
rect 42168 369826 42288 369854
rect 42168 369444 42196 369826
rect 41786 368520 41842 368529
rect 41786 368455 41842 368464
rect 41800 368249 41828 368455
rect 42352 367622 42380 379486
rect 42614 373280 42670 373289
rect 42614 373215 42670 373224
rect 42182 367594 42380 367622
rect 42430 367024 42486 367033
rect 42182 366968 42430 366975
rect 42182 366959 42486 366968
rect 42182 366947 42472 366959
rect 42628 365922 42656 373215
rect 42536 365894 42656 365922
rect 42338 365800 42394 365809
rect 42182 365758 42338 365786
rect 42338 365735 42394 365744
rect 42154 364984 42210 364993
rect 42154 364919 42210 364928
rect 42168 364548 42196 364919
rect 42536 364426 42564 365894
rect 42812 365809 42840 379630
rect 43456 379514 43484 590271
rect 44468 581097 44496 591903
rect 44454 581088 44510 581097
rect 44454 581023 44510 581032
rect 44744 556481 44772 599247
rect 44928 557297 44956 600063
rect 45112 598913 45140 636398
rect 45204 634814 45232 636511
rect 45388 634814 45416 640863
rect 45204 634786 45324 634814
rect 45388 634786 45508 634814
rect 45296 625297 45324 634786
rect 45282 625288 45338 625297
rect 45282 625223 45338 625232
rect 45480 612082 45508 634786
rect 45388 612054 45508 612082
rect 45098 598904 45154 598913
rect 45098 598839 45154 598848
rect 45098 598496 45154 598505
rect 45098 598431 45154 598440
rect 44914 557288 44970 557297
rect 44914 557223 44970 557232
rect 44730 556472 44786 556481
rect 44730 556407 44786 556416
rect 44638 556064 44694 556073
rect 44638 555999 44694 556008
rect 44362 554432 44418 554441
rect 44362 554367 44418 554376
rect 44178 549128 44234 549137
rect 44178 549063 44234 549072
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43640 379514 43668 547703
rect 43810 547088 43866 547097
rect 43810 547023 43866 547032
rect 43456 379486 43576 379514
rect 43640 379486 43760 379514
rect 43350 375456 43406 375465
rect 43350 375391 43406 375400
rect 42798 365800 42854 365809
rect 42798 365735 42854 365744
rect 42536 364398 42656 364426
rect 42430 364304 42486 364313
rect 42430 364239 42486 364248
rect 42444 363950 42472 364239
rect 42182 363922 42472 363950
rect 41786 363624 41842 363633
rect 41786 363559 41842 363568
rect 41800 363256 41828 363559
rect 42628 362794 42656 364398
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362766 42656 362794
rect 42536 362726 42564 362766
rect 42260 362698 42564 362726
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42168 359638 42288 359666
rect 42168 359584 42196 359638
rect 42260 359598 42288 359638
rect 42260 359570 42472 359598
rect 41786 359408 41842 359417
rect 41786 359343 41842 359352
rect 41800 358972 41828 359343
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42444 357377 42472 359570
rect 42430 357368 42486 357377
rect 42430 357303 42486 357312
rect 42062 356960 42118 356969
rect 42062 356895 42118 356904
rect 42076 356592 42104 356895
rect 42430 356144 42486 356153
rect 42430 356079 42486 356088
rect 42444 355926 42472 356079
rect 42182 355898 42472 355926
rect 43364 355881 43392 375391
rect 43350 355872 43406 355881
rect 43350 355807 43406 355816
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 43548 355314 43576 379486
rect 43732 355586 43760 379486
rect 43824 355722 43852 547023
rect 44192 537577 44220 549063
rect 44178 537568 44234 537577
rect 44178 537503 44234 537512
rect 44178 428496 44234 428505
rect 44178 428431 44234 428440
rect 43994 419520 44050 419529
rect 43994 419455 44050 419464
rect 44008 355858 44036 419455
rect 44192 385665 44220 428431
rect 44376 427281 44404 554367
rect 44652 428913 44680 555999
rect 45112 555665 45140 598431
rect 45388 598097 45416 612054
rect 45572 611930 45600 764215
rect 46216 756401 46244 870810
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 46386 763056 46442 763065
rect 46386 762991 46442 763000
rect 46202 756392 46258 756401
rect 46202 756327 46258 756336
rect 45742 676696 45798 676705
rect 45742 676631 45798 676640
rect 45560 611924 45612 611930
rect 45560 611866 45612 611872
rect 45756 611318 45784 676631
rect 46018 637800 46074 637809
rect 46018 637735 46074 637744
rect 46032 615641 46060 637735
rect 46202 637120 46258 637129
rect 46202 637055 46258 637064
rect 46216 618497 46244 637055
rect 46202 618488 46258 618497
rect 46202 618423 46258 618432
rect 46018 615632 46074 615641
rect 46018 615567 46074 615576
rect 46400 612406 46428 762991
rect 46938 719944 46994 719953
rect 46938 719879 46994 719888
rect 46388 612400 46440 612406
rect 46388 612342 46440 612348
rect 46952 611726 46980 719879
rect 47596 712201 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47582 712192 47638 712201
rect 47582 712127 47638 712136
rect 47214 677920 47270 677929
rect 47214 677855 47270 677864
rect 46940 611720 46992 611726
rect 46940 611662 46992 611668
rect 45744 611312 45796 611318
rect 45744 611254 45796 611260
rect 47228 611114 47256 677855
rect 48976 669361 49004 767314
rect 50356 730561 50384 805938
rect 53116 799105 53144 923238
rect 53300 892265 53328 990218
rect 54496 892537 54524 992870
rect 55864 991500 55916 991506
rect 55864 991442 55916 991448
rect 55876 892809 55904 991442
rect 95896 990282 95924 1001914
rect 96080 991778 96108 1002322
rect 97264 1002108 97316 1002114
rect 97264 1002050 97316 1002056
rect 97276 994537 97304 1002050
rect 97460 997257 97488 1002458
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 97446 997248 97502 997257
rect 97446 997183 97502 997192
rect 98656 994702 98684 1002594
rect 100298 1002552 100354 1002561
rect 100298 1002487 100300 1002496
rect 100352 1002487 100354 1002496
rect 100300 1002458 100352 1002464
rect 99102 1002416 99158 1002425
rect 99102 1002351 99104 1002360
rect 99156 1002351 99158 1002360
rect 99104 1002322 99156 1002328
rect 101126 1002280 101182 1002289
rect 98828 1002244 98880 1002250
rect 101126 1002215 101128 1002224
rect 98828 1002186 98880 1002192
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 98840 995897 98868 1002186
rect 99470 1002144 99526 1002153
rect 99470 1002079 99472 1002088
rect 99524 1002079 99526 1002088
rect 100024 1002108 100076 1002114
rect 99472 1002050 99524 1002056
rect 100024 1002050 100076 1002056
rect 99012 1001972 99064 1001978
rect 99012 1001914 99064 1001920
rect 99024 999190 99052 1001914
rect 99012 999184 99064 999190
rect 99012 999126 99064 999132
rect 100036 998442 100064 1002050
rect 101126 1002008 101182 1002017
rect 101126 1001943 101128 1001952
rect 101180 1001943 101182 1001952
rect 101128 1001914 101180 1001920
rect 100024 998436 100076 998442
rect 100024 998378 100076 998384
rect 98826 995888 98882 995897
rect 98826 995823 98882 995832
rect 101416 995353 101444 1006130
rect 101600 997694 101628 1006402
rect 103978 1006224 104034 1006233
rect 103978 1006159 103980 1006168
rect 104032 1006159 104034 1006168
rect 106002 1006224 106058 1006233
rect 106002 1006159 106004 1006168
rect 103980 1006130 104032 1006136
rect 106056 1006159 106058 1006168
rect 106004 1006130 106056 1006136
rect 102322 1006088 102378 1006097
rect 102322 1006023 102324 1006032
rect 102376 1006023 102378 1006032
rect 108486 1006088 108542 1006097
rect 108486 1006023 108488 1006032
rect 102324 1005994 102376 1006000
rect 108540 1006023 108542 1006032
rect 108488 1005994 108540 1006000
rect 102784 1005304 102836 1005310
rect 108856 1005304 108908 1005310
rect 102784 1005246 102836 1005252
rect 108854 1005272 108856 1005281
rect 108908 1005272 108910 1005281
rect 101954 1002688 102010 1002697
rect 101954 1002623 101956 1002632
rect 102008 1002623 102010 1002632
rect 101956 1002594 102008 1002600
rect 101588 997688 101640 997694
rect 101588 997630 101640 997636
rect 101402 995344 101458 995353
rect 101402 995279 101458 995288
rect 98644 994696 98696 994702
rect 98644 994638 98696 994644
rect 97262 994528 97318 994537
rect 97262 994463 97318 994472
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 990276 95936 990282
rect 95884 990218 95936 990224
rect 89628 986128 89680 986134
rect 89628 986070 89680 986076
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 986070
rect 102796 985998 102824 1005246
rect 108854 1005207 108910 1005216
rect 108486 1004728 108542 1004737
rect 106188 1004692 106240 1004698
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 103152 1003944 103204 1003950
rect 103150 1003912 103152 1003921
rect 103204 1003912 103206 1003921
rect 103150 1003847 103206 1003856
rect 105634 1002280 105690 1002289
rect 105634 1002215 105636 1002224
rect 105688 1002215 105690 1002224
rect 105636 1002186 105688 1002192
rect 103150 1002144 103206 1002153
rect 103150 1002079 103152 1002088
rect 103204 1002079 103206 1002088
rect 103152 1002050 103204 1002056
rect 104806 1002008 104862 1002017
rect 104176 1001966 104806 1001994
rect 104176 994838 104204 1001966
rect 104806 1001943 104862 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 104164 994832 104216 994838
rect 104164 994774 104216 994780
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1004634
rect 107658 1002416 107714 1002425
rect 107658 1002351 107660 1002360
rect 107712 1002351 107714 1002360
rect 109500 1002380 109552 1002386
rect 107660 1002322 107712 1002328
rect 109500 1002322 109552 1002328
rect 108026 1002280 108082 1002289
rect 107844 1002244 107896 1002250
rect 108026 1002215 108028 1002224
rect 107844 1002186 107896 1002192
rect 108080 1002215 108082 1002224
rect 108028 1002186 108080 1002192
rect 106830 1002144 106886 1002153
rect 106830 1002079 106832 1002088
rect 106884 1002079 106886 1002088
rect 107856 1002096 107884 1002186
rect 109040 1002108 109092 1002114
rect 107856 1002068 108160 1002096
rect 106832 1002050 106884 1002056
rect 107752 1001972 107804 1001978
rect 107752 1001914 107804 1001920
rect 107764 993206 107792 1001914
rect 107752 993200 107804 993206
rect 107752 993142 107804 993148
rect 108132 990146 108160 1002068
rect 109040 1002050 109092 1002056
rect 109052 993070 109080 1002050
rect 109512 997626 109540 1002322
rect 110420 1002244 110472 1002250
rect 110420 1002186 110472 1002192
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 997620 109552 997626
rect 109500 997562 109552 997568
rect 109040 993064 109092 993070
rect 109040 993006 109092 993012
rect 110432 991642 110460 1002186
rect 111800 1002108 111852 1002114
rect 111800 1002050 111852 1002056
rect 110420 991636 110472 991642
rect 110420 991578 110472 991584
rect 108120 990140 108172 990146
rect 108120 990082 108172 990088
rect 111812 986134 111840 1002050
rect 113836 997762 113864 1007354
rect 425518 1007176 425574 1007185
rect 425518 1007111 425520 1007120
rect 425572 1007111 425574 1007120
rect 425520 1007082 425572 1007088
rect 359738 1007040 359794 1007049
rect 359738 1006975 359740 1006984
rect 359792 1006975 359794 1006984
rect 371240 1007004 371292 1007010
rect 359740 1006946 359792 1006952
rect 371240 1006946 371292 1006952
rect 359370 1006904 359426 1006913
rect 359370 1006839 359372 1006848
rect 359424 1006839 359426 1006848
rect 367376 1006868 367428 1006874
rect 359372 1006810 359424 1006816
rect 367376 1006810 367428 1006816
rect 361394 1006768 361450 1006777
rect 161756 1006732 161808 1006738
rect 161756 1006674 161808 1006680
rect 164884 1006732 164936 1006738
rect 361394 1006703 361396 1006712
rect 164884 1006674 164936 1006680
rect 361448 1006703 361450 1006712
rect 361396 1006674 361448 1006680
rect 153750 1006632 153806 1006641
rect 145564 1006596 145616 1006602
rect 153750 1006567 153752 1006576
rect 145564 1006538 145616 1006544
rect 153804 1006567 153806 1006576
rect 157430 1006632 157486 1006641
rect 157430 1006567 157432 1006576
rect 153752 1006538 153804 1006544
rect 157484 1006567 157486 1006576
rect 157432 1006538 157484 1006544
rect 144276 1006324 144328 1006330
rect 144276 1006266 144328 1006272
rect 124864 1006188 124916 1006194
rect 124864 1006130 124916 1006136
rect 121736 997892 121788 997898
rect 121736 997834 121788 997840
rect 113824 997756 113876 997762
rect 113824 997698 113876 997704
rect 117136 997756 117188 997762
rect 117136 997698 117188 997704
rect 116124 997620 116176 997626
rect 116124 997562 116176 997568
rect 116136 996985 116164 997562
rect 117148 997257 117176 997698
rect 117134 997248 117190 997257
rect 117134 997183 117190 997192
rect 116122 996976 116178 996985
rect 116122 996911 116178 996920
rect 111800 986128 111852 986134
rect 111800 986070 111852 986076
rect 105846 983606 106228 983634
rect 121748 983634 121776 997834
rect 124876 995081 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 126256 996305 126284 1005994
rect 144000 998436 144052 998442
rect 144000 998378 144052 998384
rect 143816 997756 143868 997762
rect 143816 997698 143868 997704
rect 143828 997257 143856 997698
rect 143814 997248 143870 997257
rect 143814 997183 143870 997192
rect 143724 996940 143776 996946
rect 143724 996882 143776 996888
rect 143736 996826 143764 996882
rect 143644 996798 143764 996826
rect 126242 996296 126298 996305
rect 126242 996231 126298 996240
rect 140792 995858 140820 995860
rect 140780 995852 140832 995858
rect 140780 995794 140832 995800
rect 131854 995752 131910 995761
rect 131606 995710 131854 995738
rect 131854 995687 131910 995696
rect 132958 995752 133014 995761
rect 136730 995752 136786 995761
rect 133014 995710 133446 995738
rect 136482 995710 136730 995738
rect 132958 995687 133014 995696
rect 140410 995752 140466 995761
rect 140162 995710 140410 995738
rect 136730 995687 136786 995696
rect 143644 995738 143672 996798
rect 143816 996668 143868 996674
rect 143816 996610 143868 996616
rect 140410 995687 140466 995696
rect 143460 995710 143672 995738
rect 141790 995616 141846 995625
rect 141450 995574 141790 995602
rect 141790 995551 141846 995560
rect 137374 995480 137430 995489
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994838 128492 995452
rect 128452 994832 128504 994838
rect 128452 994774 128504 994780
rect 129108 994702 129136 995452
rect 129096 994696 129148 994702
rect 129096 994638 129148 994644
rect 129752 994566 129780 995452
rect 132144 994809 132172 995452
rect 132802 995438 133184 995466
rect 132406 995344 132462 995353
rect 132406 995279 132462 995288
rect 132130 994800 132186 994809
rect 132130 994735 132186 994744
rect 129740 994560 129792 994566
rect 129740 994502 129792 994508
rect 132420 994430 132448 995279
rect 132408 994424 132460 994430
rect 132408 994366 132460 994372
rect 133156 994129 133184 995438
rect 134892 994560 134944 994566
rect 134892 994502 134944 994508
rect 134904 994294 134932 994502
rect 135916 994401 135944 995452
rect 137126 995438 137374 995466
rect 137374 995415 137430 995424
rect 135902 994392 135958 994401
rect 135902 994327 135958 994336
rect 134892 994288 134944 994294
rect 134892 994230 134944 994236
rect 133142 994120 133198 994129
rect 133142 994055 133198 994064
rect 137560 993880 137612 993886
rect 137558 993848 137560 993857
rect 137612 993848 137614 993857
rect 137558 993783 137614 993792
rect 137756 993721 137784 995452
rect 138966 995438 139348 995466
rect 142646 995438 143028 995466
rect 139320 995058 139348 995438
rect 143000 995330 143028 995438
rect 143460 995330 143488 995710
rect 143000 995302 143488 995330
rect 139320 995030 139440 995058
rect 139214 994120 139270 994129
rect 139214 994055 139270 994064
rect 137742 993712 137798 993721
rect 137742 993647 137798 993656
rect 139228 993449 139256 994055
rect 139412 993993 139440 995030
rect 142114 994696 142166 994702
rect 142166 994644 142384 994650
rect 142114 994638 142384 994644
rect 142126 994622 142384 994638
rect 142158 994528 142214 994537
rect 141804 994486 142158 994514
rect 139398 993984 139454 993993
rect 139398 993919 139454 993928
rect 141804 993886 141832 994486
rect 142158 994463 142214 994472
rect 141974 994392 142030 994401
rect 141974 994327 142030 994336
rect 141988 994022 142016 994327
rect 142158 994256 142214 994265
rect 142158 994191 142214 994200
rect 141976 994016 142028 994022
rect 141976 993958 142028 993964
rect 141792 993880 141844 993886
rect 141792 993822 141844 993828
rect 142172 993721 142200 994191
rect 142356 994158 142384 994622
rect 142344 994152 142396 994158
rect 142344 994094 142396 994100
rect 142344 994016 142396 994022
rect 142344 993958 142396 993964
rect 142356 993721 142384 993958
rect 142158 993712 142214 993721
rect 142158 993647 142214 993656
rect 142342 993712 142398 993721
rect 142342 993647 142398 993656
rect 143828 993449 143856 996610
rect 144012 995858 144040 998378
rect 144288 995897 144316 1006266
rect 144736 1006188 144788 1006194
rect 144736 1006130 144788 1006136
rect 144748 1001894 144776 1006130
rect 144656 1001866 144776 1001894
rect 144656 996713 144684 1001866
rect 144828 997620 144880 997626
rect 144828 997562 144880 997568
rect 144840 996985 144868 997562
rect 144826 996976 144882 996985
rect 144826 996911 144882 996920
rect 144642 996704 144698 996713
rect 144642 996639 144698 996648
rect 144552 996532 144604 996538
rect 144552 996474 144604 996480
rect 144564 996305 144592 996474
rect 144550 996296 144606 996305
rect 144550 996231 144606 996240
rect 144274 995888 144330 995897
rect 144000 995852 144052 995858
rect 144274 995823 144330 995832
rect 144000 995794 144052 995800
rect 145576 994809 145604 1006538
rect 152922 1006496 152978 1006505
rect 145748 1006460 145800 1006466
rect 152922 1006431 152924 1006440
rect 145748 1006402 145800 1006408
rect 152976 1006431 152978 1006440
rect 158258 1006496 158314 1006505
rect 158258 1006431 158260 1006440
rect 152924 1006402 152976 1006408
rect 158312 1006431 158314 1006440
rect 158260 1006402 158312 1006408
rect 145562 994800 145618 994809
rect 145562 994735 145618 994744
rect 145760 993993 145788 1006402
rect 158626 1006360 158682 1006369
rect 158626 1006295 158628 1006304
rect 158680 1006295 158682 1006304
rect 158628 1006266 158680 1006272
rect 151266 1006224 151322 1006233
rect 151266 1006159 151268 1006168
rect 151320 1006159 151322 1006168
rect 152094 1006224 152150 1006233
rect 152094 1006159 152096 1006168
rect 151268 1006130 151320 1006136
rect 152148 1006159 152150 1006168
rect 160282 1006224 160338 1006233
rect 161768 1006194 161796 1006674
rect 162308 1006596 162360 1006602
rect 162308 1006538 162360 1006544
rect 162492 1006596 162544 1006602
rect 162492 1006538 162544 1006544
rect 162320 1006194 162348 1006538
rect 162504 1006330 162532 1006538
rect 162492 1006324 162544 1006330
rect 162492 1006266 162544 1006272
rect 160282 1006159 160284 1006168
rect 152096 1006130 152148 1006136
rect 160336 1006159 160338 1006168
rect 161756 1006188 161808 1006194
rect 160284 1006130 160336 1006136
rect 161756 1006130 161808 1006136
rect 162308 1006188 162360 1006194
rect 162308 1006130 162360 1006136
rect 147126 1006088 147182 1006097
rect 147126 1006023 147182 1006032
rect 148874 1006088 148930 1006097
rect 148874 1006023 148876 1006032
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145746 993984 145802 993993
rect 145746 993919 145802 993928
rect 139214 993440 139270 993449
rect 139214 993375 139270 993384
rect 143814 993440 143870 993449
rect 143814 993375 143870 993384
rect 138296 991636 138348 991642
rect 138296 991578 138348 991584
rect 121748 983606 122130 983634
rect 138308 983620 138336 991578
rect 146956 991506 146984 1001914
rect 147140 995625 147168 1006023
rect 148928 1006023 148930 1006032
rect 150070 1006088 150126 1006097
rect 158258 1006088 158314 1006097
rect 150070 1006023 150072 1006032
rect 148876 1005994 148928 1006000
rect 150124 1006023 150126 1006032
rect 153936 1006052 153988 1006058
rect 150072 1005994 150124 1006000
rect 158258 1006023 158260 1006032
rect 153936 1005994 153988 1006000
rect 158312 1006023 158314 1006032
rect 159454 1006088 159510 1006097
rect 159454 1006023 159456 1006032
rect 158260 1005994 158312 1006000
rect 159508 1006023 159510 1006032
rect 159456 1005994 159508 1006000
rect 152922 1005136 152978 1005145
rect 149888 1005100 149940 1005106
rect 152922 1005071 152924 1005080
rect 149888 1005042 149940 1005048
rect 152976 1005071 152978 1005080
rect 152924 1005042 152976 1005048
rect 149704 1004828 149756 1004834
rect 149704 1004770 149756 1004776
rect 148508 1002380 148560 1002386
rect 148508 1002322 148560 1002328
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 147126 995616 147182 995625
rect 147126 995551 147182 995560
rect 148336 992934 148364 1002050
rect 148520 994265 148548 1002322
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149060 996532 149112 996538
rect 149060 996474 149112 996480
rect 149072 994362 149100 996474
rect 149716 994634 149744 1004770
rect 149900 996674 149928 1005042
rect 153750 1005000 153806 1005009
rect 151084 1004964 151136 1004970
rect 153750 1004935 153752 1004944
rect 151084 1004906 151136 1004912
rect 153804 1004935 153806 1004944
rect 153752 1004906 153804 1004912
rect 150898 1002416 150954 1002425
rect 150898 1002351 150900 1002360
rect 150952 1002351 150954 1002360
rect 150900 1002322 150952 1002328
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 149888 996668 149940 996674
rect 149888 996610 149940 996616
rect 149704 994628 149756 994634
rect 149704 994570 149756 994576
rect 149060 994356 149112 994362
rect 149060 994298 149112 994304
rect 148506 994256 148562 994265
rect 148506 994191 148562 994200
rect 151096 994158 151124 1004906
rect 151726 1004864 151782 1004873
rect 151726 1004799 151728 1004808
rect 151780 1004799 151782 1004808
rect 151728 1004770 151780 1004776
rect 151268 1004692 151320 1004698
rect 151268 1004634 151320 1004640
rect 151280 996946 151308 1004634
rect 152464 1002108 152516 1002114
rect 152464 1002050 152516 1002056
rect 151268 996940 151320 996946
rect 151268 996882 151320 996888
rect 151084 994152 151136 994158
rect 151084 994094 151136 994100
rect 152476 993721 152504 1002050
rect 153948 997626 153976 1005994
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 160704 1004799 160706 1004808
rect 163136 1004828 163188 1004834
rect 160652 1004770 160704 1004776
rect 163136 1004770 163188 1004776
rect 154118 1004728 154174 1004737
rect 154118 1004663 154120 1004672
rect 154172 1004663 154174 1004672
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 154120 1004634 154172 1004640
rect 161164 1004663 161166 1004672
rect 162952 1004692 163004 1004698
rect 161112 1004634 161164 1004640
rect 162952 1004634 163004 1004640
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 157340 1002244 157392 1002250
rect 155776 1002186 155828 1002192
rect 157340 1002186 157392 1002192
rect 154578 1002144 154634 1002153
rect 154578 1002079 154580 1002088
rect 154632 1002079 154634 1002088
rect 154580 1002050 154632 1002056
rect 154946 1002008 155002 1002017
rect 154592 1001966 154946 1001994
rect 153936 997620 153988 997626
rect 153936 997562 153988 997568
rect 153016 996872 153068 996878
rect 153016 996814 153068 996820
rect 153028 994498 153056 996814
rect 154302 995752 154358 995761
rect 154302 995687 154358 995696
rect 154316 995081 154344 995687
rect 154302 995072 154358 995081
rect 154302 995007 154358 995016
rect 154592 994537 154620 1001966
rect 154946 1001943 155002 1001952
rect 155774 1002008 155830 1002017
rect 156602 1002008 156658 1002017
rect 155830 1001966 156000 1001994
rect 155774 1001943 155830 1001952
rect 155972 998442 156000 1001966
rect 156602 1001943 156604 1001952
rect 156656 1001943 156658 1001952
rect 156604 1001914 156656 1001920
rect 155960 998436 156012 998442
rect 155960 998378 156012 998384
rect 157352 994838 157380 1002186
rect 157798 1002144 157854 1002153
rect 157798 1002079 157800 1002088
rect 157852 1002079 157854 1002088
rect 160100 1002108 160152 1002114
rect 157800 1002050 157852 1002056
rect 160100 1002050 160152 1002056
rect 158720 1001972 158772 1001978
rect 158720 1001914 158772 1001920
rect 158732 996878 158760 1001914
rect 160112 997762 160140 1002050
rect 160100 997756 160152 997762
rect 160100 997698 160152 997704
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 158720 996872 158772 996878
rect 158720 996814 158772 996820
rect 157340 994832 157392 994838
rect 157340 994774 157392 994780
rect 154578 994528 154634 994537
rect 153016 994492 153068 994498
rect 154578 994463 154634 994472
rect 153016 994434 153068 994440
rect 152462 993712 152518 993721
rect 152462 993647 152518 993656
rect 148324 992928 148376 992934
rect 148324 992870 148376 992876
rect 146944 991500 146996 991506
rect 146944 991442 146996 991448
rect 160756 985726 160784 997154
rect 163148 991642 163176 1004770
rect 163136 991636 163188 991642
rect 163136 991578 163188 991584
rect 164896 990894 164924 1006674
rect 173164 1006596 173216 1006602
rect 173164 1006538 173216 1006544
rect 171784 1006460 171836 1006466
rect 171784 1006402 171836 1006408
rect 171796 996130 171824 1006402
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 169392 995988 169444 995994
rect 169392 995930 169444 995936
rect 171692 995988 171744 995994
rect 171692 995930 171744 995936
rect 169404 994226 169432 995930
rect 170680 995852 170732 995858
rect 170680 995794 170732 995800
rect 171232 995852 171284 995858
rect 171232 995794 171284 995800
rect 170496 994764 170548 994770
rect 170496 994706 170548 994712
rect 169392 994220 169444 994226
rect 169392 994162 169444 994168
rect 170508 993682 170536 994706
rect 170692 994498 170720 995794
rect 170864 995580 170916 995586
rect 170864 995522 170916 995528
rect 170876 994634 170904 995522
rect 171046 995208 171102 995217
rect 171046 995143 171102 995152
rect 171060 994770 171088 995143
rect 171244 995111 171272 995794
rect 171704 995335 171732 995930
rect 171692 995329 171744 995335
rect 171692 995271 171744 995277
rect 171508 995217 171560 995223
rect 171506 995208 171508 995217
rect 171560 995208 171562 995217
rect 171506 995143 171562 995152
rect 171232 995105 171284 995111
rect 173176 995081 173204 1006538
rect 256146 1006496 256202 1006505
rect 247868 1006460 247920 1006466
rect 307758 1006496 307814 1006505
rect 256146 1006431 256148 1006440
rect 247868 1006402 247920 1006408
rect 256200 1006431 256202 1006440
rect 301504 1006460 301556 1006466
rect 256148 1006402 256200 1006408
rect 307758 1006431 307760 1006440
rect 301504 1006402 301556 1006408
rect 307812 1006431 307814 1006440
rect 360566 1006496 360622 1006505
rect 360566 1006431 360568 1006440
rect 307760 1006402 307812 1006408
rect 360620 1006431 360622 1006440
rect 367008 1006460 367060 1006466
rect 360568 1006402 360620 1006408
rect 367008 1006402 367060 1006408
rect 210422 1006224 210478 1006233
rect 175924 1006188 175976 1006194
rect 210422 1006159 210424 1006168
rect 175924 1006130 175976 1006136
rect 210476 1006159 210478 1006168
rect 228364 1006188 228416 1006194
rect 210424 1006130 210476 1006136
rect 228364 1006130 228416 1006136
rect 175936 996033 175964 1006130
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 198188 1006052 198240 1006058
rect 201038 1006023 201040 1006032
rect 198188 1005994 198240 1006000
rect 201092 1006023 201094 1006032
rect 208398 1006088 208454 1006097
rect 208398 1006023 208400 1006032
rect 201040 1005994 201092 1006000
rect 208452 1006023 208454 1006032
rect 208400 1005994 208452 1006000
rect 175922 996024 175978 996033
rect 175922 995959 175978 995968
rect 177316 995353 177344 1005994
rect 195152 1001972 195204 1001978
rect 195152 1001914 195204 1001920
rect 195164 997121 195192 1001914
rect 195520 1001224 195572 1001230
rect 195520 1001166 195572 1001172
rect 195150 997112 195206 997121
rect 195150 997047 195206 997056
rect 195058 996840 195114 996849
rect 195058 996775 195114 996784
rect 188066 995752 188122 995761
rect 187864 995710 188066 995738
rect 189446 995752 189502 995761
rect 189152 995710 189446 995738
rect 188066 995687 188122 995696
rect 191746 995752 191802 995761
rect 191544 995710 191746 995738
rect 189446 995687 189502 995696
rect 192482 995752 192538 995761
rect 192188 995710 192482 995738
rect 191746 995687 191802 995696
rect 192482 995687 192538 995696
rect 195072 995625 195100 996775
rect 195244 996396 195296 996402
rect 195244 996338 195296 996344
rect 192298 995616 192354 995625
rect 194322 995616 194378 995625
rect 192354 995574 192832 995602
rect 194028 995574 194322 995602
rect 192298 995551 192354 995560
rect 194322 995551 194378 995560
rect 195058 995616 195114 995625
rect 195058 995551 195114 995560
rect 194876 995512 194928 995518
rect 179860 995438 180196 995466
rect 180504 995438 180748 995466
rect 181148 995438 181484 995466
rect 177302 995344 177358 995353
rect 177302 995279 177358 995288
rect 180168 995110 180196 995438
rect 180720 995382 180748 995438
rect 180708 995376 180760 995382
rect 180708 995318 180760 995324
rect 180156 995104 180208 995110
rect 171232 995047 171284 995053
rect 173162 995072 173218 995081
rect 180156 995046 180208 995052
rect 173162 995007 173218 995016
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 171048 994764 171100 994770
rect 171048 994706 171100 994712
rect 170864 994628 170916 994634
rect 170864 994570 170916 994576
rect 170680 994492 170732 994498
rect 170680 994434 170732 994440
rect 171244 993818 171272 994823
rect 181456 994022 181484 995438
rect 182974 995246 183002 995452
rect 183540 995438 183876 995466
rect 184184 995438 184520 995466
rect 184828 995438 184888 995466
rect 187312 995438 187648 995466
rect 188508 995438 188844 995466
rect 190348 995438 190592 995466
rect 194876 995454 194928 995460
rect 182962 995240 183014 995246
rect 182962 995182 183014 995188
rect 183848 994974 183876 995438
rect 183836 994968 183888 994974
rect 183836 994910 183888 994916
rect 184492 994022 184520 995438
rect 184860 994809 184888 995438
rect 184846 994800 184902 994809
rect 184846 994735 184902 994744
rect 186134 994392 186190 994401
rect 186502 994392 186558 994401
rect 186134 994327 186136 994336
rect 186188 994327 186190 994336
rect 186274 994356 186326 994362
rect 186136 994298 186188 994304
rect 186502 994327 186558 994336
rect 186274 994298 186326 994304
rect 186286 994242 186314 994298
rect 186148 994214 186314 994242
rect 186148 994022 186176 994214
rect 181444 994016 181496 994022
rect 184296 994016 184348 994022
rect 181444 993958 181496 993964
rect 184294 993984 184296 993993
rect 184480 994016 184532 994022
rect 184348 993984 184350 993993
rect 184480 993958 184532 993964
rect 186136 994016 186188 994022
rect 186274 994016 186326 994022
rect 186136 993958 186188 993964
rect 186272 993984 186274 993993
rect 186326 993984 186328 993993
rect 184294 993919 184350 993928
rect 186272 993919 186328 993928
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 170496 993676 170548 993682
rect 170496 993618 170548 993624
rect 164884 990888 164936 990894
rect 164884 990830 164936 990836
rect 170772 990888 170824 990894
rect 170772 990830 170824 990836
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 154500 983620 154528 985662
rect 170784 983620 170812 990830
rect 186516 983634 186544 994327
rect 187620 993886 187648 995438
rect 188816 994537 188844 995438
rect 188802 994528 188858 994537
rect 188802 994463 188858 994472
rect 187608 993880 187660 993886
rect 187422 993848 187478 993857
rect 187608 993822 187660 993828
rect 187422 993783 187424 993792
rect 187476 993783 187478 993792
rect 187424 993754 187476 993760
rect 190564 993546 190592 995438
rect 191104 994016 191156 994022
rect 190748 993964 191104 993970
rect 190748 993958 191156 993964
rect 190748 993942 191144 993958
rect 190748 993886 190776 993942
rect 190736 993880 190788 993886
rect 190736 993822 190788 993828
rect 194888 993546 194916 995454
rect 195256 993857 195284 996338
rect 195532 995518 195560 1001166
rect 196808 998708 196860 998714
rect 196808 998650 196860 998656
rect 196624 998572 196676 998578
rect 196624 998514 196676 998520
rect 195704 997824 195756 997830
rect 195704 997766 195756 997772
rect 195716 996169 195744 997766
rect 195702 996160 195758 996169
rect 195702 996095 195758 996104
rect 195520 995512 195572 995518
rect 195520 995454 195572 995460
rect 195518 995344 195574 995353
rect 195518 995279 195574 995288
rect 195532 994809 195560 995279
rect 195518 994800 195574 994809
rect 195518 994735 195574 994744
rect 195796 994356 195848 994362
rect 195796 994298 195848 994304
rect 195242 993848 195298 993857
rect 195808 993834 195836 994298
rect 196636 994265 196664 998514
rect 196622 994256 196678 994265
rect 196622 994191 196678 994200
rect 195808 993806 195974 993834
rect 195242 993783 195298 993792
rect 195946 993750 195974 993806
rect 196820 993750 196848 998650
rect 197360 998096 197412 998102
rect 197360 998038 197412 998044
rect 195934 993744 195986 993750
rect 195934 993686 195986 993692
rect 196808 993744 196860 993750
rect 196808 993686 196860 993692
rect 197372 993682 197400 998038
rect 198004 997960 198056 997966
rect 198004 997902 198056 997908
rect 198016 996402 198044 997902
rect 198200 996441 198228 1005994
rect 204904 1005304 204956 1005310
rect 212080 1005304 212132 1005310
rect 204904 1005246 204956 1005252
rect 212078 1005272 212080 1005281
rect 212132 1005272 212134 1005281
rect 203340 1002244 203392 1002250
rect 203340 1002186 203392 1002192
rect 202694 1002008 202750 1002017
rect 202694 1001943 202696 1001952
rect 202748 1001943 202750 1001952
rect 202696 1001914 202748 1001920
rect 200856 998368 200908 998374
rect 200856 998310 200908 998316
rect 200028 998232 200080 998238
rect 200028 998174 200080 998180
rect 200040 997801 200068 998174
rect 200672 997960 200724 997966
rect 200670 997928 200672 997937
rect 200724 997928 200726 997937
rect 200670 997863 200726 997872
rect 198738 997792 198794 997801
rect 198738 997727 198794 997736
rect 200026 997792 200082 997801
rect 200868 997754 200896 998310
rect 202696 998232 202748 998238
rect 202694 998200 202696 998209
rect 202748 998200 202750 998209
rect 202694 998135 202750 998144
rect 201868 998096 201920 998102
rect 201866 998064 201868 998073
rect 202328 998096 202380 998102
rect 201920 998064 201922 998073
rect 202328 998038 202380 998044
rect 201866 997999 201922 998008
rect 202144 997960 202196 997966
rect 202144 997902 202196 997908
rect 200026 997727 200082 997736
rect 198752 997121 198780 997727
rect 200776 997726 200896 997754
rect 198738 997112 198794 997121
rect 198738 997047 198794 997056
rect 200212 996872 200264 996878
rect 200210 996840 200212 996849
rect 200264 996840 200266 996849
rect 200210 996775 200266 996784
rect 198186 996432 198242 996441
rect 198004 996396 198056 996402
rect 198186 996367 198242 996376
rect 198004 996338 198056 996344
rect 200776 994537 200804 997726
rect 202156 994974 202184 997902
rect 202340 995382 202368 998038
rect 203352 997754 203380 1002186
rect 203708 1001972 203760 1001978
rect 203708 1001914 203760 1001920
rect 203522 998608 203578 998617
rect 203522 998543 203524 998552
rect 203576 998543 203578 998552
rect 203524 998514 203576 998520
rect 203524 998368 203576 998374
rect 203522 998336 203524 998345
rect 203576 998336 203578 998345
rect 203522 998271 203578 998280
rect 203352 997726 203564 997754
rect 202972 995920 203024 995926
rect 202970 995888 202972 995897
rect 203024 995888 203026 995897
rect 202970 995823 203026 995832
rect 203154 995888 203210 995897
rect 203154 995823 203210 995832
rect 202328 995376 202380 995382
rect 203168 995353 203196 995823
rect 202328 995318 202380 995324
rect 203154 995344 203210 995353
rect 203154 995279 203210 995288
rect 202144 994968 202196 994974
rect 202144 994910 202196 994916
rect 200762 994528 200818 994537
rect 200762 994463 200818 994472
rect 203536 994022 203564 997726
rect 203720 996878 203748 1001914
rect 203892 1001224 203944 1001230
rect 203890 1001192 203892 1001201
rect 203944 1001192 203946 1001201
rect 203890 1001127 203946 1001136
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 204720 997960 204772 997966
rect 204718 997928 204720 997937
rect 204772 997928 204774 997937
rect 204718 997863 204774 997872
rect 203708 996872 203760 996878
rect 203708 996814 203760 996820
rect 203524 994016 203576 994022
rect 203524 993958 203576 993964
rect 197360 993676 197412 993682
rect 197360 993618 197412 993624
rect 190552 993540 190604 993546
rect 190552 993482 190604 993488
rect 194876 993540 194928 993546
rect 194876 993482 194928 993488
rect 204916 986678 204944 1005246
rect 212078 1005207 212134 1005216
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 211250 1004864 211306 1004873
rect 211250 1004799 211252 1004808
rect 211304 1004799 211306 1004808
rect 211252 1004770 211304 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 211160 1004692 211212 1004698
rect 209228 1004634 209280 1004640
rect 211160 1004634 211212 1004640
rect 206374 1002280 206430 1002289
rect 206374 1002215 206376 1002224
rect 206428 1002215 206430 1002224
rect 206742 1002280 206798 1002289
rect 206742 1002215 206744 1002224
rect 206376 1002186 206428 1002192
rect 206796 1002215 206798 1002224
rect 208584 1002244 208636 1002250
rect 206744 1002186 206796 1002192
rect 208584 1002186 208636 1002192
rect 207202 1002144 207258 1002153
rect 205088 1002108 205140 1002114
rect 207202 1002079 207204 1002088
rect 205088 1002050 205140 1002056
rect 207256 1002079 207258 1002088
rect 207204 1002050 207256 1002056
rect 205100 995926 205128 1002050
rect 205546 1002008 205602 1002017
rect 206742 1002008 206798 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 206296 1001966 206742 1001994
rect 205548 1001914 205600 1001920
rect 205548 998096 205600 998102
rect 205546 998064 205548 998073
rect 205600 998064 205602 998073
rect 205546 997999 205602 998008
rect 205088 995920 205140 995926
rect 205088 995862 205140 995868
rect 206296 995110 206324 1001966
rect 207570 1002008 207626 1002017
rect 206742 1001943 206798 1001952
rect 207032 1001966 207570 1001994
rect 206284 995104 206336 995110
rect 206284 995046 206336 995052
rect 207032 993886 207060 1001966
rect 207570 1001943 207626 1001952
rect 208398 995888 208454 995897
rect 208398 995823 208454 995832
rect 208412 995081 208440 995823
rect 208596 995246 208624 1002186
rect 210882 1002144 210938 1002153
rect 210882 1002079 210884 1002088
rect 210936 1002079 210938 1002088
rect 210884 1002050 210936 1002056
rect 211172 996130 211200 1004634
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211816 995450 211844 1004906
rect 215944 1004828 215996 1004834
rect 215944 1004770 215996 1004776
rect 213184 1002108 213236 1002114
rect 213184 1002050 213236 1002056
rect 212538 1002008 212594 1002017
rect 212538 1001943 212540 1001952
rect 212592 1001943 212594 1001952
rect 212540 1001914 212592 1001920
rect 213196 995994 213224 1002050
rect 214564 1001972 214616 1001978
rect 214564 1001914 214616 1001920
rect 213184 995988 213236 995994
rect 213184 995930 213236 995936
rect 211804 995444 211856 995450
rect 211804 995386 211856 995392
rect 208584 995240 208636 995246
rect 208584 995182 208636 995188
rect 208398 995072 208454 995081
rect 208398 995007 208454 995016
rect 207020 993880 207072 993886
rect 207020 993822 207072 993828
rect 214576 991234 214604 1001914
rect 214564 991228 214616 991234
rect 214564 991170 214616 991176
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 204904 986672 204956 986678
rect 204904 986614 204956 986620
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1004770
rect 226340 997824 226392 997830
rect 226340 997766 226392 997772
rect 226352 994294 226380 997766
rect 228376 996130 228404 1006130
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 228364 996124 228416 996130
rect 228364 996066 228416 996072
rect 229756 995858 229784 1005994
rect 247316 1003944 247368 1003950
rect 247316 1003886 247368 1003892
rect 246580 1002584 246632 1002590
rect 246580 1002526 246632 1002532
rect 246592 997754 246620 1002526
rect 247132 999796 247184 999802
rect 247132 999738 247184 999744
rect 246764 998300 246816 998306
rect 246764 998242 246816 998248
rect 246500 997726 246620 997754
rect 229744 995852 229796 995858
rect 229744 995794 229796 995800
rect 234526 995752 234582 995761
rect 234416 995710 234526 995738
rect 234526 995687 234582 995696
rect 238574 995752 238630 995761
rect 240046 995752 240102 995761
rect 238630 995710 238740 995738
rect 239936 995710 240046 995738
rect 238574 995687 238630 995696
rect 243450 995752 243506 995761
rect 242972 995710 243450 995738
rect 240046 995687 240102 995696
rect 243818 995752 243874 995761
rect 243616 995710 243818 995738
rect 243450 995687 243506 995696
rect 243818 995687 243874 995696
rect 244094 995752 244150 995761
rect 244150 995710 244260 995738
rect 244094 995687 244150 995696
rect 240874 995616 240930 995625
rect 240580 995574 240874 995602
rect 240874 995551 240930 995560
rect 243266 995616 243322 995625
rect 243266 995551 243322 995560
rect 246212 995580 246264 995586
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 234968 995438 235304 995466
rect 235612 995438 235948 995466
rect 231596 995110 231624 995438
rect 231584 995104 231636 995110
rect 231584 995046 231636 995052
rect 232240 994974 232268 995438
rect 232228 994968 232280 994974
rect 232228 994910 232280 994916
rect 226340 994288 226392 994294
rect 226340 994230 226392 994236
rect 232884 994022 232912 995438
rect 235276 994809 235304 995438
rect 235920 995081 235948 995438
rect 236242 995246 236270 995452
rect 239292 995438 239628 995466
rect 241776 995438 242112 995466
rect 236230 995240 236282 995246
rect 236230 995182 236282 995188
rect 239600 995081 239628 995438
rect 242084 995353 242112 995438
rect 241886 995344 241942 995353
rect 241886 995279 241942 995288
rect 242070 995344 242126 995353
rect 242070 995279 242126 995288
rect 235906 995072 235962 995081
rect 235906 995007 235962 995016
rect 239586 995072 239642 995081
rect 239586 995007 239642 995016
rect 235262 994800 235318 994809
rect 235262 994735 235318 994744
rect 241900 994537 241928 995279
rect 243280 994838 243308 995551
rect 246212 995522 246264 995528
rect 245456 995438 245792 995466
rect 245764 995330 245792 995438
rect 246224 995330 246252 995522
rect 245764 995302 246252 995330
rect 246500 995081 246528 997726
rect 246776 995761 246804 998242
rect 246948 997552 247000 997558
rect 246948 997494 247000 997500
rect 246960 996985 246988 997494
rect 246946 996976 247002 996985
rect 246946 996911 247002 996920
rect 246762 995752 246818 995761
rect 246762 995687 246818 995696
rect 247144 995586 247172 999738
rect 247328 996033 247356 1003886
rect 247500 998436 247552 998442
rect 247500 998378 247552 998384
rect 247512 997257 247540 998378
rect 247684 997824 247736 997830
rect 247684 997766 247736 997772
rect 247498 997248 247554 997257
rect 247498 997183 247554 997192
rect 247314 996024 247370 996033
rect 247314 995959 247370 995968
rect 247132 995580 247184 995586
rect 247132 995522 247184 995528
rect 246486 995072 246542 995081
rect 246486 995007 246542 995016
rect 246670 995072 246726 995081
rect 246670 995007 246726 995016
rect 246684 994838 246712 995007
rect 243268 994832 243320 994838
rect 243268 994774 243320 994780
rect 246672 994832 246724 994838
rect 246672 994774 246724 994780
rect 243084 994764 243136 994770
rect 243084 994706 243136 994712
rect 241886 994528 241942 994537
rect 241886 994463 241942 994472
rect 232872 994016 232924 994022
rect 232872 993958 232924 993964
rect 243096 993886 243124 994706
rect 247696 993886 247724 997766
rect 247880 994537 247908 1006402
rect 258998 1006360 259054 1006369
rect 255964 1006324 256016 1006330
rect 258998 1006295 259000 1006304
rect 255964 1006266 256016 1006272
rect 259052 1006295 259054 1006304
rect 300492 1006324 300544 1006330
rect 259000 1006266 259052 1006272
rect 300492 1006266 300544 1006272
rect 252466 1006088 252522 1006097
rect 249064 1006052 249116 1006058
rect 252466 1006023 252522 1006032
rect 249064 1005994 249116 1006000
rect 248052 997688 248104 997694
rect 248052 997630 248104 997636
rect 248064 996713 248092 997630
rect 249076 997257 249104 1005994
rect 251824 1002380 251876 1002386
rect 251824 1002322 251876 1002328
rect 250628 998164 250680 998170
rect 250628 998106 250680 998112
rect 250444 997960 250496 997966
rect 250444 997902 250496 997908
rect 249062 997248 249118 997257
rect 249062 997183 249118 997192
rect 248050 996704 248106 996713
rect 248050 996639 248106 996648
rect 247866 994528 247922 994537
rect 250456 994498 250484 997902
rect 250640 995081 250668 998106
rect 251836 995246 251864 1002322
rect 252480 998306 252508 1006023
rect 255320 1003944 255372 1003950
rect 255318 1003912 255320 1003921
rect 255372 1003912 255374 1003921
rect 255318 1003847 255374 1003856
rect 253112 1002720 253164 1002726
rect 253112 1002662 253164 1002668
rect 252468 998300 252520 998306
rect 252468 998242 252520 998248
rect 252468 997824 252520 997830
rect 252466 997792 252468 997801
rect 252520 997792 252522 997801
rect 252466 997727 252522 997736
rect 251824 995240 251876 995246
rect 251824 995182 251876 995188
rect 250626 995072 250682 995081
rect 250626 995007 250682 995016
rect 253124 994809 253152 1002662
rect 254124 1002584 254176 1002590
rect 254122 1002552 254124 1002561
rect 254176 1002552 254178 1002561
rect 254122 1002487 254178 1002496
rect 254490 1002416 254546 1002425
rect 254490 1002351 254492 1002360
rect 254544 1002351 254546 1002360
rect 254492 1002322 254544 1002328
rect 254584 1002244 254636 1002250
rect 254584 1002186 254636 1002192
rect 253388 1002108 253440 1002114
rect 253388 1002050 253440 1002056
rect 253400 995353 253428 1002050
rect 253662 998200 253718 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 253664 998106 253716 998112
rect 253664 997960 253716 997966
rect 253662 997928 253664 997937
rect 253716 997928 253718 997937
rect 253662 997863 253718 997872
rect 253386 995344 253442 995353
rect 253386 995279 253442 995288
rect 254596 994974 254624 1002186
rect 255318 1002144 255374 1002153
rect 255318 1002079 255320 1002088
rect 255372 1002079 255374 1002088
rect 255320 1002050 255372 1002056
rect 254768 1001972 254820 1001978
rect 254768 1001914 254820 1001920
rect 254780 999802 254808 1001914
rect 254768 999796 254820 999802
rect 254768 999738 254820 999744
rect 255976 997558 256004 1006266
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 262732 1006159 262734 1006168
rect 269764 1006188 269816 1006194
rect 262680 1006130 262732 1006136
rect 269764 1006130 269816 1006136
rect 298744 1006188 298796 1006194
rect 298744 1006130 298796 1006136
rect 257342 1006088 257398 1006097
rect 257342 1006023 257344 1006032
rect 257396 1006023 257398 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 257344 1005994 257396 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 258170 1005136 258226 1005145
rect 257356 1005094 258170 1005122
rect 256148 1002720 256200 1002726
rect 256146 1002688 256148 1002697
rect 256200 1002688 256202 1002697
rect 256146 1002623 256202 1002632
rect 256514 1002280 256570 1002289
rect 256514 1002215 256516 1002224
rect 256568 1002215 256570 1002224
rect 256516 1002186 256568 1002192
rect 256974 1002008 257030 1002017
rect 256974 1001943 256976 1001952
rect 257028 1001943 257030 1001952
rect 256976 1001914 257028 1001920
rect 255964 997552 256016 997558
rect 255964 997494 256016 997500
rect 257356 995110 257384 1005094
rect 258170 1005071 258226 1005080
rect 263046 1005000 263102 1005009
rect 263046 1004935 263048 1004944
rect 263100 1004935 263102 1004944
rect 268384 1004964 268436 1004970
rect 263048 1004906 263100 1004912
rect 268384 1004906 268436 1004912
rect 258170 1004864 258226 1004873
rect 258170 1004799 258172 1004808
rect 258224 1004799 258226 1004808
rect 259460 1004828 259512 1004834
rect 258172 1004770 258224 1004776
rect 259460 1004770 259512 1004776
rect 258998 1002008 259054 1002017
rect 258092 1001966 258998 1001994
rect 257344 995104 257396 995110
rect 257344 995046 257396 995052
rect 254584 994968 254636 994974
rect 254584 994910 254636 994916
rect 253110 994800 253166 994809
rect 253110 994735 253166 994744
rect 247866 994463 247922 994472
rect 250444 994492 250496 994498
rect 250444 994434 250496 994440
rect 251456 994288 251508 994294
rect 251456 994230 251508 994236
rect 243084 993880 243136 993886
rect 243084 993822 243136 993828
rect 247684 993880 247736 993886
rect 247684 993822 247736 993828
rect 219440 991228 219492 991234
rect 219440 991170 219492 991176
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 991170
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 994230
rect 258092 994022 258120 1001966
rect 258998 1001943 259054 1001952
rect 259472 997694 259500 1004770
rect 261022 1002552 261078 1002561
rect 261022 1002487 261024 1002496
rect 261076 1002487 261078 1002496
rect 264244 1002516 264296 1002522
rect 261024 1002458 261076 1002464
rect 264244 1002458 264296 1002464
rect 260194 1002416 260250 1002425
rect 260194 1002351 260196 1002360
rect 260248 1002351 260250 1002360
rect 262864 1002380 262916 1002386
rect 260196 1002322 260248 1002328
rect 262864 1002322 262916 1002328
rect 259826 1002280 259882 1002289
rect 259826 1002215 259828 1002224
rect 259880 1002215 259882 1002224
rect 262220 1002244 262272 1002250
rect 259828 1002186 259880 1002192
rect 262220 1002186 262272 1002192
rect 261022 1002144 261078 1002153
rect 261022 1002079 261024 1002088
rect 261076 1002079 261078 1002088
rect 261024 1002050 261076 1002056
rect 260194 1002008 260250 1002017
rect 261850 1002008 261906 1002017
rect 260194 1001943 260196 1001952
rect 260248 1001943 260250 1001952
rect 260932 1001972 260984 1001978
rect 260196 1001914 260248 1001920
rect 260932 1001914 260984 1001920
rect 261128 1001966 261850 1001994
rect 259460 997688 259512 997694
rect 259460 997630 259512 997636
rect 260944 995450 260972 1001914
rect 261128 995994 261156 1001966
rect 261850 1001943 261906 1001952
rect 261116 995988 261168 995994
rect 261116 995930 261168 995936
rect 262232 995858 262260 1002186
rect 262876 996334 262904 1002322
rect 263506 1002144 263562 1002153
rect 263506 1002079 263508 1002088
rect 263560 1002079 263562 1002088
rect 263508 1002050 263560 1002056
rect 263874 1002008 263930 1002017
rect 263600 1001972 263652 1001978
rect 263874 1001943 263876 1001952
rect 263600 1001914 263652 1001920
rect 263928 1001943 263930 1001952
rect 263876 1001914 263928 1001920
rect 262864 996328 262916 996334
rect 262864 996270 262916 996276
rect 263612 996130 263640 1001914
rect 264256 996130 264284 1002458
rect 265624 1002108 265676 1002114
rect 265624 1002050 265676 1002056
rect 263600 996124 263652 996130
rect 263600 996066 263652 996072
rect 264244 996124 264296 996130
rect 264244 996066 264296 996072
rect 262220 995852 262272 995858
rect 262220 995794 262272 995800
rect 260932 995444 260984 995450
rect 260932 995386 260984 995392
rect 258080 994016 258132 994022
rect 258080 993958 258132 993964
rect 265636 990894 265664 1002050
rect 267004 1001972 267056 1001978
rect 267004 1001914 267056 1001920
rect 267016 991506 267044 1001914
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1004906
rect 269776 995994 269804 1006130
rect 279424 1006052 279476 1006058
rect 279424 1005994 279476 1006000
rect 279240 997756 279292 997762
rect 279240 997698 279292 997704
rect 270408 996328 270460 996334
rect 270408 996270 270460 996276
rect 269764 995988 269816 995994
rect 269764 995930 269816 995936
rect 270420 995081 270448 996270
rect 270406 995072 270462 995081
rect 270406 995007 270462 995016
rect 279252 994430 279280 997698
rect 279436 995353 279464 1005994
rect 298756 1001894 298784 1006130
rect 298928 1006052 298980 1006058
rect 298928 1005994 298980 1006000
rect 298756 1001866 298876 1001894
rect 298284 1000544 298336 1000550
rect 298284 1000486 298336 1000492
rect 298098 998880 298154 998889
rect 298098 998815 298154 998824
rect 298112 996033 298140 998815
rect 298098 996024 298154 996033
rect 298098 995959 298154 995968
rect 298296 995761 298324 1000486
rect 298650 997792 298706 997801
rect 298468 997756 298520 997762
rect 298650 997727 298706 997736
rect 298468 997698 298520 997704
rect 298480 996441 298508 997698
rect 298466 996432 298522 996441
rect 298466 996367 298522 996376
rect 282734 995752 282790 995761
rect 286782 995752 286838 995761
rect 282790 995710 282854 995738
rect 286534 995710 286782 995738
rect 282734 995687 282790 995696
rect 293590 995752 293646 995761
rect 293342 995710 293590 995738
rect 286782 995687 286838 995696
rect 295338 995752 295394 995761
rect 295182 995710 295338 995738
rect 293590 995687 293646 995696
rect 297270 995752 297326 995761
rect 297022 995710 297270 995738
rect 295338 995687 295394 995696
rect 297270 995687 297326 995696
rect 298282 995752 298338 995761
rect 298282 995687 298338 995696
rect 293222 995616 293278 995625
rect 293222 995551 293278 995560
rect 295522 995616 295578 995625
rect 295522 995551 295578 995560
rect 296902 995616 296958 995625
rect 298466 995616 298522 995625
rect 296902 995551 296958 995560
rect 297824 995580 297876 995586
rect 279422 995344 279478 995353
rect 279422 995279 279478 995288
rect 283484 995110 283512 995452
rect 283472 995104 283524 995110
rect 283472 995046 283524 995052
rect 284128 994974 284156 995452
rect 284116 994968 284168 994974
rect 284116 994910 284168 994916
rect 285968 994537 285996 995452
rect 285954 994528 286010 994537
rect 285954 994463 286010 994472
rect 279240 994424 279292 994430
rect 279240 994366 279292 994372
rect 287164 994265 287192 995452
rect 287808 994809 287836 995452
rect 290306 995438 290688 995466
rect 290660 995382 290688 995438
rect 290648 995376 290700 995382
rect 290648 995318 290700 995324
rect 290844 995246 290872 995452
rect 290832 995240 290884 995246
rect 290832 995182 290884 995188
rect 291488 994809 291516 995452
rect 287794 994800 287850 994809
rect 287794 994735 287850 994744
rect 291474 994800 291530 994809
rect 291474 994735 291530 994744
rect 292132 994265 292160 995452
rect 293236 994838 293264 995551
rect 293224 994832 293276 994838
rect 293224 994774 293276 994780
rect 294524 994294 294552 995452
rect 295536 995246 295564 995551
rect 295826 995438 296208 995466
rect 296180 995314 296208 995438
rect 296916 995330 296944 995551
rect 298466 995551 298522 995560
rect 297824 995522 297876 995528
rect 297836 995330 297864 995522
rect 296168 995308 296220 995314
rect 296916 995302 297864 995330
rect 296168 995250 296220 995256
rect 295524 995240 295576 995246
rect 295524 995182 295576 995188
rect 298480 994838 298508 995551
rect 298664 995314 298692 997727
rect 298652 995308 298704 995314
rect 298652 995250 298704 995256
rect 298468 994832 298520 994838
rect 298468 994774 298520 994780
rect 294512 994288 294564 994294
rect 287150 994256 287206 994265
rect 287150 994191 287206 994200
rect 292118 994256 292174 994265
rect 294512 994230 294564 994236
rect 292118 994191 292174 994200
rect 298848 994158 298876 1001866
rect 298940 997754 298968 1005994
rect 300308 1003332 300360 1003338
rect 300308 1003274 300360 1003280
rect 299386 1002280 299442 1002289
rect 299386 1002215 299442 1002224
rect 298940 997726 299060 997754
rect 299032 996130 299060 997726
rect 299204 997620 299256 997626
rect 299204 997562 299256 997568
rect 299216 996985 299244 997562
rect 299202 996976 299258 996985
rect 299202 996911 299258 996920
rect 299020 996124 299072 996130
rect 299020 996066 299072 996072
rect 299400 995586 299428 1002215
rect 300124 1002108 300176 1002114
rect 300124 1002050 300176 1002056
rect 299388 995580 299440 995586
rect 299388 995522 299440 995528
rect 300136 994634 300164 1002050
rect 300124 994628 300176 994634
rect 300124 994570 300176 994576
rect 300320 994265 300348 1003274
rect 300504 998889 300532 1006266
rect 300490 998880 300546 998889
rect 300490 998815 300546 998824
rect 301516 995625 301544 1006402
rect 306930 1006360 306986 1006369
rect 306930 1006295 306932 1006304
rect 306984 1006295 306986 1006304
rect 314658 1006360 314714 1006369
rect 314658 1006295 314660 1006304
rect 306932 1006266 306984 1006272
rect 314712 1006295 314714 1006304
rect 319444 1006324 319496 1006330
rect 314660 1006266 314712 1006272
rect 319444 1006266 319496 1006272
rect 354864 1006324 354916 1006330
rect 354864 1006266 354916 1006272
rect 360844 1006324 360896 1006330
rect 360844 1006266 360896 1006272
rect 304906 1006224 304962 1006233
rect 304906 1006159 304908 1006168
rect 304960 1006159 304962 1006168
rect 304908 1006130 304960 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301700 997801 301728 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311808 1006032
rect 304080 1005994 304132 1006000
rect 311860 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 314658 1006023 314660 1006032
rect 311808 1005994 311860 1006000
rect 314712 1006023 314714 1006032
rect 314660 1005994 314712 1006000
rect 307298 1005272 307354 1005281
rect 304264 1005236 304316 1005242
rect 307298 1005207 307300 1005216
rect 304264 1005178 304316 1005184
rect 307352 1005207 307354 1005216
rect 307300 1005178 307352 1005184
rect 302240 1002652 302292 1002658
rect 302240 1002594 302292 1002600
rect 301686 997792 301742 997801
rect 301686 997727 301742 997736
rect 302252 996713 302280 1002594
rect 303250 1002280 303306 1002289
rect 303250 1002215 303252 1002224
rect 303304 1002215 303306 1002224
rect 303252 1002186 303304 1002192
rect 304078 1002144 304134 1002153
rect 304078 1002079 304080 1002088
rect 304132 1002079 304134 1002088
rect 304080 1002050 304132 1002056
rect 302884 1001972 302936 1001978
rect 302884 1001914 302936 1001920
rect 302896 997257 302924 1001914
rect 302882 997248 302938 997257
rect 302882 997183 302938 997192
rect 302238 996704 302294 996713
rect 302238 996639 302294 996648
rect 301502 995616 301558 995625
rect 301502 995551 301558 995560
rect 304276 994537 304304 1005178
rect 308954 1005136 309010 1005145
rect 305828 1005100 305880 1005106
rect 308954 1005071 308956 1005080
rect 305828 1005042 305880 1005048
rect 309008 1005071 309010 1005080
rect 308956 1005042 309008 1005048
rect 305644 1004828 305696 1004834
rect 305644 1004770 305696 1004776
rect 304908 1004692 304960 1004698
rect 304908 1004634 304960 1004640
rect 304920 1002658 304948 1004634
rect 305274 1003368 305330 1003377
rect 305274 1003303 305276 1003312
rect 305328 1003303 305330 1003312
rect 305276 1003274 305328 1003280
rect 304908 1002652 304960 1002658
rect 304908 1002594 304960 1002600
rect 305656 995110 305684 1004770
rect 305840 1000550 305868 1005042
rect 308126 1004864 308182 1004873
rect 308126 1004799 308128 1004808
rect 308180 1004799 308182 1004808
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 308128 1004770 308180 1004776
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 306930 1004728 306986 1004737
rect 306930 1004663 306932 1004672
rect 306984 1004663 306986 1004672
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 306932 1004634 306984 1004640
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 310610 1002552 310666 1002561
rect 310610 1002487 310666 1002496
rect 310624 1002402 310652 1002487
rect 310440 1002374 310652 1002402
rect 306102 1002280 306158 1002289
rect 306102 1002215 306104 1002224
rect 306156 1002215 306158 1002224
rect 308404 1002244 308456 1002250
rect 306104 1002186 306156 1002192
rect 308404 1002186 308456 1002192
rect 306102 1002008 306158 1002017
rect 306102 1001943 306104 1001952
rect 306156 1001943 306158 1001952
rect 307024 1001972 307076 1001978
rect 306104 1001914 306156 1001920
rect 307024 1001914 307076 1001920
rect 305828 1000544 305880 1000550
rect 305828 1000486 305880 1000492
rect 307036 995246 307064 1001914
rect 307024 995240 307076 995246
rect 307024 995182 307076 995188
rect 305644 995104 305696 995110
rect 305644 995046 305696 995052
rect 308416 994974 308444 1002186
rect 308954 1002008 309010 1002017
rect 309782 1002008 309838 1002017
rect 308954 1001943 308956 1001952
rect 309008 1001943 309010 1001952
rect 309152 1001966 309782 1001994
rect 308956 1001914 309008 1001920
rect 308770 995616 308826 995625
rect 308770 995551 308826 995560
rect 308784 995081 308812 995551
rect 308770 995072 308826 995081
rect 308770 995007 308826 995016
rect 308404 994968 308456 994974
rect 308404 994910 308456 994916
rect 309152 994809 309180 1001966
rect 309782 1001943 309838 1001952
rect 310150 1002008 310206 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 310152 1001914 310204 1001920
rect 310440 1001894 310468 1002374
rect 310610 1002280 310666 1002289
rect 310610 1002215 310612 1002224
rect 310664 1002215 310666 1002224
rect 310612 1002186 310664 1002192
rect 311900 1001972 311952 1001978
rect 311900 1001914 311952 1001920
rect 310440 1001866 310560 1001894
rect 310532 997626 310560 1001866
rect 311912 997762 311940 1001914
rect 311900 997756 311952 997762
rect 311900 997698 311952 997704
rect 310520 997620 310572 997626
rect 310520 997562 310572 997568
rect 316052 995994 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316040 995988 316092 995994
rect 316040 995930 316092 995936
rect 309138 994800 309194 994809
rect 309138 994735 309194 994744
rect 304262 994528 304318 994537
rect 304262 994463 304318 994472
rect 316408 994424 316460 994430
rect 316408 994366 316460 994372
rect 300306 994256 300362 994265
rect 300306 994191 300362 994200
rect 298836 994152 298888 994158
rect 298836 994094 298888 994100
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994366
rect 318076 993070 318104 1004634
rect 318064 993064 318116 993070
rect 318064 993006 318116 993012
rect 319456 992934 319484 1006266
rect 354876 1006097 354904 1006266
rect 357714 1006224 357770 1006233
rect 357714 1006159 357716 1006168
rect 357768 1006159 357770 1006168
rect 357716 1006130 357768 1006136
rect 354862 1006088 354918 1006097
rect 320824 1006052 320876 1006058
rect 354862 1006023 354918 1006032
rect 355690 1006088 355746 1006097
rect 355690 1006023 355692 1006032
rect 320824 1005994 320876 1006000
rect 355744 1006023 355746 1006032
rect 359464 1006052 359516 1006058
rect 355692 1005994 355744 1006000
rect 359464 1005994 359516 1006000
rect 320836 997082 320864 1005994
rect 356520 1005304 356572 1005310
rect 356518 1005272 356520 1005281
rect 356572 1005272 356574 1005281
rect 356518 1005207 356574 1005216
rect 355690 1005000 355746 1005009
rect 353208 1004964 353260 1004970
rect 355690 1004935 355692 1004944
rect 353208 1004906 353260 1004912
rect 355744 1004935 355746 1004944
rect 355692 1004906 355744 1004912
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998578 351868 1001914
rect 353220 1001230 353248 1004906
rect 356518 1004864 356574 1004873
rect 354588 1004828 354640 1004834
rect 356518 1004799 356520 1004808
rect 354588 1004770 354640 1004776
rect 356572 1004799 356574 1004808
rect 356520 1004770 356572 1004776
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998572 351880 998578
rect 351828 998514 351880 998520
rect 320824 997076 320876 997082
rect 320824 997018 320876 997024
rect 332600 997076 332652 997082
rect 332600 997018 332652 997024
rect 319444 992928 319496 992934
rect 319444 992870 319496 992876
rect 332612 983634 332640 997018
rect 354600 995994 354628 1004770
rect 358542 1002280 358598 1002289
rect 355324 1002244 355376 1002250
rect 358542 1002215 358544 1002224
rect 355324 1002186 355376 1002192
rect 358596 1002215 358598 1002224
rect 358544 1002186 358596 1002192
rect 355336 998442 355364 1002186
rect 357714 1002144 357770 1002153
rect 355784 1002108 355836 1002114
rect 357714 1002079 357716 1002088
rect 355784 1002050 355836 1002056
rect 357768 1002079 357770 1002088
rect 357716 1002050 357768 1002056
rect 355324 998436 355376 998442
rect 355324 998378 355376 998384
rect 355796 997762 355824 1002050
rect 356886 1002008 356942 1002017
rect 356072 1001966 356886 1001994
rect 355784 997756 355836 997762
rect 355784 997698 355836 997704
rect 356072 997082 356100 1001966
rect 358542 1002008 358598 1002017
rect 356886 1001943 356942 1001952
rect 357452 1001966 358542 1001994
rect 357452 998714 357480 1001966
rect 358542 1001943 358598 1001952
rect 357440 998708 357492 998714
rect 357440 998650 357492 998656
rect 356060 997076 356112 997082
rect 356060 997018 356112 997024
rect 354588 995988 354640 995994
rect 354588 995930 354640 995936
rect 359476 995897 359504 1005994
rect 360568 1005440 360620 1005446
rect 360566 1005408 360568 1005417
rect 360620 1005408 360622 1005417
rect 360566 1005343 360622 1005352
rect 360198 1002008 360254 1002017
rect 360198 1001943 360200 1001952
rect 360252 1001943 360254 1001952
rect 360200 1001914 360252 1001920
rect 359462 995888 359518 995897
rect 359462 995823 359518 995832
rect 360856 994906 360884 1006266
rect 365074 1006224 365130 1006233
rect 362224 1006188 362276 1006194
rect 365074 1006159 365076 1006168
rect 362224 1006130 362276 1006136
rect 365128 1006159 365130 1006168
rect 365076 1006130 365128 1006136
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 362236 995314 362264 1006130
rect 363418 1006088 363474 1006097
rect 363418 1006023 363420 1006032
rect 363472 1006023 363474 1006032
rect 363420 1005994 363472 1006000
rect 367020 1005582 367048 1006402
rect 367388 1006330 367416 1006810
rect 367376 1006324 367428 1006330
rect 367376 1006266 367428 1006272
rect 367744 1006188 367796 1006194
rect 367744 1006130 367796 1006136
rect 367008 1005576 367060 1005582
rect 367008 1005518 367060 1005524
rect 365074 1005136 365130 1005145
rect 365074 1005071 365076 1005080
rect 365128 1005071 365130 1005080
rect 365076 1005042 365128 1005048
rect 364984 1004964 365036 1004970
rect 364984 1004906 365036 1004912
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 363604 1001972 363656 1001978
rect 363604 1001914 363656 1001920
rect 362224 995308 362276 995314
rect 362224 995250 362276 995256
rect 363616 995042 363644 1001914
rect 364996 995858 365024 1004906
rect 365168 1004828 365220 1004834
rect 365168 1004770 365220 1004776
rect 365180 997626 365208 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365168 997620 365220 997626
rect 365168 997562 365220 997568
rect 364984 995852 365036 995858
rect 364984 995794 365036 995800
rect 366376 995450 366404 1004634
rect 366364 995444 366416 995450
rect 366364 995386 366416 995392
rect 363604 995036 363656 995042
rect 363604 994978 363656 994984
rect 360844 994900 360896 994906
rect 360844 994842 360896 994848
rect 349160 993064 349212 993070
rect 349160 993006 349212 993012
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 993006
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 364996 983634 365024 992870
rect 367756 991506 367784 1006130
rect 370504 1005100 370556 1005106
rect 370504 1005042 370556 1005048
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 369136 991642 369164 1001914
rect 369124 991636 369176 991642
rect 369124 991578 369176 991584
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 370516 985998 370544 1005042
rect 371252 1002998 371280 1006946
rect 428372 1006936 428424 1006942
rect 428370 1006904 428372 1006913
rect 507860 1006936 507912 1006942
rect 428424 1006904 428426 1006913
rect 428370 1006839 428426 1006848
rect 507858 1006904 507860 1006913
rect 507912 1006904 507914 1006913
rect 507858 1006839 507914 1006848
rect 520924 1006868 520976 1006874
rect 520924 1006810 520976 1006816
rect 429200 1006800 429252 1006806
rect 429198 1006768 429200 1006777
rect 431868 1006800 431920 1006806
rect 429252 1006768 429254 1006777
rect 376024 1006732 376076 1006738
rect 431868 1006742 431920 1006748
rect 440240 1006800 440292 1006806
rect 440240 1006742 440292 1006748
rect 505006 1006768 505062 1006777
rect 429198 1006703 429254 1006712
rect 376024 1006674 376076 1006680
rect 373264 1005304 373316 1005310
rect 373264 1005246 373316 1005252
rect 371240 1002992 371292 1002998
rect 371240 1002934 371292 1002940
rect 372344 997756 372396 997762
rect 372344 997698 372396 997704
rect 372356 996713 372384 997698
rect 372528 997620 372580 997626
rect 372528 997562 372580 997568
rect 372540 996985 372568 997562
rect 372712 997076 372764 997082
rect 372712 997018 372764 997024
rect 372526 996976 372582 996985
rect 372526 996911 372582 996920
rect 372342 996704 372398 996713
rect 372342 996639 372398 996648
rect 372724 994770 372752 997018
rect 373276 996033 373304 1005246
rect 374368 1002992 374420 1002998
rect 374368 1002934 374420 1002940
rect 373262 996024 373318 996033
rect 373262 995959 373318 995968
rect 374380 995042 374408 1002934
rect 376036 998345 376064 1006674
rect 431684 1006664 431736 1006670
rect 431682 1006632 431684 1006641
rect 431736 1006632 431738 1006641
rect 431682 1006567 431738 1006576
rect 429198 1006496 429254 1006505
rect 402244 1006460 402296 1006466
rect 429198 1006431 429200 1006440
rect 402244 1006402 402296 1006408
rect 429252 1006431 429254 1006440
rect 429200 1006402 429252 1006408
rect 380164 1006324 380216 1006330
rect 380164 1006266 380216 1006272
rect 377404 1005576 377456 1005582
rect 377404 1005518 377456 1005524
rect 376022 998336 376078 998345
rect 376022 998271 376078 998280
rect 374368 995036 374420 995042
rect 374368 994978 374420 994984
rect 372712 994764 372764 994770
rect 372712 994706 372764 994712
rect 377416 994634 377444 1005518
rect 378784 1005440 378836 1005446
rect 378784 1005382 378836 1005388
rect 378796 998646 378824 1005382
rect 378784 998640 378836 998646
rect 378784 998582 378836 998588
rect 378600 998572 378652 998578
rect 378600 998514 378652 998520
rect 378612 998306 378640 998514
rect 378600 998300 378652 998306
rect 378600 998242 378652 998248
rect 380176 995586 380204 1006266
rect 382924 1006052 382976 1006058
rect 382924 1005994 382976 1006000
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 380912 996033 380940 1001166
rect 382280 998300 382332 998306
rect 382280 998242 382332 998248
rect 381542 996296 381598 996305
rect 381542 996231 381598 996240
rect 380898 996024 380954 996033
rect 381556 995994 381584 996231
rect 380898 995959 380954 995968
rect 381544 995988 381596 995994
rect 381544 995930 381596 995936
rect 382292 995761 382320 998242
rect 382936 996062 382964 1005994
rect 383292 998776 383344 998782
rect 383292 998718 383344 998724
rect 382924 996056 382976 996062
rect 382924 995998 382976 996004
rect 382278 995752 382334 995761
rect 382278 995687 382334 995696
rect 383304 995586 383332 998718
rect 383568 998640 383620 998646
rect 383620 998588 383700 998594
rect 383568 998582 383700 998588
rect 383580 998566 383700 998582
rect 383476 998436 383528 998442
rect 383476 998378 383528 998384
rect 380164 995580 380216 995586
rect 380164 995522 380216 995528
rect 383108 995580 383160 995586
rect 383108 995522 383160 995528
rect 383292 995580 383344 995586
rect 383292 995522 383344 995528
rect 377404 994628 377456 994634
rect 377404 994570 377456 994576
rect 383120 994498 383148 995522
rect 383488 995489 383516 998378
rect 383474 995480 383530 995489
rect 383474 995415 383530 995424
rect 383672 995330 383700 998566
rect 399944 997688 399996 997694
rect 399944 997630 399996 997636
rect 399956 996985 399984 997630
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 400876 995858 400904 1005994
rect 400864 995852 400916 995858
rect 400864 995794 400916 995800
rect 388718 995752 388774 995761
rect 388774 995710 389022 995738
rect 388718 995687 388774 995696
rect 384764 995580 384816 995586
rect 384764 995522 384816 995528
rect 385408 995580 385460 995586
rect 385408 995522 385460 995528
rect 386972 995580 387024 995586
rect 386972 995522 387024 995528
rect 384776 995466 384804 995522
rect 384316 995438 384698 995466
rect 384776 995438 385342 995466
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 384304 995172 384356 995178
rect 384304 995114 384356 995120
rect 384316 995024 384344 995114
rect 385420 995047 385448 995522
rect 384672 995036 384724 995042
rect 384316 994996 384672 995024
rect 384672 994978 384724 994984
rect 385406 995038 385462 995047
rect 385406 994973 385462 994982
rect 385972 994945 386000 995452
rect 386984 995330 387012 995522
rect 388166 995480 388222 995489
rect 386984 995302 387656 995330
rect 385958 994936 386014 994945
rect 387628 994922 387656 995302
rect 387812 995042 387840 995452
rect 392398 995480 392454 995489
rect 388222 995438 388378 995466
rect 389376 995438 389666 995466
rect 388166 995415 388222 995424
rect 389376 995042 389404 995438
rect 392136 995178 392164 995452
rect 393686 995480 393742 995489
rect 392454 995438 392702 995466
rect 392398 995415 392454 995424
rect 392124 995172 392176 995178
rect 392124 995114 392176 995120
rect 387800 995036 387852 995042
rect 387800 994978 387852 994984
rect 387984 995036 388036 995042
rect 387984 994978 388036 994984
rect 389364 995036 389416 995042
rect 389364 994978 389416 994984
rect 389548 995036 389600 995042
rect 389548 994978 389600 994984
rect 387996 994922 388024 994978
rect 387628 994894 388024 994922
rect 385958 994871 386014 994880
rect 389560 994498 389588 994978
rect 393332 994770 393360 995452
rect 396538 995480 396594 995489
rect 393742 995438 393990 995466
rect 394620 995438 395186 995466
rect 396382 995438 396538 995466
rect 393686 995415 393742 995424
rect 394620 995314 394648 995438
rect 396538 995415 396594 995424
rect 394608 995308 394660 995314
rect 394608 995250 394660 995256
rect 393320 994764 393372 994770
rect 393320 994706 393372 994712
rect 397012 994634 397040 995452
rect 397656 994770 397684 995452
rect 398852 995042 398880 995452
rect 402256 995450 402284 1006402
rect 431880 1006398 431908 1006742
rect 431868 1006392 431920 1006398
rect 423494 1006360 423550 1006369
rect 431868 1006334 431920 1006340
rect 423494 1006295 423496 1006304
rect 423548 1006295 423550 1006304
rect 429108 1006324 429160 1006330
rect 423496 1006266 423548 1006272
rect 429108 1006266 429160 1006272
rect 421838 1006088 421894 1006097
rect 421838 1006023 421894 1006032
rect 423494 1006088 423550 1006097
rect 423494 1006023 423496 1006032
rect 420828 1004828 420880 1004834
rect 420828 1004770 420880 1004776
rect 419448 1001972 419500 1001978
rect 419448 1001914 419500 1001920
rect 414478 996432 414534 996441
rect 414478 996367 414534 996376
rect 402244 995444 402296 995450
rect 402244 995386 402296 995392
rect 402796 995376 402848 995382
rect 402796 995318 402848 995324
rect 402980 995376 403032 995382
rect 402980 995318 403032 995324
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 402808 994770 402836 995318
rect 402992 994906 403020 995318
rect 402980 994900 403032 994906
rect 402980 994842 403032 994848
rect 397644 994764 397696 994770
rect 397644 994706 397696 994712
rect 402796 994764 402848 994770
rect 402796 994706 402848 994712
rect 397000 994628 397052 994634
rect 397000 994570 397052 994576
rect 383108 994492 383160 994498
rect 383108 994434 383160 994440
rect 389548 994492 389600 994498
rect 389548 994434 389600 994440
rect 414492 994294 414520 996367
rect 416134 995752 416190 995761
rect 416134 995687 416190 995696
rect 415398 995480 415454 995489
rect 415398 995415 415400 995424
rect 415452 995415 415454 995424
rect 415400 995386 415452 995392
rect 416148 995293 416176 995687
rect 416136 995287 416188 995293
rect 416136 995229 416188 995235
rect 419460 994702 419488 1001914
rect 420840 994974 420868 1004770
rect 421852 1003950 421880 1006023
rect 423548 1006023 423550 1006032
rect 423496 1005994 423548 1006000
rect 426348 1005712 426400 1005718
rect 426346 1005680 426348 1005689
rect 426400 1005680 426402 1005689
rect 426346 1005615 426402 1005624
rect 425520 1005576 425572 1005582
rect 425518 1005544 425520 1005553
rect 425572 1005544 425574 1005553
rect 425518 1005479 425574 1005488
rect 424324 1005440 424376 1005446
rect 424322 1005408 424324 1005417
rect 424376 1005408 424378 1005417
rect 424322 1005343 424378 1005352
rect 425152 1005304 425204 1005310
rect 425150 1005272 425152 1005281
rect 425204 1005272 425206 1005281
rect 425150 1005207 425206 1005216
rect 429120 1005174 429148 1006266
rect 431682 1006088 431738 1006097
rect 430304 1006052 430356 1006058
rect 431682 1006023 431684 1006032
rect 430304 1005994 430356 1006000
rect 431736 1006023 431738 1006032
rect 431684 1005994 431736 1006000
rect 429476 1005848 429528 1005854
rect 429476 1005790 429528 1005796
rect 429488 1005446 429516 1005790
rect 429476 1005440 429528 1005446
rect 429476 1005382 429528 1005388
rect 429108 1005168 429160 1005174
rect 429108 1005110 429160 1005116
rect 428004 1005032 428056 1005038
rect 428002 1005000 428004 1005009
rect 428056 1005000 428058 1005009
rect 428002 1004935 428058 1004944
rect 422666 1004864 422722 1004873
rect 422666 1004799 422668 1004808
rect 422720 1004799 422722 1004808
rect 422668 1004770 422720 1004776
rect 426348 1004080 426400 1004086
rect 426346 1004048 426348 1004057
rect 426400 1004048 426402 1004057
rect 426346 1003983 426402 1003992
rect 421840 1003944 421892 1003950
rect 421840 1003886 421892 1003892
rect 427174 1002144 427230 1002153
rect 427174 1002079 427230 1002088
rect 421470 1002008 421526 1002017
rect 424322 1002008 424378 1002017
rect 421470 1001943 421472 1001952
rect 421524 1001943 421526 1001952
rect 423588 1001972 423640 1001978
rect 421472 1001914 421524 1001920
rect 424322 1001943 424324 1001952
rect 423588 1001914 423640 1001920
rect 424376 1001943 424378 1001952
rect 424324 1001914 424376 1001920
rect 423600 1001230 423628 1001914
rect 423588 1001224 423640 1001230
rect 423588 1001166 423640 1001172
rect 427188 1000550 427216 1002079
rect 427544 1002040 427596 1002046
rect 427542 1002008 427544 1002017
rect 427596 1002008 427598 1002017
rect 427542 1001943 427598 1001952
rect 427176 1000544 427228 1000550
rect 427176 1000486 427228 1000492
rect 430316 999802 430344 1005994
rect 431868 1005848 431920 1005854
rect 431868 1005790 431920 1005796
rect 431880 1005038 431908 1005790
rect 431868 1005032 431920 1005038
rect 431868 1004974 431920 1004980
rect 432878 1004728 432934 1004737
rect 432878 1004663 432880 1004672
rect 432932 1004663 432934 1004672
rect 438124 1004692 438176 1004698
rect 432880 1004634 432932 1004640
rect 438124 1004634 438176 1004640
rect 431868 1002040 431920 1002046
rect 431868 1001982 431920 1001988
rect 430488 1000544 430540 1000550
rect 430488 1000486 430540 1000492
rect 430304 999796 430356 999802
rect 430304 999738 430356 999744
rect 428370 998880 428426 998889
rect 428370 998815 428372 998824
rect 428424 998815 428426 998824
rect 428372 998786 428424 998792
rect 430500 998714 430528 1000486
rect 430488 998708 430540 998714
rect 430488 998650 430540 998656
rect 430854 998608 430910 998617
rect 430854 998543 430856 998552
rect 430908 998543 430910 998552
rect 430856 998514 430908 998520
rect 431880 998442 431908 1001982
rect 436100 998844 436152 998850
rect 436100 998786 436152 998792
rect 436112 998578 436140 998786
rect 433984 998572 434036 998578
rect 433984 998514 434036 998520
rect 436100 998572 436152 998578
rect 436100 998514 436152 998520
rect 431868 998436 431920 998442
rect 431868 998378 431920 998384
rect 430026 998336 430082 998345
rect 430026 998271 430028 998280
rect 430080 998271 430082 998280
rect 432604 998300 432656 998306
rect 430028 998242 430080 998248
rect 432604 998242 432656 998248
rect 431222 998200 431278 998209
rect 431222 998135 431224 998144
rect 431276 998135 431278 998144
rect 431224 998106 431276 998112
rect 432050 998064 432106 998073
rect 432050 997999 432052 998008
rect 432104 997999 432106 998008
rect 432052 997970 432104 997976
rect 430028 997824 430080 997830
rect 430026 997792 430028 997801
rect 432052 997824 432104 997830
rect 430080 997792 430082 997801
rect 432052 997766 432104 997772
rect 430026 997727 430082 997736
rect 432064 997694 432092 997766
rect 432052 997688 432104 997694
rect 432052 997630 432104 997636
rect 432616 997626 432644 998242
rect 433524 998164 433576 998170
rect 433524 998106 433576 998112
rect 432604 997620 432656 997626
rect 432604 997562 432656 997568
rect 433536 996130 433564 998106
rect 433996 997762 434024 998514
rect 436744 998028 436796 998034
rect 436744 997970 436796 997976
rect 435362 997792 435418 997801
rect 433984 997756 434036 997762
rect 435362 997727 435418 997736
rect 433984 997698 434036 997704
rect 433524 996124 433576 996130
rect 433524 996066 433576 996072
rect 420828 994968 420880 994974
rect 420828 994910 420880 994916
rect 419448 994696 419500 994702
rect 419448 994638 419500 994644
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 414480 994288 414532 994294
rect 414480 994230 414532 994236
rect 370504 985992 370556 985998
rect 370504 985934 370556 985940
rect 381188 983634 381216 994230
rect 414112 991636 414164 991642
rect 414112 991578 414164 991584
rect 397828 985992 397880 985998
rect 397828 985934 397880 985940
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 985934
rect 414124 983620 414152 991578
rect 435376 991506 435404 997727
rect 430304 991500 430356 991506
rect 430304 991442 430356 991448
rect 435364 991500 435416 991506
rect 435364 991442 435416 991448
rect 430316 983620 430344 991442
rect 436756 985998 436784 997970
rect 438136 986134 438164 1004634
rect 440252 1002590 440280 1006742
rect 505006 1006703 505008 1006712
rect 505060 1006703 505062 1006712
rect 518164 1006732 518216 1006738
rect 505008 1006674 505060 1006680
rect 518164 1006674 518216 1006680
rect 501326 1006632 501382 1006641
rect 467104 1006596 467156 1006602
rect 501326 1006567 501328 1006576
rect 467104 1006538 467156 1006544
rect 501380 1006567 501382 1006576
rect 514760 1006596 514812 1006602
rect 501328 1006538 501380 1006544
rect 514760 1006538 514812 1006544
rect 453304 1005848 453356 1005854
rect 453304 1005790 453356 1005796
rect 445024 1005712 445076 1005718
rect 445024 1005654 445076 1005660
rect 440240 1002584 440292 1002590
rect 440240 1002526 440292 1002532
rect 440240 1001224 440292 1001230
rect 440240 1001166 440292 1001172
rect 439688 997756 439740 997762
rect 439688 997698 439740 997704
rect 439700 997257 439728 997698
rect 439872 997620 439924 997626
rect 439872 997562 439924 997568
rect 439686 997248 439742 997257
rect 439686 997183 439742 997192
rect 439884 996985 439912 997562
rect 440252 997218 440280 1001166
rect 443644 999796 443696 999802
rect 443644 999738 443696 999744
rect 440240 997212 440292 997218
rect 440240 997154 440292 997160
rect 443656 997082 443684 999738
rect 443644 997076 443696 997082
rect 443644 997018 443696 997024
rect 439870 996976 439926 996985
rect 439870 996911 439926 996920
rect 445036 996305 445064 1005654
rect 447784 1005168 447836 1005174
rect 447784 1005110 447836 1005116
rect 445668 997212 445720 997218
rect 445668 997154 445720 997160
rect 445022 996296 445078 996305
rect 445022 996231 445078 996240
rect 445680 994265 445708 997154
rect 447796 994537 447824 1005110
rect 453316 998850 453344 1005790
rect 457444 1005576 457496 1005582
rect 457444 1005518 457496 1005524
rect 455880 1004080 455932 1004086
rect 455880 1004022 455932 1004028
rect 453304 998844 453356 998850
rect 453304 998786 453356 998792
rect 453856 997076 453908 997082
rect 453856 997018 453908 997024
rect 453868 994838 453896 997018
rect 455892 995110 455920 1004022
rect 457456 998986 457484 1005518
rect 462964 1005440 463016 1005446
rect 462964 1005382 463016 1005388
rect 457444 998980 457496 998986
rect 457444 998922 457496 998928
rect 456800 998708 456852 998714
rect 456800 998650 456852 998656
rect 456812 995353 456840 998650
rect 462976 995625 463004 1005382
rect 464344 1003944 464396 1003950
rect 464344 1003886 464396 1003892
rect 462962 995616 463018 995625
rect 462962 995551 463018 995560
rect 456798 995344 456854 995353
rect 456798 995279 456854 995288
rect 455880 995104 455932 995110
rect 455880 995046 455932 995052
rect 453856 994832 453908 994838
rect 464356 994809 464384 1003886
rect 466368 1002584 466420 1002590
rect 466368 1002526 466420 1002532
rect 466380 996033 466408 1002526
rect 467116 998714 467144 1006538
rect 505374 1006360 505430 1006369
rect 505374 1006295 505376 1006304
rect 505428 1006295 505430 1006304
rect 505376 1006266 505428 1006272
rect 507030 1006224 507086 1006233
rect 469864 1006188 469916 1006194
rect 507030 1006159 507032 1006168
rect 469864 1006130 469916 1006136
rect 507084 1006159 507086 1006168
rect 509700 1006188 509752 1006194
rect 507032 1006130 507084 1006136
rect 509700 1006130 509752 1006136
rect 468484 1005304 468536 1005310
rect 468484 1005246 468536 1005252
rect 467104 998708 467156 998714
rect 467104 998650 467156 998656
rect 466366 996024 466422 996033
rect 466366 995959 466422 995968
rect 453856 994774 453908 994780
rect 464342 994800 464398 994809
rect 464342 994735 464398 994744
rect 447782 994528 447838 994537
rect 447782 994463 447838 994472
rect 468496 994430 468524 1005246
rect 469876 995081 469904 1006130
rect 498842 1006088 498898 1006097
rect 471244 1006052 471296 1006058
rect 471244 1005994 471296 1006000
rect 496728 1006052 496780 1006058
rect 498842 1006023 498844 1006032
rect 496728 1005994 496780 1006000
rect 498896 1006023 498898 1006032
rect 502522 1006088 502578 1006097
rect 506202 1006088 506258 1006097
rect 502522 1006023 502524 1006032
rect 498844 1005994 498896 1006000
rect 502576 1006023 502578 1006032
rect 505744 1006052 505796 1006058
rect 502524 1005994 502576 1006000
rect 506202 1006023 506204 1006032
rect 505744 1005994 505796 1006000
rect 506256 1006023 506258 1006032
rect 509054 1006088 509110 1006097
rect 509054 1006023 509056 1006032
rect 506204 1005994 506256 1006000
rect 509108 1006023 509110 1006032
rect 509240 1006052 509292 1006058
rect 509056 1005994 509108 1006000
rect 509240 1005994 509292 1006000
rect 471256 997754 471284 1005994
rect 472624 998980 472676 998986
rect 472624 998922 472676 998928
rect 472636 998866 472664 998922
rect 472440 998844 472492 998850
rect 472636 998838 472756 998866
rect 472440 998786 472492 998792
rect 472452 998730 472480 998786
rect 471980 998708 472032 998714
rect 472452 998702 472664 998730
rect 471980 998650 472032 998656
rect 471796 998436 471848 998442
rect 471796 998378 471848 998384
rect 471256 997726 471652 997754
rect 471150 996296 471206 996305
rect 471150 996231 471206 996240
rect 471164 995874 471192 996231
rect 471426 995888 471482 995897
rect 471164 995846 471426 995874
rect 471426 995823 471482 995832
rect 469862 995072 469918 995081
rect 469862 995007 469918 995016
rect 468484 994424 468536 994430
rect 468484 994366 468536 994372
rect 471624 994294 471652 997726
rect 446128 994288 446180 994294
rect 445666 994256 445722 994265
rect 446128 994230 446180 994236
rect 471612 994288 471664 994294
rect 471612 994230 471664 994236
rect 445666 994191 445722 994200
rect 438124 986128 438176 986134
rect 438124 986070 438176 986076
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 994230
rect 471808 994158 471836 998378
rect 471796 994152 471848 994158
rect 471796 994094 471848 994100
rect 471992 994022 472020 998650
rect 472440 998572 472492 998578
rect 472440 998514 472492 998520
rect 472452 995081 472480 998514
rect 472636 998458 472664 998702
rect 472544 998430 472664 998458
rect 472544 995330 472572 998430
rect 472728 995586 472756 998838
rect 489276 998096 489328 998102
rect 489276 998038 489328 998044
rect 493968 998096 494020 998102
rect 493968 998038 494020 998044
rect 489092 997756 489144 997762
rect 489092 997698 489144 997704
rect 488908 997620 488960 997626
rect 488908 997562 488960 997568
rect 488920 997257 488948 997562
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 489104 996985 489132 997698
rect 489090 996976 489146 996985
rect 489090 996911 489146 996920
rect 478326 995752 478382 995761
rect 473280 995710 473662 995738
rect 472716 995580 472768 995586
rect 472716 995522 472768 995528
rect 473280 995330 473308 995710
rect 478970 995752 479026 995761
rect 478382 995710 478630 995738
rect 478326 995687 478382 995696
rect 478970 995687 479026 995696
rect 485778 995752 485834 995761
rect 485834 995710 485990 995738
rect 485778 995687 485834 995696
rect 477682 995616 477738 995625
rect 474016 995586 474306 995602
rect 474004 995580 474306 995586
rect 474056 995574 474306 995580
rect 477738 995574 477986 995602
rect 477682 995551 477738 995560
rect 474004 995522 474056 995528
rect 478984 995518 479012 995687
rect 475936 995512 475988 995518
rect 472544 995302 473308 995330
rect 474752 995438 474950 995466
rect 475936 995454 475988 995460
rect 476396 995512 476448 995518
rect 476948 995512 477000 995518
rect 476448 995460 476790 995466
rect 476396 995454 476790 995460
rect 476948 995454 477000 995460
rect 478972 995512 479024 995518
rect 489288 995489 489316 998038
rect 489734 996704 489790 996713
rect 489734 996639 489790 996648
rect 489918 996704 489974 996713
rect 489918 996639 489974 996648
rect 485686 995480 485742 995489
rect 478972 995454 479024 995460
rect 474752 995081 474780 995438
rect 472254 995072 472310 995081
rect 472254 995007 472310 995016
rect 472438 995072 472494 995081
rect 472438 995007 472494 995016
rect 474738 995072 474794 995081
rect 474738 995007 474794 995016
rect 474922 995072 474978 995081
rect 474922 995007 474978 995016
rect 472268 994566 472296 995007
rect 474936 994566 474964 995007
rect 472256 994560 472308 994566
rect 472256 994502 472308 994508
rect 474924 994560 474976 994566
rect 474924 994502 474976 994508
rect 475948 994158 475976 995454
rect 476408 995438 476790 995454
rect 476960 995330 476988 995454
rect 476132 995302 476988 995330
rect 476132 995081 476160 995302
rect 476118 995072 476174 995081
rect 476118 995007 476174 995016
rect 476302 995072 476358 995081
rect 476302 995007 476358 995016
rect 476316 994294 476344 995007
rect 476304 994288 476356 994294
rect 476304 994230 476356 994236
rect 475936 994152 475988 994158
rect 475936 994094 475988 994100
rect 477328 994022 477356 995452
rect 480824 995438 481114 995466
rect 480824 995353 480852 995438
rect 480810 995344 480866 995353
rect 480810 995279 480866 995288
rect 481652 994566 481680 995452
rect 481928 995438 482310 995466
rect 481640 994560 481692 994566
rect 481640 994502 481692 994508
rect 481928 994265 481956 995438
rect 482940 994537 482968 995452
rect 482926 994528 482982 994537
rect 482926 994463 482982 994472
rect 484136 994430 484164 995452
rect 485346 995438 485686 995466
rect 489274 995480 489330 995489
rect 485686 995415 485742 995424
rect 486620 994809 486648 995452
rect 487816 995110 487844 995452
rect 489274 995415 489330 995424
rect 487804 995104 487856 995110
rect 487804 995046 487856 995052
rect 486606 994800 486662 994809
rect 486606 994735 486662 994744
rect 489748 994566 489776 996639
rect 489932 994838 489960 996639
rect 493980 995586 494008 998038
rect 493968 995580 494020 995586
rect 493968 995522 494020 995528
rect 496740 994838 496768 1005994
rect 498844 1005304 498896 1005310
rect 498842 1005272 498844 1005281
rect 498896 1005272 498898 1005281
rect 498842 1005207 498898 1005216
rect 500498 1005000 500554 1005009
rect 497924 1004964 497976 1004970
rect 500498 1004935 500500 1004944
rect 497924 1004906 497976 1004912
rect 500552 1004935 500554 1004944
rect 500500 1004906 500552 1004912
rect 497936 998442 497964 1004906
rect 499670 1004864 499726 1004873
rect 498108 1004828 498160 1004834
rect 499670 1004799 499672 1004808
rect 498108 1004770 498160 1004776
rect 499724 1004799 499726 1004808
rect 499672 1004770 499724 1004776
rect 498120 1001230 498148 1004770
rect 500498 1004728 500554 1004737
rect 499488 1004692 499540 1004698
rect 500498 1004663 500500 1004672
rect 499488 1004634 499540 1004640
rect 500552 1004663 500554 1004672
rect 500500 1004634 500552 1004640
rect 498108 1001224 498160 1001230
rect 498108 1001166 498160 1001172
rect 497924 998436 497976 998442
rect 497924 998378 497976 998384
rect 489920 994832 489972 994838
rect 489920 994774 489972 994780
rect 496728 994832 496780 994838
rect 496728 994774 496780 994780
rect 499500 994566 499528 1004634
rect 504546 1004456 504602 1004465
rect 504546 1004391 504548 1004400
rect 504600 1004391 504602 1004400
rect 504548 1004362 504600 1004368
rect 501694 1003368 501750 1003377
rect 501694 1003303 501696 1003312
rect 501748 1003303 501750 1003312
rect 504732 1003332 504784 1003338
rect 501696 1003274 501748 1003280
rect 504732 1003274 504784 1003280
rect 503350 1002416 503406 1002425
rect 503350 1002351 503352 1002360
rect 503404 1002351 503406 1002360
rect 503352 1002322 503404 1002328
rect 503350 1002144 503406 1002153
rect 503350 1002079 503352 1002088
rect 503404 1002079 503406 1002088
rect 503352 1002050 503404 1002056
rect 501694 1002008 501750 1002017
rect 500868 1001972 500920 1001978
rect 502522 1002008 502578 1002017
rect 501694 1001943 501696 1001952
rect 500868 1001914 500920 1001920
rect 501748 1001943 501750 1001952
rect 502156 1001972 502208 1001978
rect 501696 1001914 501748 1001920
rect 504178 1002008 504234 1002017
rect 502578 1001966 503024 1001994
rect 502522 1001943 502578 1001952
rect 502156 1001914 502208 1001920
rect 500880 998578 500908 1001914
rect 502168 998782 502196 1001914
rect 502156 998776 502208 998782
rect 502156 998718 502208 998724
rect 500868 998572 500920 998578
rect 500868 998514 500920 998520
rect 502996 997082 503024 1001966
rect 504178 1001943 504180 1001952
rect 504232 1001943 504234 1001952
rect 504180 1001914 504232 1001920
rect 504744 998986 504772 1003274
rect 505374 1002008 505430 1002017
rect 505374 1001943 505376 1001952
rect 505428 1001943 505430 1001952
rect 505376 1001914 505428 1001920
rect 504732 998980 504784 998986
rect 504732 998922 504784 998928
rect 502984 997076 503036 997082
rect 502984 997018 503036 997024
rect 489736 994560 489788 994566
rect 489736 994502 489788 994508
rect 499488 994560 499540 994566
rect 499488 994502 499540 994508
rect 505756 994430 505784 1005994
rect 509252 1005786 509280 1005994
rect 509240 1005780 509292 1005786
rect 509240 1005722 509292 1005728
rect 508226 1005136 508282 1005145
rect 508226 1005071 508228 1005080
rect 508280 1005071 508282 1005080
rect 508228 1005042 508280 1005048
rect 508226 1004864 508282 1004873
rect 508226 1004799 508228 1004808
rect 508280 1004799 508282 1004808
rect 508228 1004770 508280 1004776
rect 507398 1004728 507454 1004737
rect 507398 1004663 507400 1004672
rect 507452 1004663 507454 1004672
rect 509240 1004692 509292 1004698
rect 507400 1004634 507452 1004640
rect 509240 1004634 509292 1004640
rect 506480 1002380 506532 1002386
rect 506480 1002322 506532 1002328
rect 506296 1002108 506348 1002114
rect 506296 1002050 506348 1002056
rect 506308 998306 506336 1002050
rect 506492 999190 506520 1002322
rect 508504 1001972 508556 1001978
rect 508504 1001914 508556 1001920
rect 506480 999184 506532 999190
rect 506480 999126 506532 999132
rect 506296 998300 506348 998306
rect 506296 998242 506348 998248
rect 508516 997490 508544 1001914
rect 509252 997762 509280 1004634
rect 509712 997762 509740 1006130
rect 514024 1005780 514076 1005786
rect 514024 1005722 514076 1005728
rect 511264 1005100 511316 1005106
rect 511264 1005042 511316 1005048
rect 510804 1004828 510856 1004834
rect 510804 1004770 510856 1004776
rect 509882 1002144 509938 1002153
rect 509882 1002079 509884 1002088
rect 509936 1002079 509938 1002088
rect 509884 1002050 509936 1002056
rect 510342 1002008 510398 1002017
rect 510342 1001943 510344 1001952
rect 510396 1001943 510398 1001952
rect 510344 1001914 510396 1001920
rect 509240 997756 509292 997762
rect 509240 997698 509292 997704
rect 509700 997756 509752 997762
rect 509700 997698 509752 997704
rect 510816 997626 510844 1004770
rect 510988 1004420 511040 1004426
rect 510988 1004362 511040 1004368
rect 510804 997620 510856 997626
rect 510804 997562 510856 997568
rect 508504 997484 508556 997490
rect 508504 997426 508556 997432
rect 511000 997257 511028 1004362
rect 510986 997248 511042 997257
rect 510986 997183 511042 997192
rect 511276 996130 511304 1005042
rect 512644 1001972 512696 1001978
rect 512644 1001914 512696 1001920
rect 511264 996124 511316 996130
rect 511264 996066 511316 996072
rect 511080 995580 511132 995586
rect 511080 995522 511132 995528
rect 484124 994424 484176 994430
rect 484124 994366 484176 994372
rect 505744 994424 505796 994430
rect 505744 994366 505796 994372
rect 481914 994256 481970 994265
rect 481914 994191 481970 994200
rect 471980 994016 472032 994022
rect 471980 993958 472032 993964
rect 477316 994016 477368 994022
rect 477316 993958 477368 993964
rect 478972 991500 479024 991506
rect 478972 991442 479024 991448
rect 462780 986128 462832 986134
rect 462780 986070 462832 986076
rect 446140 983606 446522 983634
rect 462792 983620 462820 986070
rect 478984 983620 479012 991442
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 995522
rect 512656 990146 512684 1001914
rect 512644 990140 512696 990146
rect 512644 990082 512696 990088
rect 514036 985998 514064 1005722
rect 514772 999326 514800 1006538
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 515404 1002108 515456 1002114
rect 515404 1002050 515456 1002056
rect 514760 999320 514812 999326
rect 514760 999262 514812 999268
rect 515416 986134 515444 1002050
rect 516796 1001894 516824 1005246
rect 516796 1001866 517100 1001894
rect 516876 998776 516928 998782
rect 516876 998718 516928 998724
rect 516888 998617 516916 998718
rect 516874 998608 516930 998617
rect 516874 998543 516930 998552
rect 517072 998186 517100 1001866
rect 517428 999184 517480 999190
rect 517428 999126 517480 999132
rect 517244 998844 517296 998850
rect 517244 998786 517296 998792
rect 517256 998306 517284 998786
rect 517440 998714 517468 999126
rect 517704 998980 517756 998986
rect 517704 998922 517756 998928
rect 517428 998708 517480 998714
rect 517428 998650 517480 998656
rect 517520 998572 517572 998578
rect 517520 998514 517572 998520
rect 517244 998300 517296 998306
rect 517244 998242 517296 998248
rect 517072 998158 517284 998186
rect 517060 997756 517112 997762
rect 517060 997698 517112 997704
rect 516692 997484 516744 997490
rect 516692 997426 516744 997432
rect 516704 996441 516732 997426
rect 516876 997076 516928 997082
rect 516876 997018 516928 997024
rect 516690 996432 516746 996441
rect 516690 996367 516746 996376
rect 516888 995761 516916 997018
rect 517072 996985 517100 997698
rect 517058 996976 517114 996985
rect 517058 996911 517114 996920
rect 516874 995752 516930 995761
rect 516874 995687 516930 995696
rect 517256 993682 517284 998158
rect 517532 995353 517560 998514
rect 517518 995344 517574 995353
rect 517518 995279 517574 995288
rect 517716 995110 517744 998922
rect 518176 998306 518204 1006674
rect 519544 1006188 519596 1006194
rect 519544 1006130 519596 1006136
rect 518164 998300 518216 998306
rect 518164 998242 518216 998248
rect 517704 995104 517756 995110
rect 517704 995046 517756 995052
rect 519556 994430 519584 1006130
rect 520936 996033 520964 1006810
rect 555974 1006768 556030 1006777
rect 555974 1006703 555976 1006712
rect 556028 1006703 556030 1006712
rect 558828 1006732 558880 1006738
rect 555976 1006674 556028 1006680
rect 558828 1006674 558880 1006680
rect 556802 1006632 556858 1006641
rect 556802 1006567 556804 1006576
rect 556856 1006567 556858 1006576
rect 556804 1006538 556856 1006544
rect 553122 1006496 553178 1006505
rect 553122 1006431 553124 1006440
rect 553176 1006431 553178 1006440
rect 553124 1006402 553176 1006408
rect 552294 1006360 552350 1006369
rect 552294 1006295 552296 1006304
rect 552348 1006295 552350 1006304
rect 558184 1006324 558236 1006330
rect 552296 1006266 552348 1006272
rect 558184 1006266 558236 1006272
rect 551466 1006224 551522 1006233
rect 551466 1006159 551468 1006168
rect 551520 1006159 551522 1006168
rect 557448 1006188 557500 1006194
rect 551468 1006130 551520 1006136
rect 557448 1006130 557500 1006136
rect 551098 1006088 551154 1006097
rect 522304 1006052 522356 1006058
rect 551098 1006023 551154 1006032
rect 555974 1006088 556030 1006097
rect 555974 1006023 555976 1006032
rect 522304 1005994 522356 1006000
rect 521292 1001224 521344 1001230
rect 521292 1001166 521344 1001172
rect 520922 996024 520978 996033
rect 520922 995959 520978 995968
rect 519544 994424 519596 994430
rect 519544 994366 519596 994372
rect 521304 993818 521332 1001166
rect 522120 998844 522172 998850
rect 522120 998786 522172 998792
rect 522132 994158 522160 998786
rect 522316 995994 522344 1005994
rect 551112 1001366 551140 1006023
rect 556028 1006023 556030 1006032
rect 555976 1005994 556028 1006000
rect 552296 1005440 552348 1005446
rect 552294 1005408 552296 1005417
rect 552348 1005408 552350 1005417
rect 552294 1005343 552350 1005352
rect 551468 1005304 551520 1005310
rect 551466 1005272 551468 1005281
rect 551520 1005272 551522 1005281
rect 551466 1005207 551522 1005216
rect 557172 1003944 557224 1003950
rect 557170 1003912 557172 1003921
rect 557224 1003912 557226 1003921
rect 557170 1003847 557226 1003856
rect 553950 1002416 554006 1002425
rect 551928 1002380 551980 1002386
rect 553950 1002351 553952 1002360
rect 551928 1002322 551980 1002328
rect 554004 1002351 554006 1002360
rect 553952 1002322 554004 1002328
rect 551100 1001360 551152 1001366
rect 551100 1001302 551152 1001308
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 523500 999116 523552 999122
rect 523500 999058 523552 999064
rect 523512 996713 523540 999058
rect 523684 998708 523736 998714
rect 523684 998650 523736 998656
rect 523498 996704 523554 996713
rect 523498 996639 523554 996648
rect 522304 995988 522356 995994
rect 522304 995930 522356 995936
rect 523696 995330 523724 998650
rect 524052 998436 524104 998442
rect 524052 998378 524104 998384
rect 523868 998300 523920 998306
rect 523868 998242 523920 998248
rect 523880 995466 523908 998242
rect 524064 997257 524092 998378
rect 540888 997552 540940 997558
rect 540888 997494 540940 997500
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 540900 996985 540928 997494
rect 551940 997082 551968 1002322
rect 555146 1002280 555202 1002289
rect 553308 1002244 553360 1002250
rect 555146 1002215 555148 1002224
rect 553308 1002186 553360 1002192
rect 555200 1002215 555202 1002224
rect 555148 1002186 555200 1002192
rect 552664 1001972 552716 1001978
rect 552664 1001914 552716 1001920
rect 552676 997694 552704 1001914
rect 552664 997688 552716 997694
rect 552664 997630 552716 997636
rect 553320 997422 553348 1002186
rect 554318 1002008 554374 1002017
rect 554318 1001943 554320 1001952
rect 554372 1001943 554374 1001952
rect 554320 1001914 554372 1001920
rect 555148 999184 555200 999190
rect 555146 999152 555148 999161
rect 556160 999184 556212 999190
rect 555200 999152 555202 999161
rect 556160 999126 556212 999132
rect 555146 999087 555202 999096
rect 555424 998436 555476 998442
rect 555424 998378 555476 998384
rect 553952 997824 554004 997830
rect 553950 997792 553952 997801
rect 554004 997792 554006 997801
rect 553950 997727 554006 997736
rect 555436 997558 555464 998378
rect 555608 997824 555660 997830
rect 555608 997766 555660 997772
rect 555424 997552 555476 997558
rect 555424 997494 555476 997500
rect 553308 997416 553360 997422
rect 553308 997358 553360 997364
rect 555620 997218 555648 997766
rect 555608 997212 555660 997218
rect 555608 997154 555660 997160
rect 551928 997076 551980 997082
rect 551928 997018 551980 997024
rect 540886 996976 540942 996985
rect 540886 996911 540942 996920
rect 524050 996432 524106 996441
rect 524050 996367 524106 996376
rect 549442 996432 549498 996441
rect 549442 996367 549444 996376
rect 524064 995586 524092 996367
rect 549496 996367 549498 996376
rect 550640 996396 550692 996402
rect 549444 996338 549496 996344
rect 550640 996338 550692 996344
rect 529018 995752 529074 995761
rect 529662 995752 529718 995761
rect 529074 995710 529414 995738
rect 529018 995687 529074 995696
rect 529662 995687 529718 995696
rect 532238 995752 532294 995761
rect 532790 995752 532846 995761
rect 532294 995710 532542 995738
rect 532238 995687 532294 995696
rect 534630 995752 534686 995761
rect 532846 995710 533094 995738
rect 534382 995710 534630 995738
rect 532790 995687 532846 995696
rect 534630 995687 534686 995696
rect 536562 995752 536618 995761
rect 536618 995710 536774 995738
rect 538062 995710 538260 995738
rect 536562 995687 536618 995696
rect 526088 995586 526378 995602
rect 524052 995580 524104 995586
rect 524052 995522 524104 995528
rect 526076 995580 526378 995586
rect 526128 995574 526378 995580
rect 526076 995522 526128 995528
rect 523880 995438 524368 995466
rect 524340 995330 524368 995438
rect 524616 995438 525090 995466
rect 525168 995438 525734 995466
rect 527928 995438 528218 995466
rect 524616 995330 524644 995438
rect 525168 995330 525196 995438
rect 523696 995302 524276 995330
rect 524340 995302 524644 995330
rect 524708 995302 525196 995330
rect 524248 995194 524276 995302
rect 524708 995194 524736 995302
rect 524248 995166 524736 995194
rect 527928 995081 527956 995438
rect 527914 995072 527970 995081
rect 527914 995007 527970 995016
rect 528756 994294 528784 995452
rect 529676 995081 529704 995687
rect 529846 995616 529902 995625
rect 529902 995574 530058 995602
rect 529846 995551 529902 995560
rect 533724 995110 533752 995452
rect 535578 995438 535684 995466
rect 537418 995438 537800 995466
rect 535656 995353 535684 995438
rect 535642 995344 535698 995353
rect 535642 995279 535698 995288
rect 537772 995178 537800 995438
rect 537760 995172 537812 995178
rect 537760 995114 537812 995120
rect 533712 995104 533764 995110
rect 529662 995072 529718 995081
rect 533712 995046 533764 995052
rect 529662 995007 529718 995016
rect 538232 994838 538260 995710
rect 538404 995172 538456 995178
rect 538404 995114 538456 995120
rect 538220 994832 538272 994838
rect 538220 994774 538272 994780
rect 538416 994430 538444 995114
rect 538588 994560 538640 994566
rect 538586 994528 538588 994537
rect 538640 994528 538642 994537
rect 538586 994463 538642 994472
rect 538404 994424 538456 994430
rect 538404 994366 538456 994372
rect 539244 994294 539272 995452
rect 550652 994294 550680 996338
rect 556172 996334 556200 999126
rect 557460 998578 557488 1006130
rect 557448 998572 557500 998578
rect 557448 998514 557500 998520
rect 557998 998336 558054 998345
rect 557998 998271 558000 998280
rect 558052 998271 558054 998280
rect 558000 998242 558052 998248
rect 557998 998064 558054 998073
rect 557998 997999 558000 998008
rect 558052 997999 558054 998008
rect 558000 997970 558052 997976
rect 557630 997928 557686 997937
rect 557630 997863 557632 997872
rect 557684 997863 557686 997872
rect 557632 997834 557684 997840
rect 558196 997762 558224 1006266
rect 558840 1006194 558868 1006674
rect 567844 1006596 567896 1006602
rect 567844 1006538 567896 1006544
rect 558828 1006188 558880 1006194
rect 558828 1006130 558880 1006136
rect 566648 1005440 566700 1005446
rect 566648 1005382 566700 1005388
rect 560850 1004728 560906 1004737
rect 560850 1004663 560852 1004672
rect 560904 1004663 560906 1004672
rect 566464 1004692 566516 1004698
rect 560852 1004634 560904 1004640
rect 566464 1004634 566516 1004640
rect 560850 1002552 560906 1002561
rect 560850 1002487 560852 1002496
rect 560904 1002487 560906 1002496
rect 565084 1002516 565136 1002522
rect 560852 1002458 560904 1002464
rect 565084 1002458 565136 1002464
rect 560482 1002416 560538 1002425
rect 560482 1002351 560484 1002360
rect 560536 1002351 560538 1002360
rect 563060 1002380 563112 1002386
rect 560484 1002322 560536 1002328
rect 563060 1002322 563112 1002328
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 558826 998472 558882 998481
rect 558826 998407 558828 998416
rect 558880 998407 558882 998416
rect 558828 998378 558880 998384
rect 560944 998300 560996 998306
rect 560944 998242 560996 998248
rect 558826 998200 558882 998209
rect 558826 998135 558828 998144
rect 558880 998135 558882 998144
rect 558828 998106 558880 998112
rect 560300 998028 560352 998034
rect 560300 997970 560352 997976
rect 560022 997928 560078 997937
rect 559564 997892 559616 997898
rect 560022 997863 560024 997872
rect 559564 997834 559616 997840
rect 560076 997863 560078 997872
rect 560024 997834 560076 997840
rect 558184 997756 558236 997762
rect 558184 997698 558236 997704
rect 556160 996328 556212 996334
rect 556160 996270 556212 996276
rect 528744 994288 528796 994294
rect 528744 994230 528796 994236
rect 539232 994288 539284 994294
rect 539232 994230 539284 994236
rect 550640 994288 550692 994294
rect 550640 994230 550692 994236
rect 522120 994152 522172 994158
rect 522120 994094 522172 994100
rect 521292 993812 521344 993818
rect 521292 993754 521344 993760
rect 517244 993676 517296 993682
rect 517244 993618 517296 993624
rect 559576 991506 559604 997834
rect 560312 995994 560340 997970
rect 560300 995988 560352 995994
rect 560300 995930 560352 995936
rect 560956 992934 560984 998242
rect 562508 998164 562560 998170
rect 562508 998106 562560 998112
rect 562324 997892 562376 997898
rect 562324 997834 562376 997840
rect 562140 997620 562192 997626
rect 562140 997562 562192 997568
rect 562152 997354 562180 997562
rect 562140 997348 562192 997354
rect 562140 997290 562192 997296
rect 560944 992928 560996 992934
rect 560944 992870 560996 992876
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 562336 990146 562364 997834
rect 562520 993070 562548 998106
rect 562692 997756 562744 997762
rect 562692 997698 562744 997704
rect 562704 997490 562732 997698
rect 562692 997484 562744 997490
rect 562692 997426 562744 997432
rect 563072 996130 563100 1002322
rect 563704 1001972 563756 1001978
rect 563704 1001914 563756 1001920
rect 563060 996124 563112 996130
rect 563060 996066 563112 996072
rect 562508 993064 562560 993070
rect 562508 993006 562560 993012
rect 543832 990140 543884 990146
rect 543832 990082 543884 990088
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 515404 986128 515456 986134
rect 515404 986070 515456 986076
rect 527640 986128 527692 986134
rect 527640 986070 527692 986076
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 986070
rect 543844 983620 543872 990082
rect 563716 987426 563744 1001914
rect 563704 987420 563756 987426
rect 563704 987362 563756 987368
rect 565096 985998 565124 1002458
rect 566476 986134 566504 1004634
rect 566660 997762 566688 1005382
rect 566648 997756 566700 997762
rect 566648 997698 566700 997704
rect 567856 994838 567884 1006538
rect 570604 1006324 570656 1006330
rect 570604 1006266 570656 1006272
rect 569224 1005304 569276 1005310
rect 569224 1005246 569276 1005252
rect 568488 1001360 568540 1001366
rect 568488 1001302 568540 1001308
rect 568500 996946 568528 1001302
rect 568488 996940 568540 996946
rect 568488 996882 568540 996888
rect 567844 994832 567896 994838
rect 567844 994774 567896 994780
rect 569236 993954 569264 1005246
rect 570420 997212 570472 997218
rect 570420 997154 570472 997160
rect 570432 994809 570460 997154
rect 570616 996674 570644 1006266
rect 571984 1006188 572036 1006194
rect 571984 1006130 572036 1006136
rect 571248 1003944 571300 1003950
rect 571248 1003886 571300 1003892
rect 571064 996940 571116 996946
rect 571064 996882 571116 996888
rect 570604 996668 570656 996674
rect 570604 996610 570656 996616
rect 570418 994800 570474 994809
rect 570418 994735 570474 994744
rect 571076 994566 571104 996882
rect 571260 996810 571288 1003886
rect 571800 997620 571852 997626
rect 571800 997562 571852 997568
rect 571616 997484 571668 997490
rect 571616 997426 571668 997432
rect 571628 996946 571656 997426
rect 571812 997218 571840 997562
rect 571996 997490 572024 1006130
rect 573364 1006052 573416 1006058
rect 573364 1005994 573416 1006000
rect 572720 998436 572772 998442
rect 572720 998378 572772 998384
rect 571984 997484 572036 997490
rect 571984 997426 572036 997432
rect 571800 997212 571852 997218
rect 571800 997154 571852 997160
rect 571616 996940 571668 996946
rect 571616 996882 571668 996888
rect 571248 996804 571300 996810
rect 571248 996746 571300 996752
rect 572732 995110 572760 998378
rect 573376 996946 573404 1005994
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 572904 996940 572956 996946
rect 572904 996882 572956 996888
rect 573364 996940 573416 996946
rect 573364 996882 573416 996888
rect 572720 995104 572772 995110
rect 572720 995046 572772 995052
rect 571064 994560 571116 994566
rect 571064 994502 571116 994508
rect 572916 994430 572944 996882
rect 572904 994424 572956 994430
rect 572904 994366 572956 994372
rect 572720 994288 572772 994294
rect 572720 994230 572772 994236
rect 569224 993948 569276 993954
rect 569224 993890 569276 993896
rect 572732 990894 572760 994230
rect 574112 994090 574140 1001166
rect 618168 999184 618220 999190
rect 618168 999126 618220 999132
rect 625252 999184 625304 999190
rect 625252 999126 625304 999132
rect 591304 998096 591356 998102
rect 591304 998038 591356 998044
rect 591120 997960 591172 997966
rect 591120 997902 591172 997908
rect 590568 997212 590620 997218
rect 590568 997154 590620 997160
rect 590580 996985 590608 997154
rect 590566 996976 590622 996985
rect 591132 996946 591160 997902
rect 591316 997354 591344 998038
rect 592040 997824 592092 997830
rect 592040 997766 592092 997772
rect 592052 997490 592080 997766
rect 618180 997694 618208 999126
rect 618168 997688 618220 997694
rect 618168 997630 618220 997636
rect 592040 997484 592092 997490
rect 592040 997426 592092 997432
rect 591304 997348 591356 997354
rect 591304 997290 591356 997296
rect 623686 997248 623742 997257
rect 623686 997183 623742 997192
rect 623700 997082 623728 997183
rect 623688 997076 623740 997082
rect 623688 997018 623740 997024
rect 590566 996911 590622 996920
rect 591120 996940 591172 996946
rect 591120 996882 591172 996888
rect 590384 996804 590436 996810
rect 590384 996746 590436 996752
rect 590396 996690 590424 996746
rect 590566 996704 590622 996713
rect 590396 996662 590566 996690
rect 590566 996639 590622 996648
rect 590568 996464 590620 996470
rect 590566 996432 590568 996441
rect 590620 996432 590622 996441
rect 590566 996367 590622 996376
rect 590568 996260 590620 996266
rect 590568 996202 590620 996208
rect 590580 995081 590608 996202
rect 590750 995344 590806 995353
rect 590750 995279 590806 995288
rect 590566 995072 590622 995081
rect 590566 995007 590622 995016
rect 590764 994922 590792 995279
rect 590580 994894 590792 994922
rect 590580 994430 590608 994894
rect 625264 994430 625292 999126
rect 625620 998096 625672 998102
rect 625620 998038 625672 998044
rect 625436 997824 625488 997830
rect 625436 997766 625488 997772
rect 625448 996033 625476 997766
rect 625434 996024 625490 996033
rect 625434 995959 625490 995968
rect 625632 995761 625660 998038
rect 625804 997960 625856 997966
rect 625804 997902 625856 997908
rect 625618 995752 625674 995761
rect 625618 995687 625674 995696
rect 625816 995586 625844 997902
rect 627182 995752 627238 995761
rect 627918 995752 627974 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 629574 995752 629630 995761
rect 627974 995710 628176 995738
rect 627918 995687 627974 995696
rect 630310 995752 630366 995761
rect 629630 995710 630016 995738
rect 629574 995687 629630 995696
rect 633990 995752 634046 995761
rect 630366 995710 630568 995738
rect 630310 995687 630366 995696
rect 635278 995752 635334 995761
rect 634046 995710 634340 995738
rect 633990 995687 634046 995696
rect 637026 995752 637082 995761
rect 635334 995710 635536 995738
rect 635278 995687 635334 995696
rect 637082 995710 637376 995738
rect 637026 995687 637082 995696
rect 626552 995586 626888 995602
rect 625804 995580 625856 995586
rect 625804 995522 625856 995528
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 626540 995522 626592 995528
rect 630876 995438 631212 995466
rect 631520 995438 631856 995466
rect 634740 995438 634892 995466
rect 635844 995438 636180 995466
rect 638572 995438 638908 995466
rect 630876 994809 630904 995438
rect 630862 994800 630918 994809
rect 630862 994735 630918 994744
rect 631520 994430 631548 995438
rect 634740 995353 634768 995438
rect 634726 995344 634782 995353
rect 634726 995279 634782 995288
rect 635844 995110 635872 995438
rect 638880 995110 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640996 995438 641056 995466
rect 635832 995104 635884 995110
rect 635832 995046 635884 995052
rect 638868 995104 638920 995110
rect 638868 995046 638920 995052
rect 639064 994838 639092 995438
rect 639052 994832 639104 994838
rect 639052 994774 639104 994780
rect 639524 994566 639552 995438
rect 640800 995104 640852 995110
rect 640996 995081 641024 995438
rect 660304 995147 660356 995153
rect 660304 995089 660356 995095
rect 640800 995046 640852 995052
rect 640982 995072 641038 995081
rect 639512 994560 639564 994566
rect 639512 994502 639564 994508
rect 590568 994424 590620 994430
rect 590568 994366 590620 994372
rect 625252 994424 625304 994430
rect 625252 994366 625304 994372
rect 631508 994424 631560 994430
rect 631508 994366 631560 994372
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 572720 990888 572772 990894
rect 572720 990830 572772 990836
rect 576308 990888 576360 990894
rect 576308 990830 576360 990836
rect 566464 986128 566516 986134
rect 566464 986070 566516 986076
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 990830
rect 608784 987420 608836 987426
rect 608784 987362 608836 987368
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608796 983620 608824 987362
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 624988 983620 625016 985934
rect 640812 983634 640840 995046
rect 640982 995007 641038 995016
rect 660316 994702 660344 995089
rect 660304 994696 660356 994702
rect 660304 994638 660356 994644
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993682 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660960 993818 660988 994502
rect 660948 993812 661000 993818
rect 660948 993754 661000 993760
rect 660764 993676 660816 993682
rect 660764 993618 660816 993624
rect 660304 993064 660356 993070
rect 660304 993006 660356 993012
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 660316 937281 660344 993006
rect 667204 992928 667256 992934
rect 667204 992870 667256 992876
rect 664444 975724 664496 975730
rect 664444 975666 664496 975672
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660302 937272 660358 937281
rect 660302 937207 660358 937216
rect 661696 937038 661724 957743
rect 663064 948116 663116 948122
rect 663064 948058 663116 948064
rect 663076 941769 663104 948058
rect 664456 947345 664484 975666
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 664442 947336 664498 947345
rect 664442 947271 664498 947280
rect 663062 941760 663118 941769
rect 663062 941695 663118 941704
rect 665836 939865 665864 961862
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 667216 937825 667244 992870
rect 668584 990140 668636 990146
rect 668584 990082 668636 990088
rect 668596 938505 668624 990082
rect 675036 966709 675418 966737
rect 674378 966104 674434 966113
rect 674378 966039 674434 966048
rect 673366 962840 673422 962849
rect 673366 962775 673422 962784
rect 673182 962568 673238 962577
rect 673182 962503 673238 962512
rect 672998 958760 673054 958769
rect 672998 958695 673054 958704
rect 668582 938496 668638 938505
rect 668582 938431 668638 938440
rect 672170 938088 672226 938097
rect 672170 938023 672226 938032
rect 667202 937816 667258 937825
rect 667202 937751 667258 937760
rect 672184 937281 672212 938023
rect 672814 937816 672870 937825
rect 672814 937751 672870 937760
rect 672630 937544 672686 937553
rect 672630 937479 672686 937488
rect 672170 937272 672226 937281
rect 672170 937207 672226 937216
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 671802 936728 671858 936737
rect 671802 936663 671858 936672
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 671618 935776 671674 935785
rect 671618 935711 671674 935720
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 661684 921868 661736 921874
rect 661684 921810 661736 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 55862 892800 55918 892809
rect 55862 892735 55918 892744
rect 54482 892528 54538 892537
rect 54482 892463 54538 892472
rect 53286 892256 53342 892265
rect 53286 892191 53342 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62762 858664 62818 858673
rect 62762 858599 62818 858608
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799096 53158 799105
rect 53102 799031 53158 799040
rect 54496 774353 54524 844562
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 55876 772857 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62776 788633 62804 858599
rect 652390 856352 652446 856361
rect 652390 856287 652446 856296
rect 652404 855642 652432 856287
rect 652392 855636 652444 855642
rect 652392 855578 652444 855584
rect 652022 843024 652078 843033
rect 652022 842959 652078 842968
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 62946 793656 63002 793665
rect 62946 793591 63002 793600
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 55862 772848 55918 772857
rect 55862 772783 55918 772792
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 669352 49018 669361
rect 48962 669287 49018 669296
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47398 638208 47454 638217
rect 47398 638143 47454 638152
rect 47412 618905 47440 638143
rect 47398 618896 47454 618905
rect 47398 618831 47454 618840
rect 47216 611108 47268 611114
rect 47216 611050 47268 611056
rect 45374 598088 45430 598097
rect 45374 598023 45430 598032
rect 47596 582457 47624 662390
rect 50356 626657 50384 714818
rect 51736 691393 51764 753510
rect 62776 743073 62804 780399
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62960 741713 62988 793591
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 651470 776656 651526 776665
rect 651470 776591 651526 776600
rect 651484 775606 651512 776591
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62946 741704 63002 741713
rect 62946 741639 63002 741648
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 51724 674892 51776 674898
rect 51724 674834 51776 674840
rect 51736 646649 51764 674834
rect 51722 646640 51778 646649
rect 51722 646575 51778 646584
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 54484 647896 54536 647902
rect 54484 647838 54536 647844
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 50342 626648 50398 626657
rect 50342 626583 50398 626592
rect 48964 623824 49016 623830
rect 48964 623766 49016 623772
rect 48976 601361 49004 623766
rect 51736 601769 51764 636210
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 48962 601352 49018 601361
rect 48962 601287 49018 601296
rect 54496 600953 54524 647838
rect 55876 643249 55904 701014
rect 62776 697921 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 652036 718321 652064 842959
rect 652574 736808 652630 736817
rect 652574 736743 652630 736752
rect 652588 735622 652616 736743
rect 652576 735616 652628 735622
rect 652576 735558 652628 735564
rect 652022 718312 652078 718321
rect 652022 718247 652078 718256
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 652574 710288 652630 710297
rect 652574 710223 652630 710232
rect 652588 709374 652616 710223
rect 652576 709368 652628 709374
rect 652576 709310 652628 709316
rect 62762 697912 62818 697921
rect 62762 697847 62818 697856
rect 652392 696992 652444 696998
rect 652390 696960 652392 696969
rect 652444 696960 652446 696969
rect 652390 696895 652446 696904
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 652022 683632 652078 683641
rect 652022 683567 652078 683576
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 651470 670440 651526 670449
rect 651470 670375 651526 670384
rect 651484 669390 651512 670375
rect 651472 669384 651524 669390
rect 651472 669326 651524 669332
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 651470 657112 651526 657121
rect 651470 657047 651526 657056
rect 651484 656946 651512 657047
rect 651472 656940 651524 656946
rect 651472 656882 651524 656888
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 651470 630592 651526 630601
rect 651470 630527 651526 630536
rect 651484 629338 651512 630527
rect 651472 629332 651524 629338
rect 651472 629274 651524 629280
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 54482 600944 54538 600953
rect 54482 600879 54538 600888
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 582448 47638 582457
rect 47582 582383 47638 582392
rect 48976 557841 49004 597518
rect 51724 583772 51776 583778
rect 51724 583714 51776 583720
rect 48962 557832 49018 557841
rect 48962 557767 49018 557776
rect 51736 557569 51764 583714
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 51722 557560 51778 557569
rect 51722 557495 51778 557504
rect 45558 556880 45614 556889
rect 45558 556815 45614 556824
rect 45098 555656 45154 555665
rect 45098 555591 45154 555600
rect 44822 555248 44878 555257
rect 44822 555183 44878 555192
rect 44638 428904 44694 428913
rect 44638 428839 44694 428848
rect 44836 428097 44864 555183
rect 45006 551576 45062 551585
rect 45006 551511 45062 551520
rect 45020 529689 45048 551511
rect 45374 550896 45430 550905
rect 45374 550831 45430 550840
rect 45190 548720 45246 548729
rect 45190 548655 45246 548664
rect 45204 537033 45232 548655
rect 45190 537024 45246 537033
rect 45190 536959 45246 536968
rect 45388 532817 45416 550831
rect 45374 532808 45430 532817
rect 45374 532743 45430 532752
rect 45006 529680 45062 529689
rect 45006 529615 45062 529624
rect 45572 429729 45600 556815
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 45558 429720 45614 429729
rect 45558 429655 45614 429664
rect 45006 429312 45062 429321
rect 45006 429247 45062 429256
rect 44822 428088 44878 428097
rect 44822 428023 44878 428032
rect 44362 427272 44418 427281
rect 44362 427207 44418 427216
rect 44454 426864 44510 426873
rect 44454 426799 44510 426808
rect 44178 385656 44234 385665
rect 44178 385591 44234 385600
rect 44468 384033 44496 426799
rect 44638 421560 44694 421569
rect 44638 421495 44694 421504
rect 44652 407017 44680 421495
rect 44822 420744 44878 420753
rect 44822 420679 44878 420688
rect 44638 407008 44694 407017
rect 44638 406943 44694 406952
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44454 384024 44510 384033
rect 44454 383959 44510 383968
rect 44652 379514 44680 385183
rect 44836 379514 44864 420679
rect 45020 386753 45048 429247
rect 45190 427680 45246 427689
rect 45190 427615 45246 427624
rect 45006 386744 45062 386753
rect 45006 386679 45062 386688
rect 45204 384849 45232 427615
rect 45374 422376 45430 422385
rect 45374 422311 45430 422320
rect 45388 405657 45416 422311
rect 45374 405648 45430 405657
rect 45374 405583 45430 405592
rect 45374 386064 45430 386073
rect 45374 385999 45430 386008
rect 45190 384840 45246 384849
rect 45190 384775 45246 384784
rect 45006 384432 45062 384441
rect 45006 384367 45062 384376
rect 44652 379486 44772 379514
rect 44836 379486 44956 379514
rect 44454 377904 44510 377913
rect 44454 377839 44510 377848
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 44284 356697 44312 377431
rect 44468 364993 44496 377839
rect 44454 364984 44510 364993
rect 44454 364919 44510 364928
rect 44744 360194 44772 379486
rect 44744 360166 44864 360194
rect 44270 356688 44326 356697
rect 44270 356623 44326 356632
rect 44008 355830 44312 355858
rect 44284 355722 44312 355830
rect 43824 355694 44220 355722
rect 44284 355706 44680 355722
rect 44284 355700 44692 355706
rect 44284 355694 44640 355700
rect 44192 355586 44220 355694
rect 44640 355642 44692 355648
rect 43732 355558 43944 355586
rect 44192 355558 44772 355586
rect 43916 355450 43944 355558
rect 43916 355422 44128 355450
rect 43548 355286 44036 355314
rect 44008 354634 44036 355286
rect 44100 354906 44128 355422
rect 44100 354890 44615 354906
rect 44100 354884 44627 354890
rect 44100 354878 44575 354884
rect 44575 354826 44627 354832
rect 44575 354680 44627 354686
rect 44008 354628 44575 354634
rect 44008 354622 44627 354628
rect 44008 354606 44615 354622
rect 44744 354498 44772 355558
rect 44836 354634 44864 360166
rect 44928 357434 44956 379486
rect 45020 360194 45048 384367
rect 45190 383616 45246 383625
rect 45190 383551 45246 383560
rect 45204 379514 45232 383551
rect 45204 379486 45324 379514
rect 45020 360166 45232 360194
rect 44928 357406 45048 357434
rect 45020 355842 45048 357406
rect 45008 355836 45060 355842
rect 45008 355778 45060 355784
rect 44836 354606 44956 354634
rect 44744 354482 44839 354498
rect 44744 354476 44851 354482
rect 44744 354470 44799 354476
rect 44799 354418 44851 354424
rect 44686 354340 44738 354346
rect 44686 354282 44738 354288
rect 43902 354240 43958 354249
rect 44698 354226 44726 354282
rect 43958 354198 44726 354226
rect 43902 354175 43958 354184
rect 44730 353832 44786 353841
rect 44928 353818 44956 354606
rect 45204 354090 45232 360166
rect 44786 353790 44956 353818
rect 45020 354062 45232 354090
rect 44730 353767 44786 353776
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 38290 346352 38346 346361
rect 38290 346287 38346 346296
rect 38304 345098 38332 346287
rect 28908 345092 28960 345098
rect 28908 345034 28960 345040
rect 38292 345092 38344 345098
rect 38292 345034 38344 345040
rect 28920 344321 28948 345034
rect 28906 344312 28962 344321
rect 28906 344247 28962 344256
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 45020 341737 45048 354062
rect 45296 345014 45324 379486
rect 45204 344986 45324 345014
rect 45006 341728 45062 341737
rect 45006 341663 45062 341672
rect 45204 340921 45232 344986
rect 45388 343369 45416 385999
rect 45558 383208 45614 383217
rect 45558 383143 45614 383152
rect 45572 356969 45600 383143
rect 45742 379128 45798 379137
rect 45742 379063 45798 379072
rect 45756 364313 45784 379063
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 426456 46994 426465
rect 46938 426391 46994 426400
rect 46952 399809 46980 426391
rect 47122 423600 47178 423609
rect 47122 423535 47178 423544
rect 47136 400217 47164 423535
rect 47122 400208 47178 400217
rect 47122 400143 47178 400152
rect 46938 399800 46994 399809
rect 46938 399735 46994 399744
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 46938 380760 46994 380769
rect 46938 380695 46994 380704
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 45742 364304 45798 364313
rect 45742 364239 45798 364248
rect 46388 362976 46440 362982
rect 46388 362918 46440 362924
rect 45558 356960 45614 356969
rect 45558 356895 45614 356904
rect 45650 356688 45706 356697
rect 45480 356646 45650 356674
rect 45480 353274 45508 356646
rect 45650 356623 45706 356632
rect 45926 355872 45982 355881
rect 45652 355836 45704 355842
rect 45926 355807 45982 355816
rect 45652 355778 45704 355784
rect 45664 354074 45692 355778
rect 45652 354068 45704 354074
rect 45652 354010 45704 354016
rect 45940 353802 45968 355807
rect 45928 353796 45980 353802
rect 45928 353738 45980 353744
rect 45480 353258 45600 353274
rect 45480 353252 45612 353258
rect 45480 353246 45560 353252
rect 45560 353194 45612 353200
rect 45374 343360 45430 343369
rect 45374 343295 45430 343304
rect 45190 340912 45246 340921
rect 45190 340847 45246 340856
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37924 339516 37976 339522
rect 37924 339458 37976 339464
rect 35806 339008 35862 339017
rect 35806 338943 35862 338952
rect 31022 338600 31078 338609
rect 31022 338535 31078 338544
rect 31036 329089 31064 338535
rect 35820 338162 35848 338943
rect 35808 338156 35860 338162
rect 35808 338098 35860 338104
rect 36544 338156 36596 338162
rect 36544 338098 36596 338104
rect 31022 329080 31078 329089
rect 31022 329015 31078 329024
rect 36556 328409 36584 338098
rect 37936 335345 37964 339458
rect 45650 338464 45706 338473
rect 45650 338399 45706 338408
rect 45466 337240 45522 337249
rect 45466 337175 45522 337184
rect 37922 335336 37978 335345
rect 37922 335271 37978 335280
rect 42798 334656 42854 334665
rect 42798 334591 42854 334600
rect 43166 334656 43222 334665
rect 43166 334591 43222 334600
rect 44270 334656 44326 334665
rect 44270 334591 44326 334600
rect 36542 328400 36598 328409
rect 36542 328335 36598 328344
rect 41786 326768 41842 326777
rect 41786 326703 41842 326712
rect 41800 326264 41828 326703
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41786 324728 41842 324737
rect 41786 324663 41842 324672
rect 41800 324428 41828 324663
rect 42182 323734 42472 323762
rect 42246 323640 42302 323649
rect 42246 323575 42302 323584
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42260 321382 42288 323575
rect 42444 321473 42472 323734
rect 42430 321464 42486 321473
rect 42430 321399 42486 321408
rect 42182 321354 42288 321382
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 41800 320725 41828 321127
rect 42430 320104 42486 320113
rect 42182 320062 42430 320090
rect 42430 320039 42486 320048
rect 42182 319518 42472 319546
rect 42444 318889 42472 319518
rect 42430 318880 42486 318889
rect 42430 318815 42486 318824
rect 42812 318794 42840 334591
rect 42982 334384 43038 334393
rect 42982 334319 43038 334328
rect 42996 323649 43024 334319
rect 42982 323640 43038 323649
rect 42982 323575 43038 323584
rect 43180 322833 43208 334591
rect 43442 322960 43498 322969
rect 43442 322895 43498 322904
rect 43166 322824 43222 322833
rect 43166 322759 43222 322768
rect 42812 318766 43024 318794
rect 42996 317098 43024 318766
rect 42536 317070 43024 317098
rect 42536 317059 42564 317070
rect 42182 317031 42564 317059
rect 42430 316432 42486 316441
rect 42182 316390 42430 316418
rect 42430 316367 42486 316376
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 41878 315616 41934 315625
rect 41878 315551 41934 315560
rect 41892 315180 41920 315551
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42062 312624 42118 312633
rect 42062 312559 42118 312568
rect 42076 312052 42104 312559
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 42890 299704 42946 299713
rect 42890 299639 42946 299648
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 41326 296032 41382 296041
rect 41326 295967 41382 295976
rect 32402 294808 32458 294817
rect 32402 294743 32458 294752
rect 32416 284986 32444 294743
rect 41340 291394 41368 295967
rect 41800 292505 41828 296783
rect 41786 292496 41842 292505
rect 41786 292431 41842 292440
rect 41340 291366 41460 291394
rect 41432 290442 41460 291366
rect 41786 290456 41842 290465
rect 41432 290414 41786 290442
rect 41786 290391 41842 290400
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 285122 41368 290255
rect 41328 285116 41380 285122
rect 41328 285058 41380 285064
rect 41696 285116 41748 285122
rect 41748 285076 42380 285104
rect 41696 285058 41748 285064
rect 32404 284980 32456 284986
rect 32404 284922 32456 284928
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42288 284866
rect 42260 283059 42288 284838
rect 42182 283031 42288 283059
rect 42352 281874 42380 285076
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42430 278695 42486 278704
rect 42338 278488 42394 278497
rect 42338 278423 42394 278432
rect 42168 277953 42196 278188
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 42154 277944 42210 277953
rect 42154 277879 42210 277888
rect 41800 277508 41828 277879
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42062 273456 42118 273465
rect 42062 273391 42118 273400
rect 42076 273224 42104 273391
rect 42062 273048 42118 273057
rect 42062 272983 42118 272992
rect 42076 272544 42104 272983
rect 42352 272014 42380 278423
rect 42182 271986 42380 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 42430 270464 42486 270473
rect 42430 270399 42486 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 270399
rect 42182 269507 42472 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 42904 256873 42932 299639
rect 43258 298888 43314 298897
rect 43258 298823 43314 298832
rect 43074 295216 43130 295225
rect 43074 295151 43130 295160
rect 43088 276593 43116 295151
rect 43074 276584 43130 276593
rect 43074 276519 43130 276528
rect 42890 256864 42946 256873
rect 42890 256799 42946 256808
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 43272 256057 43300 298823
rect 43456 257689 43484 322895
rect 44284 320113 44312 334591
rect 44270 320104 44326 320113
rect 44270 320039 44326 320048
rect 45480 316033 45508 337175
rect 45664 318889 45692 338399
rect 45650 318880 45706 318889
rect 45650 318815 45706 318824
rect 45466 316024 45522 316033
rect 45466 315959 45522 315968
rect 44730 311536 44786 311545
rect 44730 311471 44786 311480
rect 44362 311264 44418 311273
rect 44362 311199 44418 311208
rect 44376 298489 44404 311199
rect 44546 311128 44602 311137
rect 44546 311063 44602 311072
rect 44560 299305 44588 311063
rect 44744 300121 44772 311471
rect 46400 303113 46428 362918
rect 46952 356153 46980 380695
rect 47122 379944 47178 379953
rect 47122 379879 47178 379888
rect 47136 357377 47164 379879
rect 47122 357368 47178 357377
rect 47122 357303 47178 357312
rect 46938 356144 46994 356153
rect 46938 356079 46994 356088
rect 46938 340096 46994 340105
rect 46938 340031 46994 340040
rect 46952 313721 46980 340031
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46938 313712 46994 313721
rect 46938 313647 46994 313656
rect 46386 303104 46442 303113
rect 46386 303039 46442 303048
rect 44730 300112 44786 300121
rect 44730 300047 44786 300056
rect 44546 299296 44602 299305
rect 44546 299231 44602 299240
rect 44362 298480 44418 298489
rect 44362 298415 44418 298424
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 44178 298072 44234 298081
rect 44178 298007 44234 298016
rect 43626 293992 43682 294001
rect 43626 293927 43682 293936
rect 43640 273057 43668 293927
rect 43810 293176 43866 293185
rect 43810 293111 43866 293120
rect 43824 279857 43852 293111
rect 43994 291952 44050 291961
rect 43994 291887 44050 291896
rect 43810 279848 43866 279857
rect 43810 279783 43866 279792
rect 44008 277137 44036 291887
rect 43994 277128 44050 277137
rect 43994 277063 44050 277072
rect 43626 273048 43682 273057
rect 43626 272983 43682 272992
rect 43442 257680 43498 257689
rect 43442 257615 43498 257624
rect 43626 256456 43682 256465
rect 43626 256391 43682 256400
rect 43258 256048 43314 256057
rect 43258 255983 43314 255992
rect 42982 255640 43038 255649
rect 42982 255575 43038 255584
rect 42798 254824 42854 254833
rect 42798 254759 42854 254768
rect 35438 253464 35494 253473
rect 35438 253399 35494 253408
rect 35452 252618 35480 253399
rect 35622 253056 35678 253065
rect 35622 252991 35678 253000
rect 35636 252754 35664 252991
rect 35808 252884 35860 252890
rect 35808 252826 35860 252832
rect 40684 252884 40736 252890
rect 40684 252826 40736 252832
rect 35624 252748 35676 252754
rect 35624 252690 35676 252696
rect 35820 252657 35848 252826
rect 35806 252648 35862 252657
rect 35440 252612 35492 252618
rect 35806 252583 35862 252592
rect 35440 252554 35492 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 36544 251252 36596 251258
rect 36544 251194 36596 251200
rect 36556 242894 36584 251194
rect 36544 242888 36596 242894
rect 36544 242830 36596 242836
rect 40696 242593 40724 252826
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 41328 252612 41380 252618
rect 41328 252554 41380 252560
rect 41340 252249 41368 252554
rect 41326 252240 41382 252249
rect 41326 252175 41382 252184
rect 41708 248414 41736 252690
rect 42614 252240 42670 252249
rect 42614 252175 42670 252184
rect 42628 248414 42656 252175
rect 41708 248386 42012 248414
rect 41984 244274 42012 248386
rect 42536 248386 42656 248414
rect 41984 244246 42196 244274
rect 41696 242888 41748 242894
rect 41694 242856 41696 242865
rect 41748 242856 41750 242865
rect 41694 242791 41750 242800
rect 42168 242706 42196 244246
rect 42338 242856 42394 242865
rect 42338 242791 42394 242800
rect 42168 242678 42288 242706
rect 40682 242584 40738 242593
rect 40682 242519 40738 242528
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42076 238513 42104 238649
rect 42062 238504 42118 238513
rect 42062 238439 42118 238448
rect 42260 238014 42288 242678
rect 42182 237986 42288 238014
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42154 235376 42210 235385
rect 42154 235311 42210 235320
rect 42168 234969 42196 235311
rect 42352 234614 42380 242791
rect 42536 238105 42564 248386
rect 42522 238096 42578 238105
rect 42522 238031 42578 238040
rect 42352 234586 42748 234614
rect 42182 234314 42472 234342
rect 42246 234152 42302 234161
rect 42246 234087 42302 234096
rect 42260 233695 42288 234087
rect 42444 233889 42472 234314
rect 42430 233880 42486 233889
rect 42430 233815 42486 233824
rect 42182 233667 42288 233695
rect 42338 233200 42394 233209
rect 42168 233158 42338 233186
rect 42168 233104 42196 233158
rect 42338 233135 42394 233144
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 42154 230208 42210 230217
rect 42154 230143 42210 230152
rect 42168 229976 42196 230143
rect 42430 229392 42486 229401
rect 42182 229350 42430 229378
rect 42430 229327 42486 229336
rect 42720 229094 42748 234586
rect 42536 229066 42748 229094
rect 42536 228834 42564 229066
rect 42182 228806 42564 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 40682 222864 40738 222873
rect 40682 222799 40738 222808
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214305 35572 217903
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 40696 213994 40724 222799
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 40684 213988 40736 213994
rect 40684 213930 40736 213936
rect 42812 212129 42840 254759
rect 42996 212945 43024 255575
rect 43442 251152 43498 251161
rect 43442 251087 43498 251096
rect 43258 242584 43314 242593
rect 43258 242519 43314 242528
rect 43272 229094 43300 242519
rect 43456 229094 43484 251087
rect 43640 251002 43668 256391
rect 44192 255241 44220 298007
rect 44638 297256 44694 297265
rect 44638 297191 44694 297200
rect 44362 294400 44418 294409
rect 44362 294335 44418 294344
rect 44376 270473 44404 294335
rect 44362 270464 44418 270473
rect 44362 270399 44418 270408
rect 44178 255232 44234 255241
rect 44178 255167 44234 255176
rect 44652 254425 44680 297191
rect 45480 296714 45508 298114
rect 44836 296686 45508 296714
rect 44638 254416 44694 254425
rect 44638 254351 44694 254360
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43180 229066 43300 229094
rect 43364 229066 43484 229094
rect 43548 250974 43668 251002
rect 43180 225729 43208 229066
rect 43364 226681 43392 229066
rect 43350 226672 43406 226681
rect 43350 226607 43406 226616
rect 43166 225720 43222 225729
rect 43166 225655 43222 225664
rect 43548 213761 43576 250974
rect 43718 249112 43774 249121
rect 43718 249047 43774 249056
rect 43732 231849 43760 249047
rect 43718 231840 43774 231849
rect 43718 231775 43774 231784
rect 43534 213752 43590 213761
rect 43534 213687 43590 213696
rect 42982 212936 43038 212945
rect 42982 212871 43038 212880
rect 42798 212120 42854 212129
rect 42798 212055 42854 212064
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35820 211206 35848 211375
rect 44192 211313 44220 253943
rect 44546 251968 44602 251977
rect 44546 251903 44602 251912
rect 44362 248704 44418 248713
rect 44362 248639 44418 248648
rect 44376 234161 44404 248639
rect 44362 234152 44418 234161
rect 44362 234087 44418 234096
rect 44560 233209 44588 251903
rect 44546 233200 44602 233209
rect 44546 233135 44602 233144
rect 44836 214985 44864 296686
rect 45006 293584 45062 293593
rect 45006 293519 45062 293528
rect 45020 273465 45048 293519
rect 45190 291680 45246 291689
rect 45190 291615 45246 291624
rect 45204 277953 45232 291615
rect 46202 290728 46258 290737
rect 46202 290663 46258 290672
rect 45190 277944 45246 277953
rect 45190 277879 45246 277888
rect 45006 273456 45062 273465
rect 45006 273391 45062 273400
rect 45558 250744 45614 250753
rect 45558 250679 45614 250688
rect 45006 248296 45062 248305
rect 45006 248231 45062 248240
rect 45020 235385 45048 248231
rect 45006 235376 45062 235385
rect 45006 235311 45062 235320
rect 45572 229401 45600 250679
rect 45834 250336 45890 250345
rect 45834 250271 45890 250280
rect 45848 230217 45876 250271
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 233889 46060 249455
rect 46018 233880 46074 233889
rect 46018 233815 46074 233824
rect 45834 230208 45890 230217
rect 45834 230143 45890 230152
rect 45558 229392 45614 229401
rect 45558 229327 45614 229336
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 45006 213344 45062 213353
rect 45006 213279 45062 213288
rect 44178 211304 44234 211313
rect 44178 211239 44234 211248
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 41696 211200 41748 211206
rect 41696 211142 41748 211148
rect 41708 209001 41736 211142
rect 43258 210896 43314 210905
rect 43258 210831 43314 210840
rect 42798 209400 42854 209409
rect 42798 209335 42854 209344
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 41694 208992 41750 209001
rect 41694 208927 41750 208936
rect 35820 208418 35848 208927
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 207777 40080 208354
rect 40038 207768 40094 207777
rect 40038 207703 40094 207712
rect 35622 204096 35678 204105
rect 35622 204031 35678 204040
rect 35636 202201 35664 204031
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 35622 202192 35678 202201
rect 35622 202127 35678 202136
rect 37936 197849 37964 202846
rect 37922 197840 37978 197849
rect 37922 197775 37978 197784
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 41878 195800 41934 195809
rect 41878 195735 41934 195744
rect 41892 195432 41920 195735
rect 42614 195528 42670 195537
rect 42614 195463 42670 195472
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42628 192953 42656 195463
rect 42168 192902 42288 192930
rect 42614 192944 42670 192953
rect 42614 192879 42670 192888
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41786 187232 41842 187241
rect 41786 187167 41842 187176
rect 41800 186796 41828 187167
rect 42168 186130 42196 186184
rect 42338 186144 42394 186153
rect 42168 186102 42338 186130
rect 42338 186079 42394 186088
rect 41970 185872 42026 185881
rect 41970 185807 42026 185816
rect 41984 185605 42012 185807
rect 42430 184920 42486 184929
rect 42430 184855 42486 184864
rect 42444 183779 42472 184855
rect 42182 183751 42472 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42812 182491 42840 209335
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 43272 206281 43300 210831
rect 44178 210488 44234 210497
rect 44178 210423 44234 210432
rect 43442 208040 43498 208049
rect 43442 207975 43498 207984
rect 43258 206272 43314 206281
rect 43258 206207 43314 206216
rect 43456 206122 43484 207975
rect 43994 206816 44050 206825
rect 43994 206751 44050 206760
rect 43272 206094 43484 206122
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 183161 43300 206094
rect 43810 205592 43866 205601
rect 43810 205527 43866 205536
rect 43626 205184 43682 205193
rect 43626 205119 43682 205128
rect 43442 202192 43498 202201
rect 43442 202127 43498 202136
rect 43258 183152 43314 183161
rect 43258 183087 43314 183096
rect 42182 182463 42840 182491
rect 43456 42838 43484 202127
rect 43640 191729 43668 205119
rect 43626 191720 43682 191729
rect 43626 191655 43682 191664
rect 43824 190505 43852 205527
rect 44008 193225 44036 206751
rect 43994 193216 44050 193225
rect 43994 193151 44050 193160
rect 43810 190496 43866 190505
rect 43810 190431 43866 190440
rect 44192 184929 44220 210423
rect 45020 209774 45048 213279
rect 45020 209746 45508 209774
rect 44362 208584 44418 208593
rect 44362 208519 44418 208528
rect 44376 189961 44404 208519
rect 44546 206000 44602 206009
rect 44546 205935 44602 205944
rect 44362 189952 44418 189961
rect 44362 189887 44418 189896
rect 44560 187649 44588 205935
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44546 187640 44602 187649
rect 44546 187575 44602 187584
rect 44178 184920 44234 184929
rect 44178 184855 44234 184864
rect 44836 74534 44864 204711
rect 45480 196654 45508 209746
rect 45468 196648 45520 196654
rect 45468 196590 45520 196596
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 290663
rect 46938 247072 46994 247081
rect 46938 247007 46994 247016
rect 46952 238513 46980 247007
rect 46938 238504 46994 238513
rect 46938 238439 46994 238448
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 47596 49026 47624 333095
rect 47780 300529 47808 389234
rect 48976 387025 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 49148 415472 49200 415478
rect 49148 415414 49200 415420
rect 48962 387016 49018 387025
rect 48962 386951 49018 386960
rect 49160 346361 49188 415414
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51724 375420 51776 375426
rect 51724 375362 51776 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 49146 346352 49202 346361
rect 49146 346287 49202 346296
rect 50344 336796 50396 336802
rect 50344 336738 50396 336744
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47780 53242 47808 247415
rect 47950 212528 48006 212537
rect 47950 212463 48006 212472
rect 47964 192409 47992 212463
rect 48780 196648 48832 196654
rect 48780 196590 48832 196596
rect 47950 192400 48006 192409
rect 47950 192335 48006 192344
rect 48792 190505 48820 196590
rect 48778 190496 48834 190505
rect 48778 190431 48834 190440
rect 47768 53236 47820 53242
rect 47768 53178 47820 53184
rect 48976 51746 49004 334047
rect 49146 289912 49202 289921
rect 49146 289847 49202 289856
rect 49160 51882 49188 289847
rect 50356 257825 50384 336738
rect 51736 301345 51764 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 651470 590744 651526 590753
rect 651470 590679 651472 590688
rect 651524 590679 651526 590688
rect 651472 590650 651524 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 652036 583001 652064 683567
rect 660316 625297 660344 763166
rect 661696 760481 661724 921810
rect 663064 909492 663116 909498
rect 663064 909434 663116 909440
rect 663076 760889 663104 909434
rect 671344 895688 671396 895694
rect 671344 895630 671396 895636
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868737 664484 881826
rect 669226 879200 669282 879209
rect 669226 879135 669282 879144
rect 664442 868728 664498 868737
rect 664442 868663 664498 868672
rect 668214 868184 668270 868193
rect 668214 868119 668270 868128
rect 664444 855636 664496 855642
rect 664444 855578 664496 855584
rect 663062 760880 663118 760889
rect 663062 760815 663118 760824
rect 661682 760472 661738 760481
rect 661682 760407 661738 760416
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 661684 696992 661736 696998
rect 661684 696934 661736 696940
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 660316 599593 660344 616830
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 652022 582992 652078 583001
rect 652022 582927 652078 582936
rect 661696 581097 661724 696934
rect 663076 689353 663104 723114
rect 664456 716553 664484 855578
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666282 777064 666338 777073
rect 666282 776999 666338 777008
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 661868 669384 661920 669390
rect 661868 669326 661920 669332
rect 661880 643793 661908 669326
rect 661866 643784 661922 643793
rect 661866 643719 661922 643728
rect 662052 590708 662104 590714
rect 662052 590650 662104 590656
rect 661682 581088 661738 581097
rect 661682 581023 661738 581032
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 658936 554033 658964 563042
rect 658922 554024 658978 554033
rect 658922 553959 658978 553968
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 652574 497720 652630 497729
rect 652574 497655 652630 497664
rect 652588 494766 652616 497655
rect 652576 494760 652628 494766
rect 652576 494702 652628 494708
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 54484 310548 54536 310554
rect 54484 310490 54536 310496
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 51722 289912 51778 289921
rect 51722 289847 51778 289856
rect 50342 257816 50398 257825
rect 50342 257751 50398 257760
rect 50526 247752 50582 247761
rect 50526 247687 50582 247696
rect 50342 246528 50398 246537
rect 50342 246463 50398 246472
rect 49330 208992 49386 209001
rect 49330 208927 49386 208936
rect 49344 196489 49372 208927
rect 49514 206272 49570 206281
rect 49514 206207 49570 206216
rect 49330 196480 49386 196489
rect 49330 196415 49386 196424
rect 49528 194449 49556 206207
rect 49514 194440 49570 194449
rect 49514 194375 49570 194384
rect 49148 51876 49200 51882
rect 49148 51818 49200 51824
rect 48964 51740 49016 51746
rect 48964 51682 49016 51688
rect 50356 50522 50384 246463
rect 50540 53378 50568 247687
rect 50710 203280 50766 203289
rect 50710 203215 50766 203224
rect 50528 53372 50580 53378
rect 50528 53314 50580 53320
rect 50724 52018 50752 203215
rect 50712 52012 50764 52018
rect 50712 51954 50764 51960
rect 50344 50516 50396 50522
rect 50344 50458 50396 50464
rect 51736 49162 51764 289847
rect 54496 217977 54524 310490
rect 55876 278769 55904 401610
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 652022 378176 652078 378185
rect 652022 378111 652078 378120
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 651654 364848 651710 364857
rect 651654 364783 651710 364792
rect 651668 364410 651696 364783
rect 651656 364404 651708 364410
rect 651656 364346 651708 364352
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 651470 351656 651526 351665
rect 651470 351591 651526 351600
rect 651484 350606 651512 351591
rect 651472 350600 651524 350606
rect 651472 350542 651524 350548
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 62776 267073 62804 350231
rect 651470 338328 651526 338337
rect 651470 338263 651526 338272
rect 651484 338162 651512 338263
rect 651472 338156 651524 338162
rect 651472 338098 651524 338104
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 651484 310554 651512 311743
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62946 285152 63002 285161
rect 62946 285087 63002 285096
rect 62762 267064 62818 267073
rect 62762 266999 62818 267008
rect 62764 228540 62816 228546
rect 62764 228482 62816 228488
rect 57888 227044 57940 227050
rect 57888 226986 57940 226992
rect 56508 222352 56560 222358
rect 56508 222294 56560 222300
rect 56324 218204 56376 218210
rect 56324 218146 56376 218152
rect 55680 218068 55732 218074
rect 55680 218010 55732 218016
rect 54482 217968 54538 217977
rect 54482 217903 54538 217912
rect 55692 217138 55720 218010
rect 56336 217274 56364 218146
rect 56520 218074 56548 222294
rect 57900 218074 57928 226986
rect 61292 225616 61344 225622
rect 61292 225558 61344 225564
rect 60648 224528 60700 224534
rect 60648 224470 60700 224476
rect 58992 224256 59044 224262
rect 58992 224198 59044 224204
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57336 218068 57388 218074
rect 57336 218010 57388 218016
rect 57888 218068 57940 218074
rect 57888 218010 57940 218016
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 56336 217246 56502 217274
rect 55646 217110 55720 217138
rect 55646 216988 55674 217110
rect 56474 216988 56502 217246
rect 57348 217138 57376 218010
rect 58176 217138 58204 218010
rect 59004 217274 59032 224198
rect 59820 218612 59872 218618
rect 59820 218554 59872 218560
rect 57302 217110 57376 217138
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 57302 216988 57330 217110
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218554
rect 60660 217274 60688 224470
rect 61304 218074 61332 225558
rect 61476 221604 61528 221610
rect 61476 221546 61528 221552
rect 61292 218068 61344 218074
rect 61292 218010 61344 218016
rect 61488 217274 61516 221546
rect 62304 218884 62356 218890
rect 62304 218826 62356 218832
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 61442 217246 61516 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61442 216988 61470 217246
rect 62316 217138 62344 218826
rect 62776 218210 62804 228482
rect 62960 222873 62988 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 274666 65932 277780
rect 67008 274718 67036 277780
rect 66996 274712 67048 274718
rect 65904 274638 66300 274666
rect 66996 274654 67048 274660
rect 66272 268394 66300 274638
rect 68204 271182 68232 277780
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274990 71820 277780
rect 71780 274984 71832 274990
rect 71780 274926 71832 274932
rect 71044 274712 71096 274718
rect 71044 274654 71096 274660
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 66260 268388 66312 268394
rect 66260 268330 66312 268336
rect 71056 267170 71084 274654
rect 72988 271318 73016 277780
rect 74092 275194 74120 277780
rect 75302 277766 75868 277794
rect 74080 275188 74132 275194
rect 74080 275130 74132 275136
rect 73804 274984 73856 274990
rect 73804 274926 73856 274932
rect 72976 271312 73028 271318
rect 72976 271254 73028 271260
rect 71044 267164 71096 267170
rect 71044 267106 71096 267112
rect 73816 267034 73844 274926
rect 75840 269958 75868 277766
rect 76484 275602 76512 277780
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 77208 275188 77260 275194
rect 77208 275130 77260 275136
rect 77220 273970 77248 275130
rect 77208 273964 77260 273970
rect 77208 273906 77260 273912
rect 77680 272542 77708 277780
rect 78876 272950 78904 277780
rect 78864 272944 78916 272950
rect 78864 272886 78916 272892
rect 77668 272536 77720 272542
rect 77668 272478 77720 272484
rect 80072 270094 80100 277780
rect 81268 275738 81296 277780
rect 81256 275732 81308 275738
rect 81256 275674 81308 275680
rect 82372 274106 82400 277780
rect 83582 277766 84148 277794
rect 82360 274100 82412 274106
rect 82360 274042 82412 274048
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 84120 269686 84148 277766
rect 84764 274242 84792 277780
rect 85960 275466 85988 277780
rect 86868 275596 86920 275602
rect 86868 275538 86920 275544
rect 85948 275460 86000 275466
rect 85948 275402 86000 275408
rect 84752 274236 84804 274242
rect 84752 274178 84804 274184
rect 84108 269680 84160 269686
rect 84108 269622 84160 269628
rect 86880 268938 86908 275538
rect 87156 272678 87184 277780
rect 88352 276010 88380 277780
rect 89548 277394 89576 277780
rect 89548 277366 89668 277394
rect 88340 276004 88392 276010
rect 88340 275946 88392 275952
rect 89640 275890 89668 277366
rect 89640 275862 89760 275890
rect 88984 275732 89036 275738
rect 88984 275674 89036 275680
rect 87144 272672 87196 272678
rect 87144 272614 87196 272620
rect 86868 268932 86920 268938
rect 86868 268874 86920 268880
rect 88996 267578 89024 275674
rect 89732 271454 89760 275862
rect 90652 274718 90680 277780
rect 91862 277766 92428 277794
rect 90640 274712 90692 274718
rect 90640 274654 90692 274660
rect 89720 271448 89772 271454
rect 89720 271390 89772 271396
rect 92400 268530 92428 277766
rect 93044 271726 93072 277780
rect 94240 272814 94268 277780
rect 95436 275874 95464 277780
rect 95424 275868 95476 275874
rect 95424 275810 95476 275816
rect 96632 275602 96660 277780
rect 97750 277766 97948 277794
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 96620 275596 96672 275602
rect 96620 275538 96672 275544
rect 95884 274712 95936 274718
rect 95884 274654 95936 274660
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 93032 271720 93084 271726
rect 93032 271662 93084 271668
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 95896 267714 95924 274654
rect 97920 270230 97948 277766
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 99300 268666 99328 277766
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 95884 267708 95936 267714
rect 95884 267650 95936 267656
rect 88984 267572 89036 267578
rect 88984 267514 89036 267520
rect 100680 267306 100708 277766
rect 101324 274378 101352 277780
rect 101312 274372 101364 274378
rect 101312 274314 101364 274320
rect 102520 268802 102548 277780
rect 103716 275738 103744 277780
rect 104912 277394 104940 277780
rect 104912 277366 105032 277394
rect 104808 275868 104860 275874
rect 104808 275810 104860 275816
rect 103704 275732 103756 275738
rect 103704 275674 103756 275680
rect 104820 274650 104848 275810
rect 104808 274644 104860 274650
rect 104808 274586 104860 274592
rect 105004 273086 105032 277366
rect 106016 274786 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 274780 106056 274786
rect 106004 274722 106056 274728
rect 104992 273080 105044 273086
rect 104992 273022 105044 273028
rect 102508 268796 102560 268802
rect 102508 268738 102560 268744
rect 107580 267442 107608 277766
rect 108960 269074 108988 277766
rect 110248 270366 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 110420 274780 110472 274786
rect 110420 274722 110472 274728
rect 110432 271862 110460 274722
rect 110420 271856 110472 271862
rect 110420 271798 110472 271804
rect 111996 271590 112024 277780
rect 113192 275874 113220 277780
rect 113180 275868 113232 275874
rect 113180 275810 113232 275816
rect 114296 273222 114324 277780
rect 115506 277766 115888 277794
rect 114284 273216 114336 273222
rect 114284 273158 114336 273164
rect 111984 271584 112036 271590
rect 111984 271526 112036 271532
rect 115860 270502 115888 277766
rect 116688 270638 116716 277780
rect 117898 277766 118648 277794
rect 116676 270632 116728 270638
rect 116676 270574 116728 270580
rect 115848 270496 115900 270502
rect 115848 270438 115900 270444
rect 110236 270360 110288 270366
rect 110236 270302 110288 270308
rect 118620 269414 118648 277766
rect 119080 269550 119108 277780
rect 120290 277766 120948 277794
rect 120920 271726 120948 277766
rect 121380 274514 121408 277780
rect 122590 277766 122788 277794
rect 121368 274508 121420 274514
rect 121368 274450 121420 274456
rect 120724 271720 120776 271726
rect 120724 271662 120776 271668
rect 120908 271720 120960 271726
rect 120908 271662 120960 271668
rect 119804 269680 119856 269686
rect 119804 269622 119856 269628
rect 119068 269544 119120 269550
rect 119068 269486 119120 269492
rect 118608 269408 118660 269414
rect 118608 269350 118660 269356
rect 108948 269068 109000 269074
rect 108948 269010 109000 269016
rect 107568 267436 107620 267442
rect 107568 267378 107620 267384
rect 100668 267300 100720 267306
rect 100668 267242 100720 267248
rect 73804 267028 73856 267034
rect 73804 266970 73856 266976
rect 119816 266490 119844 269622
rect 120736 266762 120764 271662
rect 122760 268258 122788 277766
rect 123772 273834 123800 277780
rect 124982 277766 125548 277794
rect 126178 277766 126928 277794
rect 123760 273828 123812 273834
rect 123760 273770 123812 273776
rect 122748 268252 122800 268258
rect 122748 268194 122800 268200
rect 125520 267986 125548 277766
rect 126900 269550 126928 277766
rect 127360 272406 127388 277780
rect 127348 272400 127400 272406
rect 127348 272342 127400 272348
rect 128556 271046 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 128544 271040 128596 271046
rect 128544 270982 128596 270988
rect 130856 270910 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 270904 130896 270910
rect 130844 270846 130896 270852
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 125508 267980 125560 267986
rect 125508 267922 125560 267928
rect 132420 266898 132448 277766
rect 133800 268122 133828 277766
rect 134444 273698 134472 277780
rect 135640 275058 135668 277780
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136548 274916 136600 274922
rect 136548 274858 136600 274864
rect 134432 273692 134484 273698
rect 134432 273634 134484 273640
rect 136560 269793 136588 274858
rect 136546 269784 136602 269793
rect 136546 269719 136602 269728
rect 136836 269278 136864 277780
rect 137940 270774 137968 277780
rect 138664 272944 138716 272950
rect 138664 272886 138716 272892
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137928 270768 137980 270774
rect 137928 270710 137980 270716
rect 136824 269272 136876 269278
rect 136824 269214 136876 269220
rect 137284 268388 137336 268394
rect 137284 268330 137336 268336
rect 133788 268116 133840 268122
rect 133788 268058 133840 268064
rect 132408 266892 132460 266898
rect 132408 266834 132460 266840
rect 120724 266756 120776 266762
rect 120724 266698 120776 266704
rect 119804 266484 119856 266490
rect 119804 266426 119856 266432
rect 137296 264316 137324 268330
rect 138112 267164 138164 267170
rect 138112 267106 138164 267112
rect 138124 264316 138152 267106
rect 138492 264330 138520 271118
rect 138676 266626 138704 272886
rect 139136 272270 139164 277780
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 139124 272264 139176 272270
rect 139124 272206 139176 272212
rect 139768 269816 139820 269822
rect 139952 269816 140004 269822
rect 139768 269758 139820 269764
rect 139950 269784 139952 269793
rect 140004 269784 140006 269793
rect 138664 266620 138716 266626
rect 138664 266562 138716 266568
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 139950 269719 140006 269728
rect 140148 264330 140176 275266
rect 140332 274786 140360 277780
rect 141542 277766 141832 277794
rect 140320 274780 140372 274786
rect 140320 274722 140372 274728
rect 141804 272950 141832 277766
rect 142724 275330 142752 277780
rect 143356 276004 143408 276010
rect 143356 275946 143408 275952
rect 142712 275324 142764 275330
rect 142712 275266 142764 275272
rect 141792 272944 141844 272950
rect 141792 272886 141844 272892
rect 141424 272264 141476 272270
rect 141424 272206 141476 272212
rect 141436 267170 141464 272206
rect 142160 271312 142212 271318
rect 142160 271254 142212 271260
rect 141424 267164 141476 267170
rect 141424 267106 141476 267112
rect 141424 267028 141476 267034
rect 141424 266970 141476 266976
rect 140148 264302 140622 264330
rect 141436 264316 141464 266970
rect 142172 264330 142200 271254
rect 143368 269958 143396 275946
rect 143540 273964 143592 273970
rect 143540 273906 143592 273912
rect 142620 269952 142672 269958
rect 142620 269894 142672 269900
rect 143356 269952 143408 269958
rect 143356 269894 143408 269900
rect 142632 267734 142660 269894
rect 142632 267706 142752 267734
rect 142724 264330 142752 267706
rect 143552 264330 143580 273906
rect 143920 272270 143948 277780
rect 144644 274780 144696 274786
rect 144644 274722 144696 274728
rect 144656 273562 144684 274722
rect 145024 273970 145052 277780
rect 146220 274786 146248 277780
rect 147430 277766 147628 277794
rect 146668 275460 146720 275466
rect 146668 275402 146720 275408
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145564 274100 145616 274106
rect 145564 274042 145616 274048
rect 145012 273964 145064 273970
rect 145012 273906 145064 273912
rect 144644 273556 144696 273562
rect 144644 273498 144696 273504
rect 145104 272536 145156 272542
rect 145104 272478 145156 272484
rect 143908 272264 143960 272270
rect 143908 272206 143960 272212
rect 144736 268932 144788 268938
rect 144736 268874 144788 268880
rect 144552 267572 144604 267578
rect 144552 267514 144604 267520
rect 144564 267170 144592 267514
rect 144552 267164 144604 267170
rect 144552 267106 144604 267112
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 268874
rect 144920 267572 144972 267578
rect 144920 267514 144972 267520
rect 144932 266490 144960 267514
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 272478
rect 145576 266558 145604 274042
rect 146680 270094 146708 275402
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 146668 270088 146720 270094
rect 146668 270030 146720 270036
rect 145564 266552 145616 266558
rect 145564 266494 145616 266500
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 147600 268394 147628 277766
rect 148324 274236 148376 274242
rect 148324 274178 148376 274184
rect 147588 268388 147640 268394
rect 147588 268330 147640 268336
rect 147588 267980 147640 267986
rect 147588 267922 147640 267928
rect 147600 267170 147628 267922
rect 147404 267164 147456 267170
rect 147404 267106 147456 267112
rect 147588 267164 147640 267170
rect 147588 267106 147640 267112
rect 147416 267050 147444 267106
rect 147416 267022 147720 267050
rect 147220 266416 147272 266422
rect 147220 266358 147272 266364
rect 147232 264316 147260 266358
rect 147692 264330 147720 267022
rect 148336 266422 148364 274178
rect 148612 271182 148640 277780
rect 149808 274922 149836 277780
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 149888 274780 149940 274786
rect 149888 274722 149940 274728
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149900 267170 149928 274722
rect 151004 271318 151032 277780
rect 152004 272672 152056 272678
rect 152004 272614 152056 272620
rect 150992 271312 151044 271318
rect 150992 271254 151044 271260
rect 151084 270632 151136 270638
rect 151084 270574 151136 270580
rect 151096 267578 151124 270574
rect 151360 270088 151412 270094
rect 151360 270030 151412 270036
rect 150532 267572 150584 267578
rect 150532 267514 150584 267520
rect 151084 267572 151136 267578
rect 151084 267514 151136 267520
rect 149060 267164 149112 267170
rect 149060 267106 149112 267112
rect 149888 267164 149940 267170
rect 149888 267106 149940 267112
rect 149072 266626 149100 267106
rect 149060 266620 149112 266626
rect 149060 266562 149112 266568
rect 148876 266552 148928 266558
rect 148876 266494 148928 266500
rect 148324 266416 148376 266422
rect 148324 266358 148376 266364
rect 147692 264302 148074 264330
rect 148888 264316 148916 266494
rect 149704 266416 149756 266422
rect 149704 266358 149756 266364
rect 149716 264316 149744 266358
rect 150544 264316 150572 267514
rect 151372 264316 151400 270030
rect 152016 264330 152044 272614
rect 152200 272542 152228 277780
rect 152188 272536 152240 272542
rect 152188 272478 152240 272484
rect 153304 272134 153332 277780
rect 153292 272128 153344 272134
rect 153292 272070 153344 272076
rect 152648 271448 152700 271454
rect 152648 271390 152700 271396
rect 152660 264330 152688 271390
rect 153844 270088 153896 270094
rect 153844 270030 153896 270036
rect 152016 264302 152214 264330
rect 152660 264302 153042 264330
rect 153856 264316 153884 270030
rect 154500 269958 154528 277780
rect 155710 277766 155908 277794
rect 154488 269952 154540 269958
rect 154488 269894 154540 269900
rect 155880 268530 155908 277766
rect 156892 276010 156920 277780
rect 156880 276004 156932 276010
rect 156880 275946 156932 275952
rect 156604 275596 156656 275602
rect 156604 275538 156656 275544
rect 156052 272808 156104 272814
rect 156052 272750 156104 272756
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 155868 268524 155920 268530
rect 155868 268466 155920 268472
rect 154672 267708 154724 267714
rect 154672 267650 154724 267656
rect 154684 264316 154712 267650
rect 155512 264316 155540 268466
rect 156064 264330 156092 272750
rect 156616 266422 156644 275538
rect 157616 274644 157668 274650
rect 157616 274586 157668 274592
rect 157156 266756 157208 266762
rect 157156 266698 157208 266704
rect 156604 266416 156656 266422
rect 156604 266358 156656 266364
rect 156064 264302 156354 264330
rect 157168 264316 157196 266698
rect 157628 264330 157656 274586
rect 158088 274106 158116 277780
rect 159298 277766 159956 277794
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159928 270094 159956 277766
rect 160100 275732 160152 275738
rect 160100 275674 160152 275680
rect 160112 274242 160140 275674
rect 160480 275466 160508 277780
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161584 274718 161612 277780
rect 162124 275188 162176 275194
rect 162124 275130 162176 275136
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 160928 274372 160980 274378
rect 160928 274314 160980 274320
rect 160100 274236 160152 274242
rect 160100 274178 160152 274184
rect 159916 270088 159968 270094
rect 159916 270030 159968 270036
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 159824 267300 159876 267306
rect 159824 267242 159876 267248
rect 159836 266490 159864 267242
rect 159824 266484 159876 266490
rect 159824 266426 159876 266432
rect 159640 266416 159692 266422
rect 159640 266358 159692 266364
rect 159652 264316 159680 266358
rect 160480 264316 160508 268602
rect 160940 264330 160968 274314
rect 162136 267714 162164 275130
rect 162780 268666 162808 277780
rect 163976 275602 164004 277780
rect 163964 275596 164016 275602
rect 163964 275538 164016 275544
rect 163136 274712 163188 274718
rect 163136 274654 163188 274660
rect 163148 268802 163176 274654
rect 164240 274236 164292 274242
rect 164240 274178 164292 274184
rect 163320 273080 163372 273086
rect 163320 273022 163372 273028
rect 162952 268796 163004 268802
rect 162952 268738 163004 268744
rect 163136 268796 163188 268802
rect 163136 268738 163188 268744
rect 162768 268660 162820 268666
rect 162768 268602 162820 268608
rect 162124 267708 162176 267714
rect 162124 267650 162176 267656
rect 162124 266484 162176 266490
rect 162124 266426 162176 266432
rect 160940 264302 161322 264330
rect 162136 264316 162164 266426
rect 162964 264316 162992 268738
rect 163332 264330 163360 273022
rect 164252 264330 164280 274178
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 164988 264330 165016 271798
rect 165172 271454 165200 277780
rect 166382 277766 166948 277794
rect 165160 271448 165212 271454
rect 165160 271390 165212 271396
rect 166920 270230 166948 277766
rect 167564 273086 167592 277780
rect 167736 275460 167788 275466
rect 167736 275402 167788 275408
rect 167552 273080 167604 273086
rect 167552 273022 167604 273028
rect 166908 270224 166960 270230
rect 166908 270166 166960 270172
rect 166908 269408 166960 269414
rect 166908 269350 166960 269356
rect 166264 269068 166316 269074
rect 166264 269010 166316 269016
rect 163332 264302 163806 264330
rect 164252 264302 164634 264330
rect 164988 264302 165462 264330
rect 166276 264316 166304 269010
rect 166920 267306 166948 269350
rect 167748 267442 167776 275402
rect 168668 272678 168696 277780
rect 169878 277766 170168 277794
rect 169944 275868 169996 275874
rect 169944 275810 169996 275816
rect 169024 273216 169076 273222
rect 169024 273158 169076 273164
rect 168656 272672 168708 272678
rect 168656 272614 168708 272620
rect 168380 271584 168432 271590
rect 168380 271526 168432 271532
rect 167920 270360 167972 270366
rect 167920 270302 167972 270308
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 167736 267436 167788 267442
rect 167736 267378 167788 267384
rect 166908 267300 166960 267306
rect 166908 267242 166960 267248
rect 167104 264316 167132 267378
rect 167932 264316 167960 270302
rect 168392 264330 168420 271526
rect 169036 266762 169064 273158
rect 169576 267708 169628 267714
rect 169576 267650 169628 267656
rect 169024 266756 169076 266762
rect 169024 266698 169076 266704
rect 168392 264302 168774 264330
rect 169588 264316 169616 267650
rect 169956 264330 169984 275810
rect 170140 274718 170168 277766
rect 171060 275466 171088 277780
rect 172270 277766 172468 277794
rect 171048 275460 171100 275466
rect 171048 275402 171100 275408
rect 170128 274712 170180 274718
rect 170128 274654 170180 274660
rect 171784 272128 171836 272134
rect 171784 272070 171836 272076
rect 171232 270496 171284 270502
rect 171232 270438 171284 270444
rect 169956 264302 170430 264330
rect 171244 264316 171272 270438
rect 171796 267714 171824 272070
rect 172440 270366 172468 277766
rect 173164 274712 173216 274718
rect 173164 274654 173216 274660
rect 173176 270502 173204 274654
rect 173452 271590 173480 277780
rect 174662 277766 175136 277794
rect 173440 271584 173492 271590
rect 173440 271526 173492 271532
rect 173164 270496 173216 270502
rect 173164 270438 173216 270444
rect 172428 270360 172480 270366
rect 172428 270302 172480 270308
rect 173716 269680 173768 269686
rect 173716 269622 173768 269628
rect 171784 267708 171836 267714
rect 171784 267650 171836 267656
rect 172888 267572 172940 267578
rect 172888 267514 172940 267520
rect 172060 266756 172112 266762
rect 172060 266698 172112 266704
rect 172072 264316 172100 266698
rect 172900 264316 172928 267514
rect 173728 264316 173756 269622
rect 175108 267306 175136 277766
rect 175844 271862 175872 277780
rect 176752 274508 176804 274514
rect 176752 274450 176804 274456
rect 175832 271856 175884 271862
rect 175832 271798 175884 271804
rect 175280 271720 175332 271726
rect 175280 271662 175332 271668
rect 174544 267300 174596 267306
rect 174544 267242 174596 267248
rect 175096 267300 175148 267306
rect 175096 267242 175148 267248
rect 174556 264316 174584 267242
rect 175292 264330 175320 271662
rect 176200 268252 176252 268258
rect 176200 268194 176252 268200
rect 175292 264302 175398 264330
rect 176212 264316 176240 268194
rect 176764 264330 176792 274450
rect 176948 274242 176976 277780
rect 178144 275738 178172 277780
rect 178132 275732 178184 275738
rect 178132 275674 178184 275680
rect 176936 274236 176988 274242
rect 176936 274178 176988 274184
rect 177488 273828 177540 273834
rect 177488 273770 177540 273776
rect 177500 264330 177528 273770
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179340 268938 179368 277780
rect 180536 272814 180564 277780
rect 181732 275874 181760 277780
rect 181720 275868 181772 275874
rect 181720 275810 181772 275816
rect 182088 275052 182140 275058
rect 182088 274994 182140 275000
rect 180524 272808 180576 272814
rect 180524 272750 180576 272756
rect 179880 272400 179932 272406
rect 179880 272342 179932 272348
rect 179328 268932 179380 268938
rect 179328 268874 179380 268880
rect 179512 266620 179564 266626
rect 179512 266562 179564 266568
rect 179524 264316 179552 266562
rect 179892 264330 179920 272342
rect 181352 271040 181404 271046
rect 181352 270982 181404 270988
rect 181168 269816 181220 269822
rect 181168 269758 181220 269764
rect 179892 264302 180366 264330
rect 181180 264316 181208 269758
rect 181364 267734 181392 270982
rect 182100 269822 182128 274994
rect 182928 274514 182956 277780
rect 184138 277766 184796 277794
rect 183468 275324 183520 275330
rect 183468 275266 183520 275272
rect 182916 274508 182968 274514
rect 182916 274450 182968 274456
rect 182456 270904 182508 270910
rect 182456 270846 182508 270852
rect 182088 269816 182140 269822
rect 182088 269758 182140 269764
rect 182180 269272 182232 269278
rect 182180 269214 182232 269220
rect 181364 267706 181576 267734
rect 181548 264330 181576 267706
rect 182192 266422 182220 269214
rect 182180 266416 182232 266422
rect 182180 266358 182232 266364
rect 182468 264330 182496 270846
rect 183480 269550 183508 275266
rect 184204 273080 184256 273086
rect 184204 273022 184256 273028
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183652 268116 183704 268122
rect 183652 268058 183704 268064
rect 181548 264302 182022 264330
rect 182468 264302 182850 264330
rect 183664 264316 183692 268058
rect 184216 267034 184244 273022
rect 184768 269686 184796 277766
rect 185228 274718 185256 277780
rect 186424 275330 186452 277780
rect 186412 275324 186464 275330
rect 186412 275266 186464 275272
rect 185584 274916 185636 274922
rect 185584 274858 185636 274864
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 185032 273692 185084 273698
rect 185032 273634 185084 273640
rect 184756 269680 184808 269686
rect 184756 269622 184808 269628
rect 184020 267028 184072 267034
rect 184020 266970 184072 266976
rect 184204 267028 184256 267034
rect 184204 266970 184256 266976
rect 184032 266762 184060 266970
rect 184480 266892 184532 266898
rect 184480 266834 184532 266840
rect 184020 266756 184072 266762
rect 184020 266698 184072 266704
rect 184492 264316 184520 266834
rect 185044 264330 185072 273634
rect 185596 269074 185624 274858
rect 187148 274712 187200 274718
rect 187148 274654 187200 274660
rect 186964 269816 187016 269822
rect 186964 269758 187016 269764
rect 185584 269068 185636 269074
rect 185584 269010 185636 269016
rect 186136 266416 186188 266422
rect 186136 266358 186188 266364
rect 185044 264302 185334 264330
rect 186148 264316 186176 266358
rect 186976 264316 187004 269758
rect 187160 267578 187188 274654
rect 187620 273086 187648 277780
rect 188816 275330 188844 277780
rect 187792 275324 187844 275330
rect 187792 275266 187844 275272
rect 188804 275324 188856 275330
rect 188804 275266 188856 275272
rect 187804 274378 187832 275266
rect 187792 274372 187844 274378
rect 187792 274314 187844 274320
rect 187792 273556 187844 273562
rect 187792 273498 187844 273504
rect 187608 273080 187660 273086
rect 187608 273022 187660 273028
rect 187804 272898 187832 273498
rect 187712 272870 187832 272898
rect 189816 272944 189868 272950
rect 189816 272886 189868 272892
rect 187332 269816 187384 269822
rect 187332 269758 187384 269764
rect 187344 269550 187372 269758
rect 187332 269544 187384 269550
rect 187332 269486 187384 269492
rect 187148 267572 187200 267578
rect 187148 267514 187200 267520
rect 187712 265674 187740 272870
rect 187884 270768 187936 270774
rect 187884 270710 187936 270716
rect 187700 265668 187752 265674
rect 187700 265610 187752 265616
rect 187896 265554 187924 270710
rect 189448 266756 189500 266762
rect 189448 266698 189500 266704
rect 188252 265668 188304 265674
rect 188252 265610 188304 265616
rect 187804 265526 187924 265554
rect 187804 264316 187832 265526
rect 188264 264330 188292 265610
rect 188264 264302 188646 264330
rect 189460 264316 189488 266698
rect 189828 264330 189856 272886
rect 190012 271046 190040 277780
rect 191208 272950 191236 277780
rect 191196 272944 191248 272950
rect 191196 272886 191248 272892
rect 190736 272264 190788 272270
rect 190736 272206 190788 272212
rect 190000 271040 190052 271046
rect 190000 270982 190052 270988
rect 190748 264330 190776 272206
rect 192312 271726 192340 277780
rect 193508 273970 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 193864 276004 193916 276010
rect 193864 275946 193916 275952
rect 192484 273964 192536 273970
rect 192484 273906 192536 273912
rect 193496 273964 193548 273970
rect 193496 273906 193548 273912
rect 192300 271720 192352 271726
rect 192300 271662 192352 271668
rect 191932 269816 191984 269822
rect 191932 269758 191984 269764
rect 189828 264302 190302 264330
rect 190748 264302 191130 264330
rect 191944 264316 191972 269758
rect 192496 264330 192524 273906
rect 193588 268388 193640 268394
rect 193588 268330 193640 268336
rect 192496 264302 192786 264330
rect 193600 264316 193628 268330
rect 193876 267034 193904 275946
rect 194612 269822 194640 277366
rect 195900 274650 195928 277780
rect 197110 277766 197308 277794
rect 198306 277766 198688 277794
rect 195888 274644 195940 274650
rect 195888 274586 195940 274592
rect 195980 271312 196032 271318
rect 195980 271254 196032 271260
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 193864 267028 193916 267034
rect 193864 266970 193916 266976
rect 194428 264316 194456 267106
rect 194796 264330 194824 271118
rect 195992 264330 196020 271254
rect 196900 269068 196952 269074
rect 196900 269010 196952 269016
rect 194796 264302 195270 264330
rect 195992 264302 196098 264330
rect 196912 264316 196940 269010
rect 197280 268394 197308 277766
rect 197544 272536 197596 272542
rect 197544 272478 197596 272484
rect 197268 268388 197320 268394
rect 197268 268330 197320 268336
rect 197556 264330 197584 272478
rect 198660 269958 198688 277766
rect 199488 272542 199516 277780
rect 200592 277394 200620 277780
rect 200500 277366 200620 277394
rect 199660 274508 199712 274514
rect 199660 274450 199712 274456
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 198188 269952 198240 269958
rect 198188 269894 198240 269900
rect 198648 269952 198700 269958
rect 198648 269894 198700 269900
rect 198200 264330 198228 269894
rect 199384 267708 199436 267714
rect 199384 267650 199436 267656
rect 197556 264302 197754 264330
rect 198200 264302 198582 264330
rect 199396 264316 199424 267650
rect 199672 267170 199700 274450
rect 200500 270910 200528 277366
rect 201788 276010 201816 277780
rect 201776 276004 201828 276010
rect 201776 275946 201828 275952
rect 202144 275596 202196 275602
rect 202144 275538 202196 275544
rect 200672 274100 200724 274106
rect 200672 274042 200724 274048
rect 200488 270904 200540 270910
rect 200488 270846 200540 270852
rect 200212 268524 200264 268530
rect 200212 268466 200264 268472
rect 199660 267164 199712 267170
rect 199660 267106 199712 267112
rect 200224 264316 200252 268466
rect 200684 264330 200712 274042
rect 201868 267028 201920 267034
rect 201868 266970 201920 266976
rect 200684 264302 201066 264330
rect 201880 264316 201908 266970
rect 202156 266422 202184 275538
rect 202696 270088 202748 270094
rect 202696 270030 202748 270036
rect 202144 266416 202196 266422
rect 202144 266358 202196 266364
rect 202708 264316 202736 270030
rect 202984 268530 203012 277780
rect 203996 277766 204194 277794
rect 205390 277766 205588 277794
rect 203996 268802 204024 277766
rect 205560 270094 205588 277766
rect 206284 274644 206336 274650
rect 206284 274586 206336 274592
rect 205732 271448 205784 271454
rect 205732 271390 205784 271396
rect 205548 270088 205600 270094
rect 205548 270030 205600 270036
rect 203524 268796 203576 268802
rect 203524 268738 203576 268744
rect 203984 268796 204036 268802
rect 203984 268738 204036 268744
rect 202972 268524 203024 268530
rect 202972 268466 203024 268472
rect 203536 264316 203564 268738
rect 205180 268660 205232 268666
rect 205180 268602 205232 268608
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 205192 264316 205220 268602
rect 205744 264330 205772 271390
rect 206296 267034 206324 274586
rect 206572 274106 206600 277780
rect 207782 277766 208348 277794
rect 206560 274100 206612 274106
rect 206560 274042 206612 274048
rect 207664 271856 207716 271862
rect 207664 271798 207716 271804
rect 207388 270224 207440 270230
rect 207388 270166 207440 270172
rect 206284 267028 206336 267034
rect 206284 266970 206336 266976
rect 206836 266416 206888 266422
rect 206836 266358 206888 266364
rect 205744 264302 206034 264330
rect 206848 264316 206876 266358
rect 207400 264330 207428 270166
rect 207676 267714 207704 271798
rect 208320 269550 208348 277766
rect 208492 272672 208544 272678
rect 208492 272614 208544 272620
rect 208308 269544 208360 269550
rect 208308 269486 208360 269492
rect 207664 267708 207716 267714
rect 207664 267650 207716 267656
rect 207400 264302 207690 264330
rect 208504 264316 208532 272614
rect 208872 271182 208900 277780
rect 210068 274514 210096 277780
rect 210792 275460 210844 275466
rect 210792 275402 210844 275408
rect 210056 274508 210108 274514
rect 210056 274450 210108 274456
rect 208860 271176 208912 271182
rect 208860 271118 208912 271124
rect 210804 270502 210832 275402
rect 211264 273086 211292 277780
rect 211988 273216 212040 273222
rect 211988 273158 212040 273164
rect 211252 273080 211304 273086
rect 211252 273022 211304 273028
rect 210148 270496 210200 270502
rect 210148 270438 210200 270444
rect 210792 270496 210844 270502
rect 210792 270438 210844 270444
rect 211804 270496 211856 270502
rect 211804 270438 211856 270444
rect 208676 270360 208728 270366
rect 208676 270302 208728 270308
rect 208688 266490 208716 270302
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 208676 266484 208728 266490
rect 208676 266426 208728 266432
rect 209332 264316 209360 266834
rect 210160 264316 210188 270438
rect 210976 266484 211028 266490
rect 210976 266426 211028 266432
rect 210988 264316 211016 266426
rect 211816 264316 211844 270438
rect 212000 267442 212028 273158
rect 212460 270366 212488 277780
rect 213670 277766 213868 277794
rect 212632 271584 212684 271590
rect 212632 271526 212684 271532
rect 212448 270360 212500 270366
rect 212448 270302 212500 270308
rect 211988 267436 212040 267442
rect 211988 267378 212040 267384
rect 212644 264316 212672 271526
rect 213840 270230 213868 277766
rect 214656 274236 214708 274242
rect 214656 274178 214708 274184
rect 213828 270224 213880 270230
rect 213828 270166 213880 270172
rect 213828 269680 213880 269686
rect 213828 269622 213880 269628
rect 213460 267708 213512 267714
rect 213460 267650 213512 267656
rect 213472 264316 213500 267650
rect 213840 266626 213868 269622
rect 214288 267300 214340 267306
rect 214288 267242 214340 267248
rect 213828 266620 213880 266626
rect 213828 266562 213880 266568
rect 214300 264316 214328 267242
rect 214668 264330 214696 274178
rect 214852 271862 214880 277780
rect 214840 271856 214892 271862
rect 214840 271798 214892 271804
rect 215956 271318 215984 277780
rect 217166 277766 217456 277794
rect 216864 275732 216916 275738
rect 216864 275674 216916 275680
rect 215944 271312 215996 271318
rect 215944 271254 215996 271260
rect 216128 271040 216180 271046
rect 216128 270982 216180 270988
rect 215944 268932 215996 268938
rect 215944 268874 215996 268880
rect 214668 264302 215142 264330
rect 215956 264316 215984 268874
rect 216140 267714 216168 270982
rect 216876 267734 216904 275674
rect 217232 272808 217284 272814
rect 217232 272750 217284 272756
rect 216128 267708 216180 267714
rect 216128 267650 216180 267656
rect 216784 267706 216904 267734
rect 216784 264316 216812 267706
rect 217244 264330 217272 272750
rect 217428 272678 217456 277766
rect 218348 275466 218376 277780
rect 218888 275868 218940 275874
rect 218888 275810 218940 275816
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217416 272672 217468 272678
rect 217416 272614 217468 272620
rect 218428 267164 218480 267170
rect 218428 267106 218480 267112
rect 217244 264302 217626 264330
rect 218440 264316 218468 267106
rect 218900 264330 218928 275810
rect 219544 268666 219572 277780
rect 220556 277766 220754 277794
rect 220556 274242 220584 277766
rect 221936 275602 221964 277780
rect 223146 277766 223528 277794
rect 223500 276026 223528 277766
rect 222108 276004 222160 276010
rect 223500 275998 223620 276026
rect 222108 275946 222160 275952
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 220912 274372 220964 274378
rect 220912 274314 220964 274320
rect 220544 274236 220596 274242
rect 220544 274178 220596 274184
rect 220084 273080 220136 273086
rect 220084 273022 220136 273028
rect 219532 268660 219584 268666
rect 219532 268602 219584 268608
rect 220096 267306 220124 273022
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 220084 266620 220136 266626
rect 220084 266562 220136 266568
rect 218900 264302 219282 264330
rect 220096 264316 220124 266562
rect 220924 264316 220952 274314
rect 222120 271862 222148 275946
rect 222844 275324 222896 275330
rect 222844 275266 222896 275272
rect 221464 271856 221516 271862
rect 221464 271798 221516 271804
rect 222108 271856 222160 271862
rect 222108 271798 222160 271804
rect 221476 267170 221504 271798
rect 221740 267572 221792 267578
rect 221740 267514 221792 267520
rect 221464 267164 221516 267170
rect 221464 267106 221516 267112
rect 221752 264316 221780 267514
rect 222568 267436 222620 267442
rect 222568 267378 222620 267384
rect 222580 264316 222608 267378
rect 222856 266422 222884 275266
rect 223592 271454 223620 275998
rect 224236 275126 224264 277780
rect 225432 275330 225460 277780
rect 225420 275324 225472 275330
rect 225420 275266 225472 275272
rect 224224 275120 224276 275126
rect 224224 275062 224276 275068
rect 226156 275120 226208 275126
rect 226156 275062 226208 275068
rect 224868 272944 224920 272950
rect 224920 272892 225000 272898
rect 224868 272886 225000 272892
rect 224880 272870 225000 272886
rect 223580 271448 223632 271454
rect 223580 271390 223632 271396
rect 224224 270904 224276 270910
rect 224224 270846 224276 270852
rect 223396 267708 223448 267714
rect 223396 267650 223448 267656
rect 222844 266416 222896 266422
rect 222844 266358 222896 266364
rect 223408 264316 223436 267650
rect 224236 267442 224264 270846
rect 224224 267436 224276 267442
rect 224224 267378 224276 267384
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 224236 264316 224264 266358
rect 224972 264330 225000 272870
rect 225512 271720 225564 271726
rect 225512 271662 225564 271668
rect 225524 264330 225552 271662
rect 226168 271590 226196 275062
rect 226340 273964 226392 273970
rect 226340 273906 226392 273912
rect 226156 271584 226208 271590
rect 226156 271526 226208 271532
rect 226352 264330 226380 273906
rect 226628 269686 226656 277780
rect 227824 277394 227852 277780
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 227824 277366 227944 277394
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 227272 264330 227300 269758
rect 227916 268802 227944 277366
rect 228836 272814 228864 277766
rect 228824 272808 228876 272814
rect 228824 272750 228876 272756
rect 230400 269958 230428 277766
rect 231412 272542 231440 277780
rect 232530 277766 233188 277794
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 230020 269952 230072 269958
rect 230020 269894 230072 269900
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 227720 268796 227772 268802
rect 227720 268738 227772 268744
rect 227904 268796 227956 268802
rect 227904 268738 227956 268744
rect 227732 267578 227760 268738
rect 229192 268388 229244 268394
rect 229192 268330 229244 268336
rect 227720 267572 227772 267578
rect 227720 267514 227772 267520
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226352 264302 226734 264330
rect 227272 264302 227562 264330
rect 228376 264316 228404 266970
rect 229204 264316 229232 268330
rect 230032 264316 230060 269894
rect 230584 264330 230612 272478
rect 232136 271856 232188 271862
rect 232136 271798 232188 271804
rect 230756 269544 230808 269550
rect 230756 269486 230808 269492
rect 230768 266422 230796 269486
rect 231676 267436 231728 267442
rect 231676 267378 231728 267384
rect 230756 266416 230808 266422
rect 230756 266358 230808 266364
rect 230584 264302 230874 264330
rect 231688 264316 231716 267378
rect 232148 264330 232176 271798
rect 233160 270502 233188 277766
rect 233148 270496 233200 270502
rect 233148 270438 233200 270444
rect 233332 268524 233384 268530
rect 233332 268466 233384 268472
rect 232148 264302 232530 264330
rect 233344 264316 233372 268466
rect 233712 268394 233740 277780
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 268388 233752 268394
rect 233700 268330 233752 268336
rect 233896 267442 233924 275538
rect 234908 273970 234936 277780
rect 236104 275602 236132 277780
rect 236092 275596 236144 275602
rect 236092 275538 236144 275544
rect 235448 274100 235500 274106
rect 235448 274042 235500 274048
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 234988 270088 235040 270094
rect 234988 270030 235040 270036
rect 234160 267572 234212 267578
rect 234160 267514 234212 267520
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234172 264316 234200 267514
rect 235000 264316 235028 270030
rect 235460 264330 235488 274042
rect 237300 270638 237328 277780
rect 237472 275460 237524 275466
rect 237472 275402 237524 275408
rect 237484 271726 237512 275402
rect 238496 274718 238524 277780
rect 238484 274712 238536 274718
rect 238484 274654 238536 274660
rect 237840 274508 237892 274514
rect 237840 274450 237892 274456
rect 237472 271720 237524 271726
rect 237472 271662 237524 271668
rect 237472 271176 237524 271182
rect 237472 271118 237524 271124
rect 237288 270632 237340 270638
rect 237288 270574 237340 270580
rect 237288 270496 237340 270502
rect 237288 270438 237340 270444
rect 237300 267034 237328 270438
rect 237288 267028 237340 267034
rect 237288 266970 237340 266976
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237484 264316 237512 271118
rect 237852 264330 237880 274450
rect 239600 274106 239628 277780
rect 239772 274712 239824 274718
rect 239772 274654 239824 274660
rect 239588 274100 239640 274106
rect 239588 274042 239640 274048
rect 239784 270094 239812 274654
rect 240600 274236 240652 274242
rect 240600 274178 240652 274184
rect 240612 270994 240640 274178
rect 240796 271182 240824 277780
rect 242006 277766 242388 277794
rect 242360 272678 242388 277766
rect 242164 272672 242216 272678
rect 242164 272614 242216 272620
rect 242348 272672 242400 272678
rect 242348 272614 242400 272620
rect 242176 271402 242204 272614
rect 242176 271374 242296 271402
rect 242072 271312 242124 271318
rect 242072 271254 242124 271260
rect 240784 271176 240836 271182
rect 240784 271118 240836 271124
rect 240612 270966 240732 270994
rect 239956 270360 240008 270366
rect 239956 270302 240008 270308
rect 239772 270088 239824 270094
rect 239772 270030 239824 270036
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 237852 264302 238326 264330
rect 239140 264316 239168 267242
rect 239968 264316 239996 270302
rect 240508 270224 240560 270230
rect 240508 270166 240560 270172
rect 240520 264330 240548 270166
rect 240704 266762 240732 270966
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 240692 266756 240744 266762
rect 240692 266698 240744 266704
rect 240520 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271254
rect 242268 266422 242296 271374
rect 243188 271318 243216 277780
rect 244384 275466 244412 277780
rect 244372 275460 244424 275466
rect 244372 275402 244424 275408
rect 245108 275324 245160 275330
rect 245108 275266 245160 275272
rect 243728 271720 243780 271726
rect 243728 271662 243780 271668
rect 243176 271312 243228 271318
rect 243176 271254 243228 271260
rect 242256 266416 242308 266422
rect 242256 266358 242308 266364
rect 243268 266416 243320 266422
rect 243268 266358 243320 266364
rect 242084 264302 242466 264330
rect 243280 264316 243308 266358
rect 243740 264330 243768 271662
rect 244924 268660 244976 268666
rect 244924 268602 244976 268608
rect 243740 264302 244122 264330
rect 244936 264316 244964 268602
rect 245120 266626 245148 275266
rect 245580 268530 245608 277780
rect 246790 277766 246988 277794
rect 245568 268524 245620 268530
rect 245568 268466 245620 268472
rect 246580 267436 246632 267442
rect 246580 267378 246632 267384
rect 245752 266756 245804 266762
rect 245752 266698 245804 266704
rect 245108 266620 245160 266626
rect 245108 266562 245160 266568
rect 245764 264316 245792 266698
rect 246592 264316 246620 267378
rect 246960 267170 246988 277766
rect 247224 271584 247276 271590
rect 247224 271526 247276 271532
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 247236 265674 247264 271526
rect 247880 271454 247908 277780
rect 249090 277766 249656 277794
rect 249064 272808 249116 272814
rect 249064 272750 249116 272756
rect 247408 271448 247460 271454
rect 247408 271390 247460 271396
rect 247868 271448 247920 271454
rect 247868 271390 247920 271396
rect 247224 265668 247276 265674
rect 247224 265610 247276 265616
rect 247420 264316 247448 271390
rect 249076 266762 249104 272750
rect 249628 270230 249656 277766
rect 250272 275330 250300 277780
rect 251088 275596 251140 275602
rect 251088 275538 251140 275544
rect 250260 275324 250312 275330
rect 250260 275266 250312 275272
rect 249616 270224 249668 270230
rect 249616 270166 249668 270172
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 249064 266756 249116 266762
rect 249064 266698 249116 266704
rect 249064 266620 249116 266626
rect 249064 266562 249116 266568
rect 247868 265668 247920 265674
rect 247868 265610 247920 265616
rect 247880 264330 247908 265610
rect 247880 264302 248262 264330
rect 249076 264316 249104 266562
rect 249904 264316 249932 269758
rect 251100 269074 251128 275538
rect 251468 269822 251496 277780
rect 252678 277766 252968 277794
rect 252940 272542 252968 277766
rect 252744 272536 252796 272542
rect 252744 272478 252796 272484
rect 252928 272536 252980 272542
rect 252928 272478 252980 272484
rect 252008 270496 252060 270502
rect 252008 270438 252060 270444
rect 251456 269816 251508 269822
rect 251456 269758 251508 269764
rect 251088 269068 251140 269074
rect 251088 269010 251140 269016
rect 250720 268796 250772 268802
rect 250720 268738 250772 268744
rect 250732 264316 250760 268738
rect 251548 266756 251600 266762
rect 251548 266698 251600 266704
rect 251560 264316 251588 266698
rect 252020 266422 252048 270438
rect 252376 269952 252428 269958
rect 252376 269894 252428 269900
rect 252008 266416 252060 266422
rect 252008 266358 252060 266364
rect 252388 264316 252416 269894
rect 252756 264330 252784 272478
rect 253860 270366 253888 277780
rect 254584 275460 254636 275466
rect 254584 275402 254636 275408
rect 253848 270360 253900 270366
rect 253848 270302 253900 270308
rect 253204 270088 253256 270094
rect 253204 270030 253256 270036
rect 253216 269686 253244 270030
rect 253204 269680 253256 269686
rect 253204 269622 253256 269628
rect 254596 267306 254624 275402
rect 255056 274666 255084 277780
rect 255056 274638 255360 274666
rect 255332 268394 255360 274638
rect 256160 273970 256188 277780
rect 257370 277766 258028 277794
rect 255504 273964 255556 273970
rect 255504 273906 255556 273912
rect 256148 273964 256200 273970
rect 256148 273906 256200 273912
rect 254860 268388 254912 268394
rect 254860 268330 254912 268336
rect 255320 268388 255372 268394
rect 255320 268330 255372 268336
rect 254584 267300 254636 267306
rect 254584 267242 254636 267248
rect 254032 267028 254084 267034
rect 254032 266970 254084 266976
rect 252756 264302 253230 264330
rect 254044 264316 254072 266970
rect 254872 264316 254900 268330
rect 255516 264330 255544 273906
rect 256516 269068 256568 269074
rect 256516 269010 256568 269016
rect 255516 264302 255714 264330
rect 256528 264316 256556 269010
rect 258000 266898 258028 277766
rect 258552 277394 258580 277780
rect 258460 277366 258580 277394
rect 258460 269958 258488 277366
rect 258632 274100 258684 274106
rect 258632 274042 258684 274048
rect 258448 269952 258500 269958
rect 258448 269894 258500 269900
rect 258172 269680 258224 269686
rect 258172 269622 258224 269628
rect 257988 266892 258040 266898
rect 257988 266834 258040 266840
rect 257344 266416 257396 266422
rect 257344 266358 257396 266364
rect 257356 264316 257384 266358
rect 258184 264316 258212 269622
rect 258644 264330 258672 274042
rect 259552 272672 259604 272678
rect 259552 272614 259604 272620
rect 259564 265674 259592 272614
rect 259748 271590 259776 277780
rect 260944 275466 260972 277780
rect 260932 275460 260984 275466
rect 260932 275402 260984 275408
rect 259736 271584 259788 271590
rect 259736 271526 259788 271532
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 259828 271176 259880 271182
rect 259828 271118 259880 271124
rect 259552 265668 259604 265674
rect 259552 265610 259604 265616
rect 258644 264302 259026 264330
rect 259840 264316 259868 271118
rect 260380 265668 260432 265674
rect 260380 265610 260432 265616
rect 260392 264330 260420 265610
rect 261036 264330 261064 271254
rect 262140 271182 262168 277780
rect 263258 277766 263548 277794
rect 264454 277766 264928 277794
rect 265650 277766 266216 277794
rect 262128 271176 262180 271182
rect 262128 271118 262180 271124
rect 263324 270224 263376 270230
rect 263324 270166 263376 270172
rect 263140 268524 263192 268530
rect 263140 268466 263192 268472
rect 262312 267300 262364 267306
rect 262312 267242 262364 267248
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262324 264316 262352 267242
rect 263152 264316 263180 268466
rect 263336 266422 263364 270166
rect 263520 268530 263548 277766
rect 264336 271448 264388 271454
rect 264336 271390 264388 271396
rect 263508 268524 263560 268530
rect 263508 268466 263560 268472
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263324 266416 263376 266422
rect 263324 266358 263376 266364
rect 263980 264316 264008 267106
rect 264348 264330 264376 271390
rect 264900 269278 264928 277766
rect 265072 270360 265124 270366
rect 265072 270302 265124 270308
rect 264888 269272 264940 269278
rect 264888 269214 264940 269220
rect 265084 266830 265112 270302
rect 266188 270094 266216 277766
rect 266832 275330 266860 277780
rect 266360 275324 266412 275330
rect 266360 275266 266412 275272
rect 266820 275324 266872 275330
rect 266820 275266 266872 275272
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 265072 266824 265124 266830
rect 265072 266766 265124 266772
rect 265624 266416 265676 266422
rect 265624 266358 265676 266364
rect 264348 264302 264822 264330
rect 265636 264316 265664 266358
rect 266372 264330 266400 275266
rect 268028 272542 268056 277780
rect 267740 272536 267792 272542
rect 267740 272478 267792 272484
rect 268016 272536 268068 272542
rect 268016 272478 268068 272484
rect 267280 269816 267332 269822
rect 267280 269758 267332 269764
rect 266372 264302 266478 264330
rect 267292 264316 267320 269758
rect 267752 264330 267780 272478
rect 269224 270230 269252 277780
rect 270420 277394 270448 277780
rect 270328 277366 270448 277394
rect 269212 270224 269264 270230
rect 269212 270166 269264 270172
rect 270328 269822 270356 277366
rect 271524 273970 271552 277780
rect 272734 277766 273116 277794
rect 270592 273964 270644 273970
rect 270592 273906 270644 273912
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270316 269816 270368 269822
rect 270316 269758 270368 269764
rect 269120 269272 269172 269278
rect 269120 269214 269172 269220
rect 268936 266824 268988 266830
rect 268936 266766 268988 266772
rect 267752 264302 268134 264330
rect 268948 264316 268976 266766
rect 269132 266422 269160 269214
rect 269764 268388 269816 268394
rect 269764 268330 269816 268336
rect 269120 266416 269172 266422
rect 269120 266358 269172 266364
rect 269776 264316 269804 268330
rect 270604 264316 270632 273906
rect 272616 271584 272668 271590
rect 272616 271526 272668 271532
rect 272248 269952 272300 269958
rect 272248 269894 272300 269900
rect 271420 267028 271472 267034
rect 271420 266970 271472 266976
rect 271432 264316 271460 266970
rect 272260 264316 272288 269894
rect 272628 264330 272656 271526
rect 273088 269958 273116 277766
rect 273916 275466 273944 277780
rect 273536 275460 273588 275466
rect 273536 275402 273588 275408
rect 273904 275460 273956 275466
rect 273904 275402 273956 275408
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 273548 264330 273576 275402
rect 275112 271318 275140 277780
rect 275100 271312 275152 271318
rect 275100 271254 275152 271260
rect 276308 271182 276336 277780
rect 276664 275324 276716 275330
rect 276664 275266 276716 275272
rect 274640 271176 274692 271182
rect 274640 271118 274692 271124
rect 276296 271176 276348 271182
rect 276296 271118 276348 271124
rect 274652 264330 274680 271118
rect 275560 268524 275612 268530
rect 275560 268466 275612 268472
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 268466
rect 276676 267034 276704 275266
rect 277504 274990 277532 277780
rect 278700 277394 278728 277780
rect 278608 277366 278728 277394
rect 277492 274984 277544 274990
rect 277492 274926 277544 274932
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276664 267028 276716 267034
rect 276664 266970 276716 266976
rect 276388 266416 276440 266422
rect 276388 266358 276440 266364
rect 276400 264316 276428 266358
rect 277228 264316 277256 270030
rect 278044 267028 278096 267034
rect 278044 266970 278096 266976
rect 278056 264316 278084 266970
rect 278608 266422 278636 277366
rect 279804 272542 279832 277780
rect 280804 273964 280856 273970
rect 280804 273906 280856 273912
rect 278780 272536 278832 272542
rect 278780 272478 278832 272484
rect 279792 272536 279844 272542
rect 279792 272478 279844 272484
rect 278596 266416 278648 266422
rect 278596 266358 278648 266364
rect 278792 264330 278820 272478
rect 279700 270224 279752 270230
rect 279700 270166 279752 270172
rect 278792 264302 278898 264330
rect 279712 264316 279740 270166
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280540 264316 280568 269758
rect 280816 267734 280844 273906
rect 281000 273766 281028 277780
rect 282210 277766 282776 277794
rect 280988 273760 281040 273766
rect 280988 273702 281040 273708
rect 282184 269952 282236 269958
rect 282184 269894 282236 269900
rect 280816 267706 280936 267734
rect 280908 264330 280936 267706
rect 280908 264302 281382 264330
rect 282196 264316 282224 269894
rect 282748 269142 282776 277766
rect 282920 275460 282972 275466
rect 282920 275402 282972 275408
rect 282736 269136 282788 269142
rect 282736 269078 282788 269084
rect 282932 264330 282960 275402
rect 283392 274854 283420 277780
rect 284588 275330 284616 277780
rect 284576 275324 284628 275330
rect 284576 275266 284628 275272
rect 284300 274984 284352 274990
rect 284300 274926 284352 274932
rect 283380 274848 283432 274854
rect 283380 274790 283432 274796
rect 283472 271312 283524 271318
rect 283472 271254 283524 271260
rect 283484 264330 283512 271254
rect 284312 265674 284340 274926
rect 285784 274718 285812 277780
rect 286888 277394 286916 277780
rect 286796 277366 286916 277394
rect 285772 274712 285824 274718
rect 285772 274654 285824 274660
rect 284484 271176 284536 271182
rect 284484 271118 284536 271124
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271118
rect 286796 269958 286824 277366
rect 286968 274712 287020 274718
rect 286968 274654 287020 274660
rect 286784 269952 286836 269958
rect 286784 269894 286836 269900
rect 286980 267034 287008 274654
rect 287520 273760 287572 273766
rect 287520 273702 287572 273708
rect 287152 272536 287204 272542
rect 287152 272478 287204 272484
rect 286968 267028 287020 267034
rect 286968 266970 287020 266976
rect 286324 266416 286376 266422
rect 286324 266358 286376 266364
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 286336 264316 286364 266358
rect 287164 264316 287192 272478
rect 287532 264330 287560 273702
rect 288084 272950 288112 277780
rect 289280 274922 289308 277780
rect 290096 275324 290148 275330
rect 290096 275266 290148 275272
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289084 274848 289136 274854
rect 289084 274790 289136 274796
rect 288072 272944 288124 272950
rect 288072 272886 288124 272892
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 287532 264302 288006 264330
rect 288820 264316 288848 269078
rect 289096 267734 289124 274790
rect 289096 267706 289216 267734
rect 289188 264330 289216 267706
rect 290108 264330 290136 275266
rect 290476 274718 290504 277780
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 290464 272944 290516 272950
rect 290464 272886 290516 272892
rect 290476 266422 290504 272886
rect 291672 270366 291700 277780
rect 292868 270502 292896 277780
rect 294064 275126 294092 277780
rect 295168 275210 295196 277780
rect 295168 275182 295380 275210
rect 294052 275120 294104 275126
rect 294052 275062 294104 275068
rect 295156 275120 295208 275126
rect 295156 275062 295208 275068
rect 293408 274916 293460 274922
rect 293408 274858 293460 274864
rect 292856 270496 292908 270502
rect 292856 270438 292908 270444
rect 291660 270360 291712 270366
rect 291660 270302 291712 270308
rect 292120 269952 292172 269958
rect 292120 269894 292172 269900
rect 291292 267028 291344 267034
rect 291292 266970 291344 266976
rect 290464 266416 290516 266422
rect 290464 266358 290516 266364
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 266970
rect 292132 264316 292160 269894
rect 292948 266416 293000 266422
rect 292948 266358 293000 266364
rect 292960 264316 292988 266358
rect 293420 264330 293448 274858
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 294156 264330 294184 274654
rect 295168 267034 295196 275062
rect 295352 269142 295380 275182
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 296260 270496 296312 270502
rect 296260 270438 296312 270444
rect 295524 270360 295576 270366
rect 295524 270302 295576 270308
rect 295340 269136 295392 269142
rect 295340 269078 295392 269084
rect 295536 267734 295564 270302
rect 295444 267706 295564 267734
rect 295156 267028 295208 267034
rect 295156 266970 295208 266976
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295444 264316 295472 267706
rect 296272 264316 296300 270438
rect 297548 269136 297600 269142
rect 297548 269078 297600 269084
rect 297088 267028 297140 267034
rect 297088 266970 297140 266976
rect 297100 264316 297128 266970
rect 297560 264330 297588 269078
rect 297928 266422 297956 277766
rect 298756 275398 298784 277780
rect 299952 275738 299980 277780
rect 300964 277766 301162 277794
rect 299940 275732 299992 275738
rect 299940 275674 299992 275680
rect 300768 275732 300820 275738
rect 300768 275674 300820 275680
rect 298744 275392 298796 275398
rect 298744 275334 298796 275340
rect 300032 275392 300084 275398
rect 300032 275334 300084 275340
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 297916 266416 297968 266422
rect 297916 266358 297968 266364
rect 298388 264330 298416 274654
rect 299572 266416 299624 266422
rect 299572 266358 299624 266364
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 266358
rect 300044 264330 300072 275334
rect 300780 267734 300808 275674
rect 300964 267734 300992 277766
rect 302344 277394 302372 277780
rect 303448 277394 303476 277780
rect 303724 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 302344 277366 302464 277394
rect 303448 277366 303568 277394
rect 300780 267706 300900 267734
rect 300964 267706 301084 267734
rect 300872 264330 300900 267706
rect 301056 266422 301084 267706
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303540 267734 303568 277366
rect 303724 267734 303752 277766
rect 303540 267706 303660 267734
rect 303724 267706 304120 267734
rect 303632 264330 303660 267706
rect 304092 264330 304120 267706
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 316052 277766 316526 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 267300 312872 267306
rect 312820 267242 312872 267248
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312360 266416 312412 266422
rect 312360 266358 312412 266364
rect 312372 264330 312400 266358
rect 312018 264302 312400 264330
rect 312832 264316 312860 267242
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313648 267572 313700 267578
rect 313648 267514 313700 267520
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313660 264316 313688 267514
rect 314488 264316 314516 269758
rect 314672 266422 314700 277766
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266416 314712 266422
rect 314660 266358 314712 266364
rect 315776 264330 315804 271254
rect 316052 267306 316080 277766
rect 317708 277394 317736 277780
rect 317708 277366 317828 277394
rect 316960 270292 317012 270298
rect 316960 270234 317012 270240
rect 316040 267300 316092 267306
rect 316040 267242 316092 267248
rect 316132 267028 316184 267034
rect 316132 266970 316184 266976
rect 315330 264302 315804 264330
rect 316144 264316 316172 266970
rect 316972 264316 317000 270234
rect 317800 267578 317828 277366
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317788 267572 317840 267578
rect 317788 267514 317840 267520
rect 317788 266416 317840 266422
rect 317788 266358 317840 266364
rect 317800 264316 317828 266358
rect 318628 264316 318656 271730
rect 318812 269822 318840 277780
rect 320008 271318 320036 277780
rect 320192 277766 321218 277794
rect 321572 277766 322414 277794
rect 323136 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318800 269816 318852 269822
rect 318800 269758 318852 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320192 267034 320220 277766
rect 321572 270298 321600 277766
rect 321560 270292 321612 270298
rect 321560 270234 321612 270240
rect 321928 270224 321980 270230
rect 321928 270166 321980 270172
rect 321100 269272 321152 269278
rect 321100 269214 321152 269220
rect 320180 267028 320232 267034
rect 320180 266970 320232 266976
rect 320272 266892 320324 266898
rect 320272 266834 320324 266840
rect 320284 264316 320312 266834
rect 321112 264316 321140 269214
rect 321940 264316 321968 270166
rect 322756 268388 322808 268394
rect 322756 268330 322808 268336
rect 322768 264316 322796 268330
rect 323136 266422 323164 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 327106 277766 327488 277794
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 325516 271312 325568 271318
rect 325516 271254 325568 271260
rect 323584 270088 323636 270094
rect 323584 270030 323636 270036
rect 323124 266416 323176 266422
rect 323124 266358 323176 266364
rect 323596 264316 323624 270030
rect 324412 267028 324464 267034
rect 324412 266970 324464 266976
rect 324424 264316 324452 266970
rect 325528 264330 325556 271254
rect 325712 269142 325740 277766
rect 326436 275460 326488 275466
rect 326436 275402 326488 275408
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275402
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327460 266898 327488 277766
rect 327920 277766 328302 277794
rect 328472 277766 329498 277794
rect 329852 277766 330694 277794
rect 331232 277766 331890 277794
rect 332612 277766 333086 277794
rect 327920 269278 327948 277766
rect 328472 270230 328500 277766
rect 329472 275324 329524 275330
rect 329472 275266 329524 275272
rect 328460 270224 328512 270230
rect 328460 270166 328512 270172
rect 327908 269272 327960 269278
rect 327908 269214 327960 269220
rect 327448 266892 327500 266898
rect 327448 266834 327500 266840
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 329484 266422 329512 275266
rect 329656 269680 329708 269686
rect 329656 269622 329708 269628
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 329472 266416 329524 266422
rect 329472 266358 329524 266364
rect 328564 264316 328592 266358
rect 329668 264330 329696 269622
rect 329852 268394 329880 277766
rect 331036 272672 331088 272678
rect 331036 272614 331088 272620
rect 329840 268388 329892 268394
rect 329840 268330 329892 268336
rect 330208 266688 330260 266694
rect 330208 266630 330260 266636
rect 329406 264302 329696 264330
rect 330220 264316 330248 266630
rect 331048 264316 331076 272614
rect 331232 270094 331260 277766
rect 332612 270494 332640 277766
rect 334176 271318 334204 277780
rect 335372 275466 335400 277780
rect 335924 277766 336582 277794
rect 336752 277766 337778 277794
rect 335360 275460 335412 275466
rect 335360 275402 335412 275408
rect 334624 271448 334676 271454
rect 334624 271390 334676 271396
rect 334164 271312 334216 271318
rect 334164 271254 334216 271260
rect 333888 271176 333940 271182
rect 333888 271118 333940 271124
rect 332520 270466 332640 270494
rect 331220 270088 331272 270094
rect 331220 270030 331272 270036
rect 331680 269952 331732 269958
rect 331680 269894 331732 269900
rect 331692 266558 331720 269894
rect 332520 267034 332548 270466
rect 333520 268524 333572 268530
rect 333520 268466 333572 268472
rect 332508 267028 332560 267034
rect 332508 266970 332560 266976
rect 331864 266824 331916 266830
rect 331864 266766 331916 266772
rect 331680 266552 331732 266558
rect 331680 266494 331732 266500
rect 331876 264316 331904 266766
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 332704 264316 332732 266358
rect 333532 264316 333560 268466
rect 333900 266422 333928 271118
rect 334348 267436 334400 267442
rect 334348 267378 334400 267384
rect 333888 266416 333940 266422
rect 333888 266358 333940 266364
rect 334360 264316 334388 267378
rect 334636 266694 334664 271390
rect 335924 269822 335952 277766
rect 336752 269958 336780 277766
rect 338960 275330 338988 277780
rect 339512 277766 340170 277794
rect 338948 275324 339000 275330
rect 338948 275266 339000 275272
rect 338948 275188 339000 275194
rect 338948 275130 339000 275136
rect 338028 272536 338080 272542
rect 338028 272478 338080 272484
rect 336740 269952 336792 269958
rect 336740 269894 336792 269900
rect 335912 269816 335964 269822
rect 335912 269758 335964 269764
rect 336832 269816 336884 269822
rect 336832 269758 336884 269764
rect 335636 269408 335688 269414
rect 335636 269350 335688 269356
rect 335176 268388 335228 268394
rect 335176 268330 335228 268336
rect 334624 266688 334676 266694
rect 334624 266630 334676 266636
rect 335188 264316 335216 268330
rect 335648 266830 335676 269350
rect 336004 267164 336056 267170
rect 336004 267106 336056 267112
rect 335636 266824 335688 266830
rect 335636 266766 335688 266772
rect 336016 264316 336044 267106
rect 336844 264316 336872 269758
rect 338040 264330 338068 272478
rect 338960 264330 338988 275130
rect 339316 270292 339368 270298
rect 339316 270234 339368 270240
rect 337686 264302 338068 264330
rect 338514 264302 338988 264330
rect 339328 264316 339356 270234
rect 339512 269686 339540 277766
rect 341352 271454 341380 277780
rect 341524 275460 341576 275466
rect 341524 275402 341576 275408
rect 341340 271448 341392 271454
rect 341340 271390 341392 271396
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 339500 269680 339552 269686
rect 339500 269622 339552 269628
rect 340616 264330 340644 271254
rect 341536 270298 341564 275402
rect 342456 272678 342484 277780
rect 343666 277766 343864 277794
rect 342904 274236 342956 274242
rect 342904 274178 342956 274184
rect 342444 272672 342496 272678
rect 342444 272614 342496 272620
rect 342168 271448 342220 271454
rect 342168 271390 342220 271396
rect 341524 270292 341576 270298
rect 341524 270234 341576 270240
rect 341800 270224 341852 270230
rect 341800 270166 341852 270172
rect 340972 266416 341024 266422
rect 340972 266358 341024 266364
rect 340170 264302 340644 264330
rect 340984 264316 341012 266358
rect 341812 264316 341840 270166
rect 342180 266422 342208 271390
rect 342916 267442 342944 274178
rect 343836 269414 343864 277766
rect 344480 277766 344862 277794
rect 345124 277766 346058 277794
rect 344480 271182 344508 277766
rect 344468 271176 344520 271182
rect 344468 271118 344520 271124
rect 344652 271176 344704 271182
rect 344652 271118 344704 271124
rect 343824 269408 343876 269414
rect 343824 269350 343876 269356
rect 342904 267436 342956 267442
rect 342904 267378 342956 267384
rect 343456 267300 343508 267306
rect 343456 267242 343508 267248
rect 342628 266892 342680 266898
rect 342628 266834 342680 266840
rect 342168 266416 342220 266422
rect 342168 266358 342220 266364
rect 342640 264316 342668 266834
rect 343468 264316 343496 267242
rect 344664 264330 344692 271118
rect 345124 268530 345152 277766
rect 347240 274242 347268 277780
rect 347792 277766 348450 277794
rect 347228 274236 347280 274242
rect 347228 274178 347280 274184
rect 346308 273964 346360 273970
rect 346308 273906 346360 273912
rect 345112 268524 345164 268530
rect 345112 268466 345164 268472
rect 345940 268524 345992 268530
rect 345940 268466 345992 268472
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 344310 264302 344692 264330
rect 345124 264316 345152 266358
rect 345952 264316 345980 268466
rect 346320 266422 346348 273906
rect 347044 273284 347096 273290
rect 347044 273226 347096 273232
rect 347056 267170 347084 273226
rect 347596 269952 347648 269958
rect 347596 269894 347648 269900
rect 347044 267164 347096 267170
rect 347044 267106 347096 267112
rect 346768 266552 346820 266558
rect 346768 266494 346820 266500
rect 346308 266416 346360 266422
rect 346308 266358 346360 266364
rect 346780 264316 346808 266494
rect 347608 264316 347636 269894
rect 347792 268394 347820 277766
rect 349632 273290 349660 277780
rect 350552 277766 350750 277794
rect 349620 273284 349672 273290
rect 349620 273226 349672 273232
rect 350264 273284 350316 273290
rect 350264 273226 350316 273232
rect 348424 270360 348476 270366
rect 348424 270302 348476 270308
rect 347780 268388 347832 268394
rect 347780 268330 347832 268336
rect 348436 264316 348464 270302
rect 350080 268388 350132 268394
rect 350080 268330 350132 268336
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 268330
rect 350276 266422 350304 273226
rect 350552 269822 350580 277766
rect 350724 275596 350776 275602
rect 350724 275538 350776 275544
rect 350736 271182 350764 275538
rect 351932 272542 351960 277780
rect 353128 275330 353156 277780
rect 354324 275466 354352 277780
rect 354312 275460 354364 275466
rect 354312 275402 354364 275408
rect 353116 275324 353168 275330
rect 353116 275266 353168 275272
rect 353944 275324 353996 275330
rect 353944 275266 353996 275272
rect 352932 272808 352984 272814
rect 352932 272750 352984 272756
rect 351920 272536 351972 272542
rect 351920 272478 351972 272484
rect 350724 271176 350776 271182
rect 350724 271118 350776 271124
rect 351828 271176 351880 271182
rect 351828 271118 351880 271124
rect 350540 269816 350592 269822
rect 350540 269758 350592 269764
rect 351644 269680 351696 269686
rect 351644 269622 351696 269628
rect 350908 267436 350960 267442
rect 350908 267378 350960 267384
rect 350264 266416 350316 266422
rect 350264 266358 350316 266364
rect 350920 264316 350948 267378
rect 351656 266558 351684 269622
rect 351644 266552 351696 266558
rect 351644 266494 351696 266500
rect 351840 265690 351868 271118
rect 351748 265662 351868 265690
rect 351748 264316 351776 265662
rect 352944 264330 352972 272750
rect 353956 267306 353984 275266
rect 355324 271720 355376 271726
rect 355324 271662 355376 271668
rect 354220 270088 354272 270094
rect 354220 270030 354272 270036
rect 353944 267300 353996 267306
rect 353944 267242 353996 267248
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 352590 264302 352972 264330
rect 353404 264316 353432 266970
rect 354232 264316 354260 270030
rect 355336 267034 355364 271662
rect 355520 271318 355548 277780
rect 356336 275324 356388 275330
rect 356336 275266 356388 275272
rect 356348 273290 356376 275266
rect 356336 273284 356388 273290
rect 356336 273226 356388 273232
rect 356520 271856 356572 271862
rect 356520 271798 356572 271804
rect 355508 271312 355560 271318
rect 355508 271254 355560 271260
rect 355876 267164 355928 267170
rect 355876 267106 355928 267112
rect 355324 267028 355376 267034
rect 355324 266970 355376 266976
rect 355048 266552 355100 266558
rect 355048 266494 355100 266500
rect 355060 264316 355088 266494
rect 355888 264316 355916 267106
rect 356532 266898 356560 271798
rect 356716 271454 356744 277780
rect 357452 277766 357926 277794
rect 356704 271448 356756 271454
rect 356704 271390 356756 271396
rect 357452 270230 357480 277766
rect 358636 272536 358688 272542
rect 358636 272478 358688 272484
rect 357440 270224 357492 270230
rect 357440 270166 357492 270172
rect 356704 269816 356756 269822
rect 356704 269758 356756 269764
rect 356520 266892 356572 266898
rect 356520 266834 356572 266840
rect 356716 264316 356744 269758
rect 358360 266756 358412 266762
rect 358360 266698 358412 266704
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 357544 264316 357572 266358
rect 358372 264316 358400 266698
rect 358648 266422 358676 272478
rect 359016 271862 359044 277780
rect 360212 275466 360240 277780
rect 361408 275602 361436 277780
rect 361396 275596 361448 275602
rect 361396 275538 361448 275544
rect 362224 275596 362276 275602
rect 362224 275538 362276 275544
rect 360200 275460 360252 275466
rect 360200 275402 360252 275408
rect 360292 274712 360344 274718
rect 360292 274654 360344 274660
rect 360108 274100 360160 274106
rect 360108 274042 360160 274048
rect 359004 271856 359056 271862
rect 359004 271798 359056 271804
rect 359740 270496 359792 270502
rect 359740 270438 359792 270444
rect 359188 266892 359240 266898
rect 359188 266834 359240 266840
rect 358636 266416 358688 266422
rect 358636 266358 358688 266364
rect 359200 264316 359228 266834
rect 359752 266558 359780 270438
rect 360120 267734 360148 274042
rect 360304 268530 360332 274654
rect 360844 271448 360896 271454
rect 360844 271390 360896 271396
rect 360292 268524 360344 268530
rect 360292 268466 360344 268472
rect 360028 267706 360148 267734
rect 359740 266552 359792 266558
rect 359740 266494 359792 266500
rect 360028 264316 360056 267706
rect 360856 266762 360884 271390
rect 361028 268524 361080 268530
rect 361028 268466 361080 268472
rect 361040 267442 361068 268466
rect 361028 267436 361080 267442
rect 361028 267378 361080 267384
rect 360844 266756 360896 266762
rect 360844 266698 360896 266704
rect 362236 266626 362264 275538
rect 362604 273970 362632 277780
rect 363052 275460 363104 275466
rect 363052 275402 363104 275408
rect 362868 274372 362920 274378
rect 362868 274314 362920 274320
rect 362592 273964 362644 273970
rect 362592 273906 362644 273912
rect 362880 267734 362908 274314
rect 363064 270366 363092 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 365732 277766 366114 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 364156 271312 364208 271318
rect 364156 271254 364208 271260
rect 363052 270360 363104 270366
rect 363052 270302 363104 270308
rect 363052 268660 363104 268666
rect 363052 268602 363104 268608
rect 363064 267734 363092 268602
rect 362788 267706 362908 267734
rect 362972 267706 363092 267734
rect 360844 266620 360896 266626
rect 360844 266562 360896 266568
rect 362224 266620 362276 266626
rect 362224 266562 362276 266568
rect 360856 264316 360884 266562
rect 362788 266490 362816 267706
rect 361672 266484 361724 266490
rect 361672 266426 361724 266432
rect 362776 266484 362828 266490
rect 362776 266426 362828 266432
rect 361684 264316 361712 266426
rect 362972 266370 363000 267706
rect 363328 267300 363380 267306
rect 363328 267242 363380 267248
rect 362880 266342 363000 266370
rect 362880 264330 362908 266342
rect 362526 264302 362908 264330
rect 363340 264316 363368 267242
rect 364168 264316 364196 271254
rect 364352 269686 364380 277766
rect 364984 270360 365036 270366
rect 364984 270302 365036 270308
rect 364340 269680 364392 269686
rect 364340 269622 364392 269628
rect 364996 264316 365024 270302
rect 365732 269958 365760 277766
rect 367296 275466 367324 277780
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 368492 275330 368520 277780
rect 369124 275460 369176 275466
rect 369124 275402 369176 275408
rect 368480 275324 368532 275330
rect 368480 275266 368532 275272
rect 367100 274712 367152 274718
rect 367100 274654 367152 274660
rect 366916 274236 366968 274242
rect 366916 274178 366968 274184
rect 365720 269952 365772 269958
rect 365720 269894 365772 269900
rect 365812 267436 365864 267442
rect 365812 267378 365864 267384
rect 365824 264316 365852 267378
rect 366928 264330 366956 274178
rect 367112 268394 367140 274654
rect 368388 272672 368440 272678
rect 368388 272614 368440 272620
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 368204 267708 368256 267714
rect 368204 267650 368256 267656
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 366956 264330
rect 367480 264316 367508 266358
rect 368216 264330 368244 267650
rect 368400 266422 368428 272614
rect 369136 267170 369164 275402
rect 369688 274718 369716 277780
rect 369872 277766 370898 277794
rect 369676 274712 369728 274718
rect 369676 274654 369728 274660
rect 369400 270224 369452 270230
rect 369400 270166 369452 270172
rect 369124 267164 369176 267170
rect 369124 267106 369176 267112
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 369412 264330 369440 270166
rect 369872 268530 369900 277766
rect 370504 275732 370556 275738
rect 370504 275674 370556 275680
rect 369860 268524 369912 268530
rect 369860 268466 369912 268472
rect 370320 268524 370372 268530
rect 370320 268466 370372 268472
rect 370332 264330 370360 268466
rect 370516 267306 370544 275674
rect 372080 271182 372108 277780
rect 373000 277766 373290 277794
rect 373000 272814 373028 277766
rect 373172 272944 373224 272950
rect 373172 272886 373224 272892
rect 372988 272808 373040 272814
rect 372988 272750 373040 272756
rect 372528 271584 372580 271590
rect 372528 271526 372580 271532
rect 372068 271176 372120 271182
rect 372068 271118 372120 271124
rect 372344 269952 372396 269958
rect 372344 269894 372396 269900
rect 370780 267572 370832 267578
rect 370780 267514 370832 267520
rect 370504 267300 370556 267306
rect 370504 267242 370556 267248
rect 368216 264302 368322 264330
rect 369150 264302 369440 264330
rect 369978 264302 370360 264330
rect 370792 264316 370820 267514
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 371620 264316 371648 266358
rect 372356 264330 372384 269894
rect 372540 266422 372568 271526
rect 373184 267734 373212 272886
rect 374380 271726 374408 277780
rect 375392 277766 375590 277794
rect 375104 275324 375156 275330
rect 375104 275266 375156 275272
rect 374368 271720 374420 271726
rect 374368 271662 374420 271668
rect 374920 268388 374972 268394
rect 374920 268330 374972 268336
rect 373092 267706 373212 267734
rect 373092 266694 373120 267706
rect 373264 267164 373316 267170
rect 373264 267106 373316 267112
rect 373080 266688 373132 266694
rect 373080 266630 373132 266636
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267106
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 268330
rect 375116 266422 375144 275266
rect 375392 270094 375420 277766
rect 376772 270502 376800 277780
rect 377968 275466 377996 277780
rect 378152 277766 379178 277794
rect 377956 275460 378008 275466
rect 377956 275402 378008 275408
rect 377772 273964 377824 273970
rect 377772 273906 377824 273912
rect 376760 270496 376812 270502
rect 376760 270438 376812 270444
rect 377588 270496 377640 270502
rect 377588 270438 377640 270444
rect 375380 270088 375432 270094
rect 375380 270030 375432 270036
rect 376576 270088 376628 270094
rect 376576 270030 376628 270036
rect 375748 267300 375800 267306
rect 375748 267242 375800 267248
rect 375104 266416 375156 266422
rect 375104 266358 375156 266364
rect 375760 264316 375788 267242
rect 376588 264316 376616 270030
rect 377600 267714 377628 270438
rect 377588 267708 377640 267714
rect 377588 267650 377640 267656
rect 377784 264330 377812 273906
rect 378152 269822 378180 277766
rect 380360 272542 380388 277780
rect 380532 272808 380584 272814
rect 380532 272750 380584 272756
rect 380348 272536 380400 272542
rect 380348 272478 380400 272484
rect 379428 271176 379480 271182
rect 379428 271118 379480 271124
rect 378140 269816 378192 269822
rect 378140 269758 378192 269764
rect 378232 267028 378284 267034
rect 378232 266970 378284 266976
rect 377430 264302 377812 264330
rect 378244 264316 378272 266970
rect 379440 264330 379468 271118
rect 380544 267734 380572 272750
rect 380716 272536 380768 272542
rect 380716 272478 380768 272484
rect 380360 267706 380572 267734
rect 380360 264330 380388 267706
rect 379086 264302 379468 264330
rect 379914 264302 380388 264330
rect 380728 264316 380756 272478
rect 381556 271454 381584 277780
rect 382004 275460 382056 275466
rect 382004 275402 382056 275408
rect 381544 271448 381596 271454
rect 381544 271390 381596 271396
rect 381544 271040 381596 271046
rect 381544 270982 381596 270988
rect 381556 267578 381584 270982
rect 381544 267572 381596 267578
rect 381544 267514 381596 267520
rect 382016 264330 382044 275402
rect 382660 272950 382688 277780
rect 383856 274106 383884 277780
rect 385052 275602 385080 277780
rect 385040 275596 385092 275602
rect 385040 275538 385092 275544
rect 386052 274712 386104 274718
rect 386052 274654 386104 274660
rect 383844 274100 383896 274106
rect 383844 274042 383896 274048
rect 384948 274100 385000 274106
rect 384948 274042 385000 274048
rect 382924 273080 382976 273086
rect 382924 273022 382976 273028
rect 382648 272944 382700 272950
rect 382648 272886 382700 272892
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 382936 267442 382964 273022
rect 384028 269680 384080 269686
rect 384028 269622 384080 269628
rect 383200 267572 383252 267578
rect 383200 267514 383252 267520
rect 382924 267436 382976 267442
rect 382924 267378 382976 267384
rect 383212 264316 383240 267514
rect 384040 264316 384068 269622
rect 384960 267734 384988 274042
rect 386064 271318 386092 274654
rect 386248 274378 386276 277780
rect 386432 277766 387458 277794
rect 386236 274372 386288 274378
rect 386236 274314 386288 274320
rect 386052 271312 386104 271318
rect 386052 271254 386104 271260
rect 385684 269816 385736 269822
rect 385684 269758 385736 269764
rect 384868 267706 384988 267734
rect 384868 264316 384896 267706
rect 385696 264316 385724 269758
rect 386432 268666 386460 277766
rect 388640 275738 388668 277780
rect 389180 276004 389232 276010
rect 389180 275946 389232 275952
rect 388628 275732 388680 275738
rect 388628 275674 388680 275680
rect 388168 275596 388220 275602
rect 388168 275538 388220 275544
rect 387708 271720 387760 271726
rect 387708 271662 387760 271668
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386420 268660 386472 268666
rect 386420 268602 386472 268608
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271662
rect 388180 269686 388208 275538
rect 389192 274242 389220 275946
rect 389744 274718 389772 277780
rect 390572 277766 390954 277794
rect 389732 274712 389784 274718
rect 389732 274654 389784 274660
rect 389180 274236 389232 274242
rect 389180 274178 389232 274184
rect 390284 274236 390336 274242
rect 390284 274178 390336 274184
rect 388628 272944 388680 272950
rect 388628 272886 388680 272892
rect 388640 272678 388668 272886
rect 388628 272672 388680 272678
rect 388628 272614 388680 272620
rect 389088 270904 389140 270910
rect 389088 270846 389140 270852
rect 388168 269680 388220 269686
rect 388168 269622 388220 269628
rect 389100 267734 389128 270846
rect 388168 267708 388220 267714
rect 388168 267650 388220 267656
rect 389008 267706 389128 267734
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 267650
rect 389008 264316 389036 267706
rect 390296 264330 390324 274178
rect 390572 270366 390600 277766
rect 392136 273086 392164 277780
rect 393332 276010 393360 277780
rect 393320 276004 393372 276010
rect 393320 275946 393372 275952
rect 393596 275868 393648 275874
rect 393596 275810 393648 275816
rect 392584 274508 392636 274514
rect 392584 274450 392636 274456
rect 392124 273080 392176 273086
rect 392124 273022 392176 273028
rect 391848 272944 391900 272950
rect 391848 272886 391900 272892
rect 390560 270360 390612 270366
rect 390560 270302 390612 270308
rect 390652 267436 390704 267442
rect 390652 267378 390704 267384
rect 389850 264302 390324 264330
rect 390664 264316 390692 267378
rect 391860 264330 391888 272886
rect 392308 270360 392360 270366
rect 392308 270302 392360 270308
rect 391506 264302 391888 264330
rect 392320 264316 392348 270302
rect 392596 267170 392624 274450
rect 393608 272678 393636 275810
rect 394528 272814 394556 277780
rect 394712 277766 395738 277794
rect 396092 277766 396934 277794
rect 397472 277766 398038 277794
rect 394516 272808 394568 272814
rect 394516 272750 394568 272756
rect 393596 272672 393648 272678
rect 393596 272614 393648 272620
rect 393964 272672 394016 272678
rect 393964 272614 394016 272620
rect 393976 267306 394004 272614
rect 394332 271856 394384 271862
rect 394332 271798 394384 271804
rect 393964 267300 394016 267306
rect 393964 267242 394016 267248
rect 392584 267164 392636 267170
rect 392584 267106 392636 267112
rect 393136 266892 393188 266898
rect 393136 266834 393188 266840
rect 393148 264316 393176 266834
rect 394344 264330 394372 271798
rect 394712 270502 394740 277766
rect 395896 274372 395948 274378
rect 395896 274314 395948 274320
rect 394700 270496 394752 270502
rect 394700 270438 394752 270444
rect 394700 269680 394752 269686
rect 394700 269622 394752 269628
rect 394712 267578 394740 269622
rect 394700 267572 394752 267578
rect 394700 267514 394752 267520
rect 394792 266552 394844 266558
rect 394792 266494 394844 266500
rect 393990 264302 394372 264330
rect 394804 264316 394832 266494
rect 395908 264330 395936 274314
rect 396092 270230 396120 277766
rect 397276 272808 397328 272814
rect 397276 272750 397328 272756
rect 397092 270496 397144 270502
rect 397092 270438 397144 270444
rect 396080 270224 396132 270230
rect 396080 270166 396132 270172
rect 397104 267714 397132 270438
rect 397092 267708 397144 267714
rect 397092 267650 397144 267656
rect 397092 267572 397144 267578
rect 397092 267514 397144 267520
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 395646 264302 395936 264330
rect 396460 264316 396488 266358
rect 397104 264330 397132 267514
rect 397288 266422 397316 272750
rect 397472 268530 397500 277766
rect 397920 271448 397972 271454
rect 397920 271390 397972 271396
rect 397460 268524 397512 268530
rect 397460 268466 397512 268472
rect 397932 266558 397960 271390
rect 399220 271046 399248 277780
rect 400416 271590 400444 277780
rect 401626 277766 401824 277794
rect 400588 276004 400640 276010
rect 400588 275946 400640 275952
rect 400404 271584 400456 271590
rect 400404 271526 400456 271532
rect 400128 271312 400180 271318
rect 400128 271254 400180 271260
rect 399208 271040 399260 271046
rect 399208 270982 399260 270988
rect 398104 267708 398156 267714
rect 398104 267650 398156 267656
rect 397920 266552 397972 266558
rect 397920 266494 397972 266500
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 267650
rect 399760 267300 399812 267306
rect 399760 267242 399812 267248
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 267242
rect 400140 266422 400168 271254
rect 400600 268938 400628 275946
rect 401324 271040 401376 271046
rect 401324 270982 401376 270988
rect 400588 268932 400640 268938
rect 400588 268874 400640 268880
rect 400588 268660 400640 268666
rect 400588 268602 400640 268608
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 268602
rect 401336 264330 401364 270982
rect 401796 269958 401824 277766
rect 402808 274514 402836 277780
rect 404004 275330 404032 277780
rect 404556 277766 405214 277794
rect 403992 275324 404044 275330
rect 403992 275266 404044 275272
rect 404268 274848 404320 274854
rect 404268 274790 404320 274796
rect 402796 274508 402848 274514
rect 402796 274450 402848 274456
rect 403992 273080 404044 273086
rect 403992 273022 404044 273028
rect 403072 270224 403124 270230
rect 403072 270166 403124 270172
rect 401784 269952 401836 269958
rect 401784 269894 401836 269900
rect 401600 269544 401652 269550
rect 401600 269486 401652 269492
rect 401612 266898 401640 269486
rect 402244 268524 402296 268530
rect 402244 268466 402296 268472
rect 401600 266892 401652 266898
rect 401600 266834 401652 266840
rect 401336 264302 401442 264330
rect 402256 264316 402284 268466
rect 403084 264316 403112 270166
rect 404004 267734 404032 273022
rect 404280 270094 404308 274790
rect 404268 270088 404320 270094
rect 404268 270030 404320 270036
rect 404360 269408 404412 269414
rect 404360 269350 404412 269356
rect 403912 267706 404032 267734
rect 403912 264316 403940 267706
rect 404372 267442 404400 269350
rect 404556 268394 404584 277766
rect 406304 272678 406332 277780
rect 407500 274854 407528 277780
rect 407488 274848 407540 274854
rect 407488 274790 407540 274796
rect 407120 274712 407172 274718
rect 407120 274654 407172 274660
rect 406844 274508 406896 274514
rect 406844 274450 406896 274456
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 404544 268388 404596 268394
rect 404544 268330 404596 268336
rect 404360 267436 404412 267442
rect 404360 267378 404412 267384
rect 404728 267164 404780 267170
rect 404728 267106 404780 267112
rect 404740 264316 404768 267106
rect 405556 266892 405608 266898
rect 405556 266834 405608 266840
rect 405568 264316 405596 266834
rect 406856 264330 406884 274450
rect 407132 271182 407160 274654
rect 408696 273970 408724 277780
rect 408684 273964 408736 273970
rect 408684 273906 408736 273912
rect 409892 273290 409920 277780
rect 410064 275732 410116 275738
rect 410064 275674 410116 275680
rect 409144 273284 409196 273290
rect 409144 273226 409196 273232
rect 409880 273284 409932 273290
rect 409880 273226 409932 273232
rect 408408 272672 408460 272678
rect 408408 272614 408460 272620
rect 407120 271176 407172 271182
rect 407120 271118 407172 271124
rect 407212 268388 407264 268394
rect 407212 268330 407264 268336
rect 406410 264302 406884 264330
rect 407224 264316 407252 268330
rect 408420 264330 408448 272614
rect 409156 267034 409184 273226
rect 410076 272950 410104 275674
rect 411088 274718 411116 277780
rect 412284 275874 412312 277780
rect 412272 275868 412324 275874
rect 412272 275810 412324 275816
rect 411260 275324 411312 275330
rect 411260 275266 411312 275272
rect 411076 274712 411128 274718
rect 411076 274654 411128 274660
rect 410064 272944 410116 272950
rect 410064 272886 410116 272892
rect 411272 271946 411300 275266
rect 412456 272944 412508 272950
rect 412456 272886 412508 272892
rect 410904 271918 411300 271946
rect 409788 271584 409840 271590
rect 409788 271526 409840 271532
rect 409604 267436 409656 267442
rect 409604 267378 409656 267384
rect 409144 267028 409196 267034
rect 409144 266970 409196 266976
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408066 264302 408448 264330
rect 408880 264316 408908 266358
rect 409616 264330 409644 267378
rect 409800 266422 409828 271526
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410904 264330 410932 271918
rect 412180 266756 412232 266762
rect 412180 266698 412232 266704
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 409616 264302 409722 264330
rect 410550 264302 410932 264330
rect 411364 264316 411392 266358
rect 412192 264316 412220 266698
rect 412468 266422 412496 272886
rect 413388 272542 413416 277780
rect 414584 275466 414612 277780
rect 415780 276010 415808 277780
rect 416792 277766 416990 277794
rect 415768 276004 415820 276010
rect 415768 275946 415820 275952
rect 415308 275868 415360 275874
rect 415308 275810 415360 275816
rect 414572 275460 414624 275466
rect 414572 275402 414624 275408
rect 413928 273964 413980 273970
rect 413928 273906 413980 273912
rect 413376 272536 413428 272542
rect 413376 272478 413428 272484
rect 413008 269952 413060 269958
rect 413008 269894 413060 269900
rect 412456 266416 412508 266422
rect 412456 266358 412508 266364
rect 413020 264316 413048 269894
rect 413940 267734 413968 273906
rect 415124 272536 415176 272542
rect 415124 272478 415176 272484
rect 413848 267706 413968 267734
rect 413848 264316 413876 267706
rect 415136 264330 415164 272478
rect 415320 270910 415348 275810
rect 416412 275460 416464 275466
rect 416412 275402 416464 275408
rect 415308 270904 415360 270910
rect 415308 270846 415360 270852
rect 416424 266422 416452 275402
rect 416596 271176 416648 271182
rect 416596 271118 416648 271124
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415164 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 271118
rect 416792 269686 416820 277766
rect 418172 275602 418200 277780
rect 418160 275596 418212 275602
rect 418160 275538 418212 275544
rect 418344 275596 418396 275602
rect 418344 275538 418396 275544
rect 418356 272814 418384 275538
rect 419368 274106 419396 277780
rect 419552 277766 420578 277794
rect 421392 277766 421682 277794
rect 422312 277766 422878 277794
rect 423692 277766 424074 277794
rect 419356 274100 419408 274106
rect 419356 274042 419408 274048
rect 419172 273216 419224 273222
rect 419172 273158 419224 273164
rect 418344 272808 418396 272814
rect 418344 272750 418396 272756
rect 417148 270088 417200 270094
rect 417148 270030 417200 270036
rect 416780 269680 416832 269686
rect 416780 269622 416832 269628
rect 416346 264302 416636 264330
rect 417160 264316 417188 270030
rect 418988 268932 419040 268938
rect 418988 268874 419040 268880
rect 419000 267306 419028 268874
rect 418988 267300 419040 267306
rect 418988 267242 419040 267248
rect 417976 266756 418028 266762
rect 417976 266698 418028 266704
rect 417988 264316 418016 266698
rect 419184 264330 419212 273158
rect 419552 269822 419580 277766
rect 420920 275188 420972 275194
rect 420920 275130 420972 275136
rect 420932 274378 420960 275130
rect 420920 274372 420972 274378
rect 420920 274314 420972 274320
rect 421392 271726 421420 277766
rect 421564 274100 421616 274106
rect 421564 274042 421616 274048
rect 421380 271720 421432 271726
rect 421380 271662 421432 271668
rect 419540 269816 419592 269822
rect 419540 269758 419592 269764
rect 420000 269816 420052 269822
rect 420000 269758 420052 269764
rect 420012 264330 420040 269758
rect 420460 268116 420512 268122
rect 420460 268058 420512 268064
rect 418830 264302 419212 264330
rect 419658 264302 420040 264330
rect 420472 264316 420500 268058
rect 421288 267300 421340 267306
rect 421288 267242 421340 267248
rect 421300 264316 421328 267242
rect 421576 266626 421604 274042
rect 421748 271720 421800 271726
rect 421748 271662 421800 271668
rect 421760 267714 421788 271662
rect 422312 269074 422340 277766
rect 423692 270502 423720 277766
rect 425256 275874 425284 277780
rect 425244 275868 425296 275874
rect 425244 275810 425296 275816
rect 426256 274848 426308 274854
rect 426256 274790 426308 274796
rect 424968 274644 425020 274650
rect 424968 274586 425020 274592
rect 423680 270496 423732 270502
rect 423680 270438 423732 270444
rect 424600 270496 424652 270502
rect 424600 270438 424652 270444
rect 422300 269068 422352 269074
rect 422300 269010 422352 269016
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 421748 267708 421800 267714
rect 421748 267650 421800 267656
rect 422312 267578 422340 268738
rect 422300 267572 422352 267578
rect 422300 267514 422352 267520
rect 422116 267028 422168 267034
rect 422116 266970 422168 266976
rect 421564 266620 421616 266626
rect 421564 266562 421616 266568
rect 422128 264316 422156 266970
rect 422944 266620 422996 266626
rect 422944 266562 422996 266568
rect 422956 264316 422984 266562
rect 423772 266416 423824 266422
rect 423772 266358 423824 266364
rect 423784 264316 423812 266358
rect 424612 264316 424640 270438
rect 424980 266422 425008 274586
rect 426072 272808 426124 272814
rect 426072 272750 426124 272756
rect 425704 271040 425756 271046
rect 425704 270982 425756 270988
rect 425716 266898 425744 270982
rect 425704 266892 425756 266898
rect 425704 266834 425756 266840
rect 424968 266416 425020 266422
rect 424968 266358 425020 266364
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426084 264330 426112 272750
rect 426268 271862 426296 274790
rect 426452 274242 426480 277780
rect 426636 277766 427662 277794
rect 426440 274236 426492 274242
rect 426440 274178 426492 274184
rect 426256 271856 426308 271862
rect 426256 271798 426308 271804
rect 426636 269414 426664 277766
rect 427820 276004 427872 276010
rect 427820 275946 427872 275952
rect 426900 273828 426952 273834
rect 426900 273770 426952 273776
rect 426624 269408 426676 269414
rect 426624 269350 426676 269356
rect 426912 266422 426940 273770
rect 427084 271856 427136 271862
rect 427084 271798 427136 271804
rect 427096 271454 427124 271798
rect 427084 271448 427136 271454
rect 427084 271390 427136 271396
rect 427268 271448 427320 271454
rect 427268 271390 427320 271396
rect 427280 271046 427308 271390
rect 427268 271040 427320 271046
rect 427268 270982 427320 270988
rect 427832 270910 427860 275946
rect 428844 275738 428872 277780
rect 429396 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275732 428884 275738
rect 428832 275674 428884 275680
rect 429200 275732 429252 275738
rect 429200 275674 429252 275680
rect 429016 273556 429068 273562
rect 429016 273498 429068 273504
rect 427820 270904 427872 270910
rect 427820 270846 427872 270852
rect 428464 270632 428516 270638
rect 428464 270574 428516 270580
rect 427360 269680 427412 269686
rect 427360 269622 427412 269628
rect 426900 266416 426952 266422
rect 426900 266358 426952 266364
rect 427372 264330 427400 269622
rect 428476 266898 428504 270574
rect 428464 266892 428516 266898
rect 428464 266834 428516 266840
rect 427912 266756 427964 266762
rect 427912 266698 427964 266704
rect 426084 264302 426282 264330
rect 427110 264302 427400 264330
rect 427924 264316 427952 266698
rect 429028 264330 429056 273498
rect 429212 273086 429240 275674
rect 429200 273080 429252 273086
rect 429200 273022 429252 273028
rect 429396 270366 429424 277766
rect 429384 270360 429436 270366
rect 429384 270302 429436 270308
rect 429568 270360 429620 270366
rect 429568 270302 429620 270308
rect 428766 264302 429056 264330
rect 429580 264316 429608 270302
rect 430592 269550 430620 277766
rect 432340 274854 432368 277780
rect 432972 275868 433024 275874
rect 432972 275810 433024 275816
rect 432328 274848 432380 274854
rect 432328 274790 432380 274796
rect 431684 271040 431736 271046
rect 431684 270982 431736 270988
rect 430580 269544 430632 269550
rect 430580 269486 430632 269492
rect 430396 267708 430448 267714
rect 430396 267650 430448 267656
rect 430408 264316 430436 267650
rect 431696 264330 431724 270982
rect 431960 267844 432012 267850
rect 431960 267786 432012 267792
rect 431972 267170 432000 267786
rect 432984 267734 433012 275810
rect 433536 271862 433564 277780
rect 434732 275194 434760 277780
rect 435928 275602 435956 277780
rect 436112 277766 437046 277794
rect 435916 275596 435968 275602
rect 435916 275538 435968 275544
rect 434720 275188 434772 275194
rect 434720 275130 434772 275136
rect 435640 274780 435692 274786
rect 435640 274722 435692 274728
rect 434628 273080 434680 273086
rect 434628 273022 434680 273028
rect 433524 271856 433576 271862
rect 433524 271798 433576 271804
rect 433156 270768 433208 270774
rect 433156 270710 433208 270716
rect 432892 267706 433012 267734
rect 431960 267164 432012 267170
rect 431960 267106 432012 267112
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267706
rect 433168 266422 433196 270710
rect 434444 269136 434496 269142
rect 434444 269078 434496 269084
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433708 266416 433760 266422
rect 433708 266358 433760 266364
rect 433720 264316 433748 266358
rect 434456 264330 434484 269078
rect 434640 266422 434668 273022
rect 435652 271318 435680 274722
rect 435640 271312 435692 271318
rect 435640 271254 435692 271260
rect 435364 270904 435416 270910
rect 435364 270846 435416 270852
rect 435376 267442 435404 270846
rect 436112 268802 436140 277766
rect 437480 275188 437532 275194
rect 437480 275130 437532 275136
rect 437492 274514 437520 275130
rect 437480 274508 437532 274514
rect 437480 274450 437532 274456
rect 438228 271726 438256 277780
rect 439424 274786 439452 277780
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439412 274780 439464 274786
rect 439412 274722 439464 274728
rect 438768 274236 438820 274242
rect 438768 274178 438820 274184
rect 438216 271720 438268 271726
rect 438216 271662 438268 271668
rect 436928 271448 436980 271454
rect 436928 271390 436980 271396
rect 436940 270910 436968 271390
rect 436928 270904 436980 270910
rect 436928 270846 436980 270852
rect 436100 268796 436152 268802
rect 436100 268738 436152 268744
rect 436192 268252 436244 268258
rect 436192 268194 436244 268200
rect 435364 267436 435416 267442
rect 435364 267378 435416 267384
rect 435180 266892 435232 266898
rect 435180 266834 435232 266840
rect 435192 266626 435220 266834
rect 435180 266620 435232 266626
rect 435180 266562 435232 266568
rect 435364 266620 435416 266626
rect 435364 266562 435416 266568
rect 434628 266416 434680 266422
rect 434628 266358 434680 266364
rect 434456 264302 434562 264330
rect 435376 264316 435404 266562
rect 436204 264316 436232 268194
rect 437848 267980 437900 267986
rect 437848 267922 437900 267928
rect 437020 266416 437072 266422
rect 437020 266358 437072 266364
rect 437032 264316 437060 266358
rect 437860 264316 437888 267922
rect 438780 267734 438808 274178
rect 439320 272400 439372 272406
rect 439320 272342 439372 272348
rect 438688 267706 438808 267734
rect 438688 264316 438716 267706
rect 439332 266898 439360 272342
rect 440252 268938 440280 277766
rect 440884 274508 440936 274514
rect 440884 274450 440936 274456
rect 440240 268932 440292 268938
rect 440240 268874 440292 268880
rect 440332 267436 440384 267442
rect 440332 267378 440384 267384
rect 439504 267164 439556 267170
rect 439504 267106 439556 267112
rect 439320 266892 439372 266898
rect 439320 266834 439372 266840
rect 439516 264316 439544 267106
rect 440344 264316 440372 267378
rect 440896 266422 440924 274450
rect 441160 268796 441212 268802
rect 441160 268738 441212 268744
rect 440884 266416 440936 266422
rect 440884 266358 440936 266364
rect 441172 264316 441200 268738
rect 441632 268666 441660 277766
rect 443012 276010 443040 277780
rect 443288 277766 444222 277794
rect 444392 277766 445326 277794
rect 443000 276004 443052 276010
rect 443000 275946 443052 275952
rect 442908 271720 442960 271726
rect 442908 271662 442960 271668
rect 441620 268660 441672 268666
rect 441620 268602 441672 268608
rect 442724 268660 442776 268666
rect 442724 268602 442776 268608
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 268602
rect 442920 266422 442948 271662
rect 443288 268530 443316 277766
rect 443736 276004 443788 276010
rect 443736 275946 443788 275952
rect 443748 271590 443776 275946
rect 443736 271584 443788 271590
rect 443736 271526 443788 271532
rect 444392 270230 444420 277766
rect 446508 275738 446536 277780
rect 447152 277766 447718 277794
rect 446496 275732 446548 275738
rect 446496 275674 446548 275680
rect 445760 275596 445812 275602
rect 445760 275538 445812 275544
rect 445024 270904 445076 270910
rect 445024 270846 445076 270852
rect 444380 270224 444432 270230
rect 444380 270166 444432 270172
rect 443644 268932 443696 268938
rect 443644 268874 443696 268880
rect 443276 268524 443328 268530
rect 443276 268466 443328 268472
rect 443460 267572 443512 267578
rect 443460 267514 443512 267520
rect 443472 267034 443500 267514
rect 443460 267028 443512 267034
rect 443460 266970 443512 266976
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 442736 264302 442842 264330
rect 443656 264316 443684 268874
rect 445036 267170 445064 270846
rect 445772 268666 445800 275538
rect 446956 270224 447008 270230
rect 446956 270166 447008 270172
rect 445760 268660 445812 268666
rect 445760 268602 445812 268608
rect 446588 268660 446640 268666
rect 446588 268602 446640 268608
rect 445024 267164 445076 267170
rect 445024 267106 445076 267112
rect 445300 267164 445352 267170
rect 445300 267106 445352 267112
rect 444472 266552 444524 266558
rect 444472 266494 444524 266500
rect 444484 264316 444512 266494
rect 445312 264316 445340 267106
rect 446600 264330 446628 268602
rect 446154 264302 446628 264330
rect 446968 264316 446996 270166
rect 447152 267850 447180 277766
rect 447784 271856 447836 271862
rect 447784 271798 447836 271804
rect 447140 267844 447192 267850
rect 447140 267786 447192 267792
rect 447796 266558 447824 271798
rect 448900 271318 448928 277780
rect 449164 275596 449216 275602
rect 449164 275538 449216 275544
rect 448888 271312 448940 271318
rect 448888 271254 448940 271260
rect 448612 268524 448664 268530
rect 448612 268466 448664 268472
rect 447784 266552 447836 266558
rect 447784 266494 447836 266500
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 447796 264316 447824 266358
rect 448624 264316 448652 268466
rect 449176 266422 449204 275538
rect 450096 275194 450124 277780
rect 451306 277766 451504 277794
rect 450084 275188 450136 275194
rect 450084 275130 450136 275136
rect 449900 275052 449952 275058
rect 449900 274994 449952 275000
rect 449912 273970 449940 274994
rect 449900 273964 449952 273970
rect 449900 273906 449952 273912
rect 451096 273964 451148 273970
rect 451096 273906 451148 273912
rect 449900 269544 449952 269550
rect 449900 269486 449952 269492
rect 449912 267578 449940 269486
rect 449900 267572 449952 267578
rect 449900 267514 449952 267520
rect 450084 267572 450136 267578
rect 450084 267514 450136 267520
rect 450096 267170 450124 267514
rect 450084 267164 450136 267170
rect 450084 267106 450136 267112
rect 450268 267164 450320 267170
rect 450268 267106 450320 267112
rect 449440 266756 449492 266762
rect 449440 266698 449492 266704
rect 449164 266416 449216 266422
rect 449164 266358 449216 266364
rect 449452 264316 449480 266698
rect 450280 264316 450308 267106
rect 451108 264316 451136 273906
rect 451476 268394 451504 277766
rect 452488 272678 452516 277780
rect 453592 276010 453620 277780
rect 453580 276004 453632 276010
rect 453580 275946 453632 275952
rect 453948 274780 454000 274786
rect 453948 274722 454000 274728
rect 453960 272950 453988 274722
rect 453948 272944 454000 272950
rect 453948 272886 454000 272892
rect 452476 272672 452528 272678
rect 452476 272614 452528 272620
rect 453856 272672 453908 272678
rect 453856 272614 453908 272620
rect 451924 272264 451976 272270
rect 451924 272206 451976 272212
rect 451464 268388 451516 268394
rect 451464 268330 451516 268336
rect 451936 267034 451964 272206
rect 453304 271584 453356 271590
rect 453304 271526 453356 271532
rect 451924 267028 451976 267034
rect 451924 266970 451976 266976
rect 452752 266688 452804 266694
rect 452752 266630 452804 266636
rect 451924 266416 451976 266422
rect 451924 266358 451976 266364
rect 451936 264316 451964 266358
rect 452764 264316 452792 266630
rect 453316 266558 453344 271526
rect 453304 266552 453356 266558
rect 453304 266494 453356 266500
rect 453868 264330 453896 272614
rect 454788 271454 454816 277780
rect 455984 275330 456012 277780
rect 456984 276004 457036 276010
rect 456984 275946 457036 275952
rect 455972 275324 456024 275330
rect 455972 275266 456024 275272
rect 456156 275324 456208 275330
rect 456156 275266 456208 275272
rect 454776 271448 454828 271454
rect 454776 271390 454828 271396
rect 454684 271312 454736 271318
rect 454684 271254 454736 271260
rect 454408 266552 454460 266558
rect 454408 266494 454460 266500
rect 453606 264302 453896 264330
rect 454420 264316 454448 266494
rect 454696 266422 454724 271254
rect 455236 267028 455288 267034
rect 455236 266970 455288 266976
rect 454684 266416 454736 266422
rect 454684 266358 454736 266364
rect 455248 264316 455276 266970
rect 456168 266694 456196 275266
rect 456800 275188 456852 275194
rect 456800 275130 456852 275136
rect 456812 273222 456840 275130
rect 456800 273216 456852 273222
rect 456800 273158 456852 273164
rect 456996 270774 457024 275946
rect 457180 274786 457208 277780
rect 457168 274780 457220 274786
rect 457168 274722 457220 274728
rect 458376 274106 458404 277780
rect 458364 274100 458416 274106
rect 458364 274042 458416 274048
rect 459376 274100 459428 274106
rect 459376 274042 459428 274048
rect 458088 272944 458140 272950
rect 458088 272886 458140 272892
rect 457444 271448 457496 271454
rect 457444 271390 457496 271396
rect 456984 270768 457036 270774
rect 456984 270710 457036 270716
rect 456432 266756 456484 266762
rect 456432 266698 456484 266704
rect 456156 266688 456208 266694
rect 456156 266630 456208 266636
rect 456444 264330 456472 266698
rect 457456 266558 457484 271390
rect 457720 269408 457772 269414
rect 457720 269350 457772 269356
rect 457444 266552 457496 266558
rect 457444 266494 457496 266500
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456090 264302 456472 264330
rect 456904 264316 456932 266358
rect 457732 264316 457760 269350
rect 458100 266422 458128 272886
rect 459192 266620 459244 266626
rect 459192 266562 459244 266568
rect 458088 266416 458140 266422
rect 458088 266358 458140 266364
rect 458548 266416 458600 266422
rect 458548 266358 458600 266364
rect 458560 264316 458588 266358
rect 459204 264330 459232 266562
rect 459388 266422 459416 274042
rect 459572 269958 459600 277780
rect 460676 275058 460704 277780
rect 460664 275052 460716 275058
rect 460664 274994 460716 275000
rect 460020 273692 460072 273698
rect 460020 273634 460072 273640
rect 459560 269952 459612 269958
rect 459560 269894 459612 269900
rect 460032 267714 460060 273634
rect 461872 272542 461900 277780
rect 463068 275466 463096 277780
rect 463988 277766 464278 277794
rect 465092 277766 465474 277794
rect 463056 275460 463108 275466
rect 463056 275402 463108 275408
rect 463516 273216 463568 273222
rect 463516 273158 463568 273164
rect 461860 272536 461912 272542
rect 461860 272478 461912 272484
rect 463332 272536 463384 272542
rect 463332 272478 463384 272484
rect 461860 269952 461912 269958
rect 461860 269894 461912 269900
rect 461032 268388 461084 268394
rect 461032 268330 461084 268336
rect 460020 267708 460072 267714
rect 460020 267650 460072 267656
rect 460204 267708 460256 267714
rect 460204 267650 460256 267656
rect 460216 267034 460244 267650
rect 460204 267028 460256 267034
rect 460204 266970 460256 266976
rect 460204 266484 460256 266490
rect 460204 266426 460256 266432
rect 459376 266416 459428 266422
rect 459376 266358 459428 266364
rect 459204 264302 459402 264330
rect 460216 264316 460244 266426
rect 461044 264316 461072 268330
rect 461872 264316 461900 269894
rect 462320 267028 462372 267034
rect 462320 266970 462372 266976
rect 462332 266762 462360 266970
rect 462320 266756 462372 266762
rect 462320 266698 462372 266704
rect 462688 266620 462740 266626
rect 462688 266562 462740 266568
rect 462700 264316 462728 266562
rect 463344 264330 463372 272478
rect 463528 266626 463556 273158
rect 463988 271182 464016 277766
rect 464344 274780 464396 274786
rect 464344 274722 464396 274728
rect 463976 271176 464028 271182
rect 463976 271118 464028 271124
rect 464356 267306 464384 274722
rect 464528 271176 464580 271182
rect 464528 271118 464580 271124
rect 464344 267300 464396 267306
rect 464344 267242 464396 267248
rect 464540 266762 464568 271118
rect 465092 270094 465120 277766
rect 465724 270768 465776 270774
rect 465724 270710 465776 270716
rect 465080 270088 465132 270094
rect 465080 270030 465132 270036
rect 465540 267708 465592 267714
rect 465540 267650 465592 267656
rect 465172 267300 465224 267306
rect 465172 267242 465224 267248
rect 464988 267028 465040 267034
rect 464988 266970 465040 266976
rect 465000 266762 465028 266970
rect 464528 266756 464580 266762
rect 464528 266698 464580 266704
rect 464988 266756 465040 266762
rect 464988 266698 465040 266704
rect 463516 266620 463568 266626
rect 463516 266562 463568 266568
rect 464344 266620 464396 266626
rect 464344 266562 464396 266568
rect 463344 264302 463542 264330
rect 464356 264316 464384 266562
rect 465184 264316 465212 267242
rect 465552 267034 465580 267650
rect 465540 267028 465592 267034
rect 465540 266970 465592 266976
rect 465736 266626 465764 270710
rect 466656 270638 466684 277780
rect 467656 275460 467708 275466
rect 467656 275402 467708 275408
rect 466644 270632 466696 270638
rect 466644 270574 466696 270580
rect 466000 270088 466052 270094
rect 466000 270030 466052 270036
rect 465724 266620 465776 266626
rect 465724 266562 465776 266568
rect 466012 264316 466040 270030
rect 466828 267708 466880 267714
rect 466828 267650 466880 267656
rect 466840 264316 466868 267650
rect 467668 264316 467696 275402
rect 467852 275194 467880 277780
rect 468036 277766 468970 277794
rect 469232 277766 470166 277794
rect 467840 275188 467892 275194
rect 467840 275130 467892 275136
rect 468036 269822 468064 277766
rect 468208 275188 468260 275194
rect 468208 275130 468260 275136
rect 468024 269816 468076 269822
rect 468024 269758 468076 269764
rect 468220 267986 468248 275130
rect 468760 269272 468812 269278
rect 468760 269214 468812 269220
rect 468208 267980 468260 267986
rect 468208 267922 468260 267928
rect 468772 264330 468800 269214
rect 469232 268274 469260 277766
rect 471348 274786 471376 277780
rect 471992 277766 472558 277794
rect 471796 274916 471848 274922
rect 471796 274858 471848 274864
rect 471336 274780 471388 274786
rect 471336 274722 471388 274728
rect 471244 274372 471296 274378
rect 471244 274314 471296 274320
rect 470968 269816 471020 269822
rect 470968 269758 471020 269764
rect 469048 268246 469260 268274
rect 469048 268122 469076 268246
rect 469036 268116 469088 268122
rect 469036 268058 469088 268064
rect 469220 268116 469272 268122
rect 469220 268058 469272 268064
rect 469232 266762 469260 268058
rect 470140 267708 470192 267714
rect 470140 267650 470192 267656
rect 469220 266756 469272 266762
rect 469220 266698 469272 266704
rect 469312 266620 469364 266626
rect 469312 266562 469364 266568
rect 468510 264302 468800 264330
rect 469324 264316 469352 266562
rect 470152 264316 470180 267650
rect 470980 264316 471008 269758
rect 471256 266898 471284 274314
rect 471808 269414 471836 274858
rect 471992 269550 472020 277766
rect 473740 272406 473768 277780
rect 474936 274650 474964 277780
rect 476146 277766 476344 277794
rect 474924 274644 474976 274650
rect 474924 274586 474976 274592
rect 475384 274644 475436 274650
rect 475384 274586 475436 274592
rect 473728 272400 473780 272406
rect 473728 272342 473780 272348
rect 474648 272400 474700 272406
rect 474648 272342 474700 272348
rect 473084 272128 473136 272134
rect 473084 272070 473136 272076
rect 471980 269544 472032 269550
rect 471980 269486 472032 269492
rect 471796 269408 471848 269414
rect 471796 269350 471848 269356
rect 471244 266892 471296 266898
rect 471244 266834 471296 266840
rect 471796 266756 471848 266762
rect 471796 266698 471848 266704
rect 471808 264316 471836 266698
rect 473096 264330 473124 272070
rect 474280 269544 474332 269550
rect 474280 269486 474332 269492
rect 473452 266620 473504 266626
rect 473452 266562 473504 266568
rect 472650 264302 473124 264330
rect 473464 264316 473492 266562
rect 474292 264316 474320 269486
rect 474660 266626 474688 272342
rect 475396 266762 475424 274586
rect 476316 270502 476344 277766
rect 477236 273834 477264 277780
rect 477224 273828 477276 273834
rect 477224 273770 477276 273776
rect 478432 272814 478460 277780
rect 478892 277766 479642 277794
rect 478420 272808 478472 272814
rect 478420 272750 478472 272756
rect 478420 271992 478472 271998
rect 478420 271934 478472 271940
rect 477500 270632 477552 270638
rect 477500 270574 477552 270580
rect 476304 270496 476356 270502
rect 476304 270438 476356 270444
rect 476764 269408 476816 269414
rect 476764 269350 476816 269356
rect 475384 266756 475436 266762
rect 475384 266698 475436 266704
rect 475936 266756 475988 266762
rect 475936 266698 475988 266704
rect 474648 266620 474700 266626
rect 474648 266562 474700 266568
rect 475108 266076 475160 266082
rect 475108 266018 475160 266024
rect 475120 264316 475148 266018
rect 475948 264316 475976 266698
rect 476776 264316 476804 269350
rect 477512 266744 477540 270574
rect 477328 266716 477540 266744
rect 477328 266626 477356 266716
rect 477316 266620 477368 266626
rect 477316 266562 477368 266568
rect 477592 266620 477644 266626
rect 477592 266562 477644 266568
rect 477604 264316 477632 266562
rect 478432 264316 478460 271934
rect 478892 269686 478920 277766
rect 480824 272270 480852 277780
rect 482020 273562 482048 277780
rect 483216 277394 483244 277780
rect 483124 277366 483244 277394
rect 482928 274780 482980 274786
rect 482928 274722 482980 274728
rect 482008 273556 482060 273562
rect 482008 273498 482060 273504
rect 481364 273420 481416 273426
rect 481364 273362 481416 273368
rect 480812 272264 480864 272270
rect 480812 272206 480864 272212
rect 479248 270496 479300 270502
rect 479248 270438 479300 270444
rect 478880 269680 478932 269686
rect 478880 269622 478932 269628
rect 479260 264316 479288 270438
rect 480996 268252 481048 268258
rect 480996 268194 481048 268200
rect 481008 268138 481036 268194
rect 480456 268122 481036 268138
rect 480444 268116 481036 268122
rect 480496 268110 481036 268116
rect 480444 268058 480496 268064
rect 480904 267300 480956 267306
rect 480904 267242 480956 267248
rect 481088 267300 481140 267306
rect 481088 267242 481140 267248
rect 480916 266898 480944 267242
rect 480904 266892 480956 266898
rect 480904 266834 480956 266840
rect 481100 266762 481128 267242
rect 481088 266756 481140 266762
rect 481088 266698 481140 266704
rect 480076 265668 480128 265674
rect 480076 265610 480128 265616
rect 480088 264316 480116 265610
rect 481376 264330 481404 273362
rect 482560 272808 482612 272814
rect 482560 272750 482612 272756
rect 481548 267572 481600 267578
rect 481548 267514 481600 267520
rect 481732 267572 481784 267578
rect 481732 267514 481784 267520
rect 481560 266762 481588 267514
rect 481548 266756 481600 266762
rect 481548 266698 481600 266704
rect 480930 264302 481404 264330
rect 481744 264316 481772 267514
rect 482572 264316 482600 272750
rect 482940 272134 482968 274722
rect 482928 272128 482980 272134
rect 482928 272070 482980 272076
rect 483124 270366 483152 277366
rect 484320 273698 484348 277780
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483388 272128 483440 272134
rect 483388 272070 483440 272076
rect 483112 270360 483164 270366
rect 483112 270302 483164 270308
rect 483400 264316 483428 272070
rect 485516 271046 485544 277780
rect 486712 276010 486740 277780
rect 486700 276004 486752 276010
rect 486700 275946 486752 275952
rect 486884 276004 486936 276010
rect 486884 275946 486936 275952
rect 486896 273222 486924 275946
rect 487908 275874 487936 277780
rect 488736 277766 489118 277794
rect 489932 277766 490314 277794
rect 487896 275868 487948 275874
rect 487896 275810 487948 275816
rect 488540 275052 488592 275058
rect 488540 274994 488592 275000
rect 487988 273692 488040 273698
rect 487988 273634 488040 273640
rect 487068 273556 487120 273562
rect 487068 273498 487120 273504
rect 486884 273216 486936 273222
rect 486884 273158 486936 273164
rect 485504 271040 485556 271046
rect 485504 270982 485556 270988
rect 486700 270360 486752 270366
rect 486700 270302 486752 270308
rect 484216 269680 484268 269686
rect 484216 269622 484268 269628
rect 484228 264316 484256 269622
rect 485732 267472 485788 267481
rect 485732 267407 485734 267416
rect 485786 267407 485788 267416
rect 485872 267436 485924 267442
rect 485734 267378 485786 267384
rect 485872 267378 485924 267384
rect 485686 266928 485742 266937
rect 485686 266863 485742 266872
rect 485700 266626 485728 266863
rect 485688 266620 485740 266626
rect 485688 266562 485740 266568
rect 485044 265940 485096 265946
rect 485044 265882 485096 265888
rect 485056 264316 485084 265882
rect 485884 264316 485912 267378
rect 486054 266928 486110 266937
rect 486054 266863 486110 266872
rect 486068 266626 486096 266863
rect 486056 266620 486108 266626
rect 486056 266562 486108 266568
rect 486712 264316 486740 270302
rect 487080 267442 487108 273498
rect 487250 267472 487306 267481
rect 487068 267436 487120 267442
rect 487250 267407 487252 267416
rect 487068 267378 487120 267384
rect 487304 267407 487306 267416
rect 487252 267378 487304 267384
rect 488000 264330 488028 273634
rect 488356 272264 488408 272270
rect 488356 272206 488408 272212
rect 487554 264302 488028 264330
rect 488368 264316 488396 272206
rect 488552 268122 488580 274994
rect 488736 273086 488764 277766
rect 488724 273080 488776 273086
rect 488724 273022 488776 273028
rect 488724 271040 488776 271046
rect 488724 270982 488776 270988
rect 488540 268116 488592 268122
rect 488540 268058 488592 268064
rect 488736 266626 488764 270982
rect 489932 269142 489960 277766
rect 491496 274378 491524 277780
rect 492600 275058 492628 277780
rect 492588 275052 492640 275058
rect 492588 274994 492640 275000
rect 493796 274514 493824 277780
rect 494532 277766 495006 277794
rect 494532 275194 494560 277766
rect 494704 276004 494756 276010
rect 494704 275946 494756 275952
rect 495440 276004 495492 276010
rect 495440 275946 495492 275952
rect 494716 275194 494744 275946
rect 494520 275188 494572 275194
rect 494520 275130 494572 275136
rect 494704 275188 494756 275194
rect 494704 275130 494756 275136
rect 494704 275052 494756 275058
rect 494704 274994 494756 275000
rect 493784 274508 493836 274514
rect 493784 274450 493836 274456
rect 491484 274372 491536 274378
rect 491484 274314 491536 274320
rect 492496 274372 492548 274378
rect 492496 274314 492548 274320
rect 491208 273828 491260 273834
rect 491208 273770 491260 273776
rect 490392 270422 490788 270450
rect 490392 270366 490420 270422
rect 490380 270360 490432 270366
rect 490380 270302 490432 270308
rect 490564 270360 490616 270366
rect 490564 270302 490616 270308
rect 490576 269686 490604 270302
rect 490760 269686 490788 270422
rect 490564 269680 490616 269686
rect 490564 269622 490616 269628
rect 490748 269680 490800 269686
rect 490748 269622 490800 269628
rect 489920 269136 489972 269142
rect 489920 269078 489972 269084
rect 489184 267844 489236 267850
rect 489184 267786 489236 267792
rect 488724 266620 488776 266626
rect 488724 266562 488776 266568
rect 489196 264316 489224 267786
rect 490012 266620 490064 266626
rect 490012 266562 490064 266568
rect 490024 264316 490052 266562
rect 491220 264330 491248 273770
rect 491484 268116 491536 268122
rect 491484 268058 491536 268064
rect 491496 267442 491524 268058
rect 492310 267880 492366 267889
rect 492310 267815 492366 267824
rect 491484 267436 491536 267442
rect 491484 267378 491536 267384
rect 491668 267436 491720 267442
rect 491668 267378 491720 267384
rect 490866 264302 491248 264330
rect 491680 264316 491708 267378
rect 492324 266762 492352 267815
rect 492508 267442 492536 274314
rect 493324 273216 493376 273222
rect 493324 273158 493376 273164
rect 492496 267436 492548 267442
rect 492496 267378 492548 267384
rect 492680 267436 492732 267442
rect 492680 267378 492732 267384
rect 492692 266898 492720 267378
rect 492680 266892 492732 266898
rect 492680 266834 492732 266840
rect 492312 266756 492364 266762
rect 492312 266698 492364 266704
rect 492496 266756 492548 266762
rect 492496 266698 492548 266704
rect 492508 264316 492536 266698
rect 493336 264316 493364 273158
rect 494150 270056 494206 270065
rect 494150 269991 494206 270000
rect 494164 264316 494192 269991
rect 494716 268122 494744 274994
rect 495452 272406 495480 275946
rect 496188 274242 496216 277780
rect 496360 274508 496412 274514
rect 496360 274450 496412 274456
rect 496176 274236 496228 274242
rect 496176 274178 496228 274184
rect 495440 272400 495492 272406
rect 495440 272342 495492 272348
rect 494704 268116 494756 268122
rect 494704 268058 494756 268064
rect 496372 267734 496400 274450
rect 496636 273080 496688 273086
rect 496636 273022 496688 273028
rect 496280 267706 496400 267734
rect 494980 265804 495032 265810
rect 494980 265746 495032 265752
rect 494992 264316 495020 265746
rect 496280 264330 496308 267706
rect 495834 264302 496308 264330
rect 496648 264316 496676 273022
rect 497384 270910 497412 277780
rect 498200 275868 498252 275874
rect 498200 275810 498252 275816
rect 497372 270904 497424 270910
rect 497372 270846 497424 270852
rect 498212 267889 498240 275810
rect 498580 275058 498608 277780
rect 499592 277766 499790 277794
rect 500512 277766 500894 277794
rect 498568 275052 498620 275058
rect 498568 274994 498620 275000
rect 499592 268802 499620 277766
rect 500512 271726 500540 277766
rect 502076 275738 502104 277780
rect 502444 277766 503286 277794
rect 502064 275732 502116 275738
rect 502064 275674 502116 275680
rect 502248 275732 502300 275738
rect 502248 275674 502300 275680
rect 502260 275618 502288 275674
rect 501800 275602 502288 275618
rect 501788 275596 502288 275602
rect 501840 275590 502288 275596
rect 501788 275538 501840 275544
rect 501972 274236 502024 274242
rect 501972 274178 502024 274184
rect 501604 272400 501656 272406
rect 501604 272342 501656 272348
rect 500500 271720 500552 271726
rect 500500 271662 500552 271668
rect 500868 271720 500920 271726
rect 500868 271662 500920 271668
rect 499580 268796 499632 268802
rect 499580 268738 499632 268744
rect 500684 268796 500736 268802
rect 500684 268738 500736 268744
rect 499120 268116 499172 268122
rect 499120 268058 499172 268064
rect 498198 267880 498254 267889
rect 498198 267815 498254 267824
rect 497464 266892 497516 266898
rect 497464 266834 497516 266840
rect 497476 264316 497504 266834
rect 498568 266348 498620 266354
rect 498568 266290 498620 266296
rect 498580 264330 498608 266290
rect 498318 264302 498608 264330
rect 499132 264316 499160 268058
rect 499578 267200 499634 267209
rect 499578 267135 499580 267144
rect 499632 267135 499634 267144
rect 499764 267164 499816 267170
rect 499580 267106 499632 267112
rect 499764 267106 499816 267112
rect 499776 266898 499804 267106
rect 499764 266892 499816 266898
rect 499764 266834 499816 266840
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499960 264316 499988 266834
rect 500696 264330 500724 268738
rect 500880 266898 500908 271662
rect 501050 267200 501106 267209
rect 501050 267135 501106 267144
rect 501064 266898 501092 267135
rect 500868 266892 500920 266898
rect 500868 266834 500920 266840
rect 501052 266892 501104 266898
rect 501052 266834 501104 266840
rect 501616 266354 501644 272342
rect 501604 266348 501656 266354
rect 501604 266290 501656 266296
rect 501984 264330 502012 274178
rect 502444 268938 502472 277766
rect 504468 277394 504496 277780
rect 504468 277366 504588 277394
rect 504364 276004 504416 276010
rect 504364 275946 504416 275952
rect 504376 275466 504404 275946
rect 504364 275460 504416 275466
rect 504364 275402 504416 275408
rect 504560 271862 504588 277366
rect 504916 276004 504968 276010
rect 504916 275946 504968 275952
rect 504548 271856 504600 271862
rect 504548 271798 504600 271804
rect 504732 271856 504784 271862
rect 504732 271798 504784 271804
rect 504178 270600 504234 270609
rect 504178 270535 504234 270544
rect 504192 270230 504220 270535
rect 504180 270224 504232 270230
rect 504180 270166 504232 270172
rect 504364 270224 504416 270230
rect 504364 270166 504416 270172
rect 504376 269686 504404 270166
rect 504364 269680 504416 269686
rect 503074 269648 503130 269657
rect 504548 269680 504600 269686
rect 504364 269622 504416 269628
rect 504546 269648 504548 269657
rect 504600 269648 504602 269657
rect 503074 269583 503130 269592
rect 504546 269583 504602 269592
rect 502432 268932 502484 268938
rect 502432 268874 502484 268880
rect 503088 267578 503116 269583
rect 503260 269068 503312 269074
rect 503260 269010 503312 269016
rect 503076 267572 503128 267578
rect 503076 267514 503128 267520
rect 502800 266348 502852 266354
rect 502800 266290 502852 266296
rect 502812 264330 502840 266290
rect 500696 264302 500802 264330
rect 501630 264302 502012 264330
rect 502458 264302 502840 264330
rect 503272 264316 503300 269010
rect 503444 268932 503496 268938
rect 503444 268874 503496 268880
rect 503456 268666 503484 268874
rect 503444 268660 503496 268666
rect 503444 268602 503496 268608
rect 504180 268660 504232 268666
rect 504180 268602 504232 268608
rect 504192 268258 504220 268602
rect 504364 268524 504416 268530
rect 504364 268466 504416 268472
rect 504376 268258 504404 268466
rect 504180 268252 504232 268258
rect 504180 268194 504232 268200
rect 504364 268252 504416 268258
rect 504364 268194 504416 268200
rect 504744 267734 504772 271798
rect 504560 267706 504772 267734
rect 504180 267572 504232 267578
rect 504180 267514 504232 267520
rect 504192 267170 504220 267514
rect 504364 267436 504416 267442
rect 504364 267378 504416 267384
rect 504376 267170 504404 267378
rect 504180 267164 504232 267170
rect 504180 267106 504232 267112
rect 504364 267164 504416 267170
rect 504364 267106 504416 267112
rect 504560 264330 504588 267706
rect 504114 264302 504588 264330
rect 504928 264316 504956 275946
rect 505664 275874 505692 277780
rect 505652 275868 505704 275874
rect 505652 275810 505704 275816
rect 506860 275058 506888 277780
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 507032 276004 507084 276010
rect 507032 275946 507084 275952
rect 507044 275058 507072 275946
rect 507216 275868 507268 275874
rect 507216 275810 507268 275816
rect 505100 275052 505152 275058
rect 505100 274994 505152 275000
rect 506848 275052 506900 275058
rect 506848 274994 506900 275000
rect 507032 275052 507084 275058
rect 507032 274994 507084 275000
rect 505112 268938 505140 274994
rect 505100 268932 505152 268938
rect 505100 268874 505152 268880
rect 506112 268660 506164 268666
rect 506112 268602 506164 268608
rect 506124 264330 506152 268602
rect 507228 267578 507256 275810
rect 507676 270904 507728 270910
rect 507676 270846 507728 270852
rect 506480 267572 506532 267578
rect 506480 267514 506532 267520
rect 507216 267572 507268 267578
rect 507216 267514 507268 267520
rect 507400 267572 507452 267578
rect 507400 267514 507452 267520
rect 506492 267050 506520 267514
rect 506400 267022 506520 267050
rect 506400 266898 506428 267022
rect 506388 266892 506440 266898
rect 506388 266834 506440 266840
rect 506572 266892 506624 266898
rect 506572 266834 506624 266840
rect 505770 264302 506152 264330
rect 506584 264316 506612 266834
rect 507412 264316 507440 267514
rect 507688 266898 507716 270846
rect 507872 270609 507900 277366
rect 508044 276004 508096 276010
rect 508044 275946 508096 275952
rect 508056 271726 508084 275946
rect 509160 275738 509188 277780
rect 509620 277766 510370 277794
rect 509148 275732 509200 275738
rect 509148 275674 509200 275680
rect 508044 271720 508096 271726
rect 508044 271662 508096 271668
rect 508964 271720 509016 271726
rect 508964 271662 509016 271668
rect 507858 270600 507914 270609
rect 507858 270535 507914 270544
rect 508504 268932 508556 268938
rect 508504 268874 508556 268880
rect 507676 266892 507728 266898
rect 507676 266834 507728 266840
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 507872 266354 507900 266834
rect 507860 266348 507912 266354
rect 507860 266290 507912 266296
rect 508516 264330 508544 268874
rect 508254 264302 508544 264330
rect 508976 264330 509004 271662
rect 509620 268258 509648 277766
rect 511552 271590 511580 277780
rect 512748 275874 512776 277780
rect 513944 277394 513972 277780
rect 513852 277366 513972 277394
rect 512736 275868 512788 275874
rect 512736 275810 512788 275816
rect 512920 275868 512972 275874
rect 512920 275810 512972 275816
rect 512184 275732 512236 275738
rect 512184 275674 512236 275680
rect 512196 275330 512224 275674
rect 512184 275324 512236 275330
rect 512184 275266 512236 275272
rect 511540 271584 511592 271590
rect 511540 271526 511592 271532
rect 511908 271584 511960 271590
rect 511908 271526 511960 271532
rect 511724 271448 511776 271454
rect 511722 271416 511724 271425
rect 511776 271416 511778 271425
rect 511722 271351 511778 271360
rect 509882 269784 509938 269793
rect 509882 269719 509938 269728
rect 509608 268252 509660 268258
rect 509608 268194 509660 268200
rect 508976 264302 509082 264330
rect 509896 264316 509924 269719
rect 510712 268252 510764 268258
rect 510712 268194 510764 268200
rect 510724 264316 510752 268194
rect 511920 264330 511948 271526
rect 512932 267034 512960 275810
rect 513852 273970 513880 277366
rect 514024 276004 514076 276010
rect 514024 275946 514076 275952
rect 514036 275058 514064 275946
rect 514024 275052 514076 275058
rect 514024 274994 514076 275000
rect 513840 273964 513892 273970
rect 513840 273906 513892 273912
rect 513194 272368 513250 272377
rect 513194 272303 513250 272312
rect 512920 267028 512972 267034
rect 512920 266970 512972 266976
rect 512368 266484 512420 266490
rect 512368 266426 512420 266432
rect 511566 264302 511948 264330
rect 512380 264316 512408 266426
rect 513208 264316 513236 272303
rect 515140 271454 515168 277780
rect 515496 275868 515548 275874
rect 515496 275810 515548 275816
rect 515128 271448 515180 271454
rect 515312 271448 515364 271454
rect 515128 271390 515180 271396
rect 515310 271416 515312 271425
rect 515364 271416 515366 271425
rect 515310 271351 515366 271360
rect 514484 271312 514536 271318
rect 514484 271254 514536 271260
rect 514024 268660 514076 268666
rect 514024 268602 514076 268608
rect 514208 268660 514260 268666
rect 514208 268602 514260 268608
rect 514036 268258 514064 268602
rect 513840 268252 513892 268258
rect 513840 268194 513892 268200
rect 514024 268252 514076 268258
rect 514024 268194 514076 268200
rect 513852 268138 513880 268194
rect 514220 268138 514248 268602
rect 513852 268110 514248 268138
rect 513380 267028 513432 267034
rect 513380 266970 513432 266976
rect 513392 266490 513420 266970
rect 513380 266484 513432 266490
rect 513380 266426 513432 266432
rect 514496 264330 514524 271254
rect 515508 267734 515536 275810
rect 516244 275738 516272 277780
rect 516428 277766 517454 277794
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 516428 272678 516456 277766
rect 516784 275868 516836 275874
rect 516784 275810 516836 275816
rect 516598 274136 516654 274145
rect 516598 274071 516600 274080
rect 516652 274071 516654 274080
rect 516600 274042 516652 274048
rect 516416 272672 516468 272678
rect 516416 272614 516468 272620
rect 516600 272672 516652 272678
rect 516600 272614 516652 272620
rect 516612 272490 516640 272614
rect 514772 267706 515536 267734
rect 516060 272462 516640 272490
rect 514772 266506 514800 267706
rect 514680 266478 514800 266506
rect 514680 266422 514708 266478
rect 514668 266416 514720 266422
rect 514668 266358 514720 266364
rect 514852 266416 514904 266422
rect 514852 266358 514904 266364
rect 514050 264302 514524 264330
rect 514864 264316 514892 266358
rect 516060 264330 516088 272462
rect 516796 266422 516824 275810
rect 518440 274236 518492 274242
rect 518440 274178 518492 274184
rect 517058 274136 517114 274145
rect 517058 274071 517114 274080
rect 517072 273970 517100 274071
rect 517060 273964 517112 273970
rect 517060 273906 517112 273912
rect 518452 272377 518480 274178
rect 518438 272368 518494 272377
rect 518438 272303 518494 272312
rect 518636 271454 518664 277780
rect 519832 276010 519860 277780
rect 520292 277766 521042 277794
rect 521856 277766 522238 277794
rect 523144 277766 523434 277794
rect 524538 277766 524736 277794
rect 519820 276004 519872 276010
rect 519820 275946 519872 275952
rect 520004 276004 520056 276010
rect 520004 275946 520056 275952
rect 519188 275862 519584 275890
rect 519188 275738 519216 275862
rect 519556 275754 519584 275862
rect 519176 275732 519228 275738
rect 519176 275674 519228 275680
rect 519360 275732 519412 275738
rect 519556 275726 519768 275754
rect 519360 275674 519412 275680
rect 519372 275330 519400 275674
rect 519740 275602 519768 275726
rect 519544 275596 519596 275602
rect 519544 275538 519596 275544
rect 519728 275596 519780 275602
rect 519728 275538 519780 275544
rect 519556 275330 519584 275538
rect 519360 275324 519412 275330
rect 519360 275266 519412 275272
rect 519544 275324 519596 275330
rect 519544 275266 519596 275272
rect 520016 271674 520044 275946
rect 519924 271646 520044 271674
rect 518624 271448 518676 271454
rect 518624 271390 518676 271396
rect 518438 268560 518494 268569
rect 518438 268495 518494 268504
rect 518990 268560 519046 268569
rect 519046 268530 519400 268546
rect 519046 268524 519412 268530
rect 519046 268518 519360 268524
rect 518990 268495 519046 268504
rect 516966 267744 517022 267753
rect 516966 267679 517022 267688
rect 516784 266416 516836 266422
rect 516784 266358 516836 266364
rect 516980 264330 517008 267679
rect 517336 266484 517388 266490
rect 517336 266426 517388 266432
rect 515706 264302 516088 264330
rect 516534 264302 517008 264330
rect 517348 264316 517376 266426
rect 518452 264330 518480 268495
rect 519360 268466 519412 268472
rect 519174 268424 519230 268433
rect 518912 268394 519174 268410
rect 518900 268388 519174 268394
rect 518952 268382 519174 268388
rect 519174 268359 519230 268368
rect 518900 268330 518952 268336
rect 518990 267744 519046 267753
rect 518808 267708 518860 267714
rect 519924 267734 519952 271646
rect 520096 271448 520148 271454
rect 520096 271390 520148 271396
rect 518990 267679 518992 267688
rect 518808 267650 518860 267656
rect 519044 267679 519046 267688
rect 519832 267706 519952 267734
rect 518992 267650 519044 267656
rect 518820 267594 518848 267650
rect 518820 267566 519032 267594
rect 519004 267306 519032 267566
rect 518808 267300 518860 267306
rect 518808 267242 518860 267248
rect 518992 267300 519044 267306
rect 518992 267242 519044 267248
rect 518820 267186 518848 267242
rect 519174 267200 519230 267209
rect 518820 267158 519174 267186
rect 519174 267135 519230 267144
rect 518808 267028 518860 267034
rect 518808 266970 518860 266976
rect 518992 267028 519044 267034
rect 518992 266970 519044 266976
rect 518820 266354 518848 266970
rect 518808 266348 518860 266354
rect 518808 266290 518860 266296
rect 518190 264302 518480 264330
rect 519004 264316 519032 266970
rect 519832 264316 519860 267706
rect 520108 267034 520136 271390
rect 520292 268394 520320 277766
rect 521106 273728 521162 273737
rect 521106 273663 521162 273672
rect 520462 268424 520518 268433
rect 520280 268388 520332 268394
rect 520462 268359 520464 268368
rect 520280 268330 520332 268336
rect 520516 268359 520518 268368
rect 520464 268330 520516 268336
rect 520096 267028 520148 267034
rect 520096 266970 520148 266976
rect 520280 267028 520332 267034
rect 520280 266970 520332 266976
rect 520292 266354 520320 266970
rect 520280 266348 520332 266354
rect 520280 266290 520332 266296
rect 521120 264330 521148 273663
rect 521856 272950 521884 277766
rect 522948 276276 523000 276282
rect 522948 276218 523000 276224
rect 522960 275602 522988 276218
rect 522948 275596 523000 275602
rect 522948 275538 523000 275544
rect 523144 274922 523172 277766
rect 523132 274916 523184 274922
rect 523132 274858 523184 274864
rect 523316 274916 523368 274922
rect 523316 274858 523368 274864
rect 521844 272944 521896 272950
rect 521844 272886 521896 272892
rect 521474 272640 521530 272649
rect 521474 272575 521530 272584
rect 521488 267866 521516 272575
rect 522028 270904 522080 270910
rect 522026 270872 522028 270881
rect 522080 270872 522082 270881
rect 522026 270807 522082 270816
rect 523328 269793 523356 274858
rect 524708 274530 524736 277766
rect 525076 277766 525734 277794
rect 524880 276140 524932 276146
rect 524880 276082 524932 276088
rect 524892 275874 524920 276082
rect 524880 275868 524932 275874
rect 524880 275810 524932 275816
rect 524432 274502 524736 274530
rect 524432 274394 524460 274502
rect 524248 274366 524460 274394
rect 524248 273970 524276 274366
rect 524236 273964 524288 273970
rect 524236 273906 524288 273912
rect 524420 273964 524472 273970
rect 524420 273906 524472 273912
rect 524432 273850 524460 273906
rect 524248 273822 524460 273850
rect 524248 273737 524276 273822
rect 524234 273728 524290 273737
rect 524234 273663 524290 273672
rect 524386 273006 524736 273034
rect 524386 272950 524414 273006
rect 524374 272944 524426 272950
rect 524374 272886 524426 272892
rect 524512 272944 524564 272950
rect 524512 272886 524564 272892
rect 524524 272678 524552 272886
rect 524328 272672 524380 272678
rect 524328 272614 524380 272620
rect 524512 272672 524564 272678
rect 524512 272614 524564 272620
rect 523958 271688 524014 271697
rect 523958 271623 524014 271632
rect 523972 271454 524000 271623
rect 523960 271448 524012 271454
rect 523960 271390 524012 271396
rect 524144 271448 524196 271454
rect 524144 271390 524196 271396
rect 523314 269784 523370 269793
rect 523314 269719 523370 269728
rect 521658 269512 521714 269521
rect 521658 269447 521714 269456
rect 521488 267838 521608 267866
rect 521580 267734 521608 267838
rect 520674 264302 521148 264330
rect 521488 267706 521608 267734
rect 521672 267734 521700 269447
rect 521672 267706 521792 267734
rect 521488 264316 521516 267706
rect 521764 267170 521792 267706
rect 521752 267164 521804 267170
rect 521752 267106 521804 267112
rect 523132 267028 523184 267034
rect 523132 266970 523184 266976
rect 522672 266348 522724 266354
rect 522672 266290 522724 266296
rect 522684 264330 522712 266290
rect 522330 264302 522712 264330
rect 523144 264316 523172 266970
rect 524156 264330 524184 271390
rect 524340 267034 524368 272614
rect 524708 272542 524736 273006
rect 524880 272672 524932 272678
rect 524878 272640 524880 272649
rect 524932 272640 524934 272649
rect 524878 272575 524934 272584
rect 524512 272536 524564 272542
rect 524512 272478 524564 272484
rect 524696 272536 524748 272542
rect 524696 272478 524748 272484
rect 524524 272377 524552 272478
rect 524510 272368 524566 272377
rect 524510 272303 524566 272312
rect 525076 271810 525104 277766
rect 526916 276282 526944 277780
rect 527192 277766 528126 277794
rect 528848 277766 529322 277794
rect 526904 276276 526956 276282
rect 526904 276218 526956 276224
rect 525798 275768 525854 275777
rect 525798 275703 525854 275712
rect 524524 271782 525104 271810
rect 524524 271182 524552 271782
rect 524694 271688 524750 271697
rect 524694 271623 524750 271632
rect 524708 271182 524736 271623
rect 524512 271176 524564 271182
rect 524512 271118 524564 271124
rect 524696 271176 524748 271182
rect 524696 271118 524748 271124
rect 524788 270904 524840 270910
rect 524786 270872 524788 270881
rect 524840 270872 524842 270881
rect 524786 270807 524842 270816
rect 525812 269226 525840 275703
rect 526258 271008 526314 271017
rect 526258 270943 526314 270952
rect 526272 270774 526300 270943
rect 526260 270768 526312 270774
rect 526260 270710 526312 270716
rect 526444 270768 526496 270774
rect 526444 270710 526496 270716
rect 525720 269198 525840 269226
rect 525522 268696 525578 268705
rect 525522 268631 525578 268640
rect 524328 267028 524380 267034
rect 524328 266970 524380 266976
rect 524788 267028 524840 267034
rect 524788 266970 524840 266976
rect 523986 264302 524184 264330
rect 524800 264316 524828 266970
rect 525536 264330 525564 268631
rect 525720 267034 525748 269198
rect 525708 267028 525760 267034
rect 525708 266970 525760 266976
rect 525892 267028 525944 267034
rect 525892 266970 525944 266976
rect 525904 266354 525932 266970
rect 525892 266348 525944 266354
rect 525892 266290 525944 266296
rect 525536 264302 525642 264330
rect 526456 264316 526484 270710
rect 527192 268546 527220 277766
rect 527362 275768 527418 275777
rect 527362 275703 527364 275712
rect 527416 275703 527418 275712
rect 527364 275674 527416 275680
rect 528006 273864 528062 273873
rect 528006 273799 528062 273808
rect 527008 268518 527220 268546
rect 527008 268394 527036 268518
rect 526996 268388 527048 268394
rect 526996 268330 527048 268336
rect 527180 268388 527232 268394
rect 527180 268330 527232 268336
rect 527192 267209 527220 268330
rect 527178 267200 527234 267209
rect 527178 267135 527234 267144
rect 527640 266348 527692 266354
rect 527640 266290 527692 266296
rect 527652 264330 527680 266290
rect 527298 264302 527680 264330
rect 528020 264330 528048 273799
rect 528652 270768 528704 270774
rect 528650 270736 528652 270745
rect 528704 270736 528706 270745
rect 528650 270671 528706 270680
rect 528848 270314 528876 277766
rect 530504 275602 530532 277780
rect 530492 275596 530544 275602
rect 530492 275538 530544 275544
rect 530768 275596 530820 275602
rect 530768 275538 530820 275544
rect 529388 271448 529440 271454
rect 529388 271390 529440 271396
rect 529020 271312 529072 271318
rect 529020 271254 529072 271260
rect 529202 271280 529258 271289
rect 529032 270774 529060 271254
rect 529202 271215 529258 271224
rect 529020 270768 529072 270774
rect 529020 270710 529072 270716
rect 528664 270286 528876 270314
rect 528468 270088 528520 270094
rect 528468 270030 528520 270036
rect 528480 269770 528508 270030
rect 528664 269958 528692 270286
rect 528928 270224 528980 270230
rect 528928 270166 528980 270172
rect 528652 269952 528704 269958
rect 528652 269894 528704 269900
rect 528940 269770 528968 270166
rect 528480 269742 528968 269770
rect 529216 264330 529244 271215
rect 529400 271182 529428 271390
rect 529388 271176 529440 271182
rect 529388 271118 529440 271124
rect 529572 271176 529624 271182
rect 529572 271118 529624 271124
rect 529584 271017 529612 271118
rect 529570 271008 529626 271017
rect 529570 270943 529626 270952
rect 530780 269958 530808 275538
rect 531608 272377 531636 277780
rect 531594 272368 531650 272377
rect 531594 272303 531650 272312
rect 532804 271182 532832 277780
rect 532988 277766 534014 277794
rect 534184 277766 535210 277794
rect 535472 277766 536406 277794
rect 532792 271176 532844 271182
rect 532792 271118 532844 271124
rect 531410 270056 531466 270065
rect 531410 269991 531466 270000
rect 529756 269952 529808 269958
rect 529756 269894 529808 269900
rect 530768 269952 530820 269958
rect 530768 269894 530820 269900
rect 530952 269952 531004 269958
rect 530952 269894 531004 269900
rect 528020 264302 528126 264330
rect 528954 264302 529244 264330
rect 529768 264316 529796 269894
rect 530964 269521 530992 269894
rect 530950 269512 531006 269521
rect 530950 269447 531006 269456
rect 530950 269104 531006 269113
rect 530950 269039 531006 269048
rect 530964 264330 530992 269039
rect 530610 264302 530992 264330
rect 531424 264316 531452 269991
rect 532988 269958 533016 277766
rect 533894 274272 533950 274281
rect 533894 274207 533950 274216
rect 533908 274106 533936 274207
rect 533896 274100 533948 274106
rect 533896 274042 533948 274048
rect 534034 274100 534086 274106
rect 534034 274042 534086 274048
rect 534046 273986 534074 274042
rect 533908 273958 534074 273986
rect 533908 273873 533936 273958
rect 533894 273864 533950 273873
rect 533894 273799 533950 273808
rect 534184 273254 534212 277766
rect 534906 275768 534962 275777
rect 534906 275703 534962 275712
rect 534920 275602 534948 275703
rect 534908 275596 534960 275602
rect 534908 275538 534960 275544
rect 535090 275088 535146 275097
rect 535090 275023 535146 275032
rect 534184 273226 534396 273254
rect 534078 272776 534134 272785
rect 534078 272711 534134 272720
rect 534092 272626 534120 272711
rect 534000 272598 534120 272626
rect 534000 272542 534028 272598
rect 533988 272536 534040 272542
rect 533710 272504 533766 272513
rect 534172 272536 534224 272542
rect 533988 272478 534040 272484
rect 534170 272504 534172 272513
rect 534224 272504 534226 272513
rect 533710 272439 533766 272448
rect 534170 272439 534226 272448
rect 533160 271176 533212 271182
rect 533160 271118 533212 271124
rect 533172 270745 533200 271118
rect 533158 270736 533214 270745
rect 533158 270671 533214 270680
rect 533528 270224 533580 270230
rect 533528 270166 533580 270172
rect 532976 269952 533028 269958
rect 532976 269894 533028 269900
rect 533540 269793 533568 270166
rect 533526 269784 533582 269793
rect 533526 269719 533582 269728
rect 532238 267064 532294 267073
rect 532238 266999 532294 267008
rect 532252 264316 532280 266999
rect 533068 265124 533120 265130
rect 533068 265066 533120 265072
rect 533080 264316 533108 265066
rect 533724 264330 533752 272439
rect 533988 270224 534040 270230
rect 533988 270166 534040 270172
rect 534000 270042 534028 270166
rect 533908 270014 534028 270042
rect 533908 269113 533936 270014
rect 534368 269793 534396 273226
rect 534354 269784 534410 269793
rect 534354 269719 534410 269728
rect 533894 269104 533950 269113
rect 533894 269039 533950 269048
rect 533894 268696 533950 268705
rect 533950 268654 534074 268682
rect 533894 268631 533950 268640
rect 534046 268530 534074 268654
rect 533896 268524 533948 268530
rect 533896 268466 533948 268472
rect 534034 268524 534086 268530
rect 534034 268466 534086 268472
rect 533908 268138 533936 268466
rect 533908 268110 534074 268138
rect 533894 268016 533950 268025
rect 534046 267986 534074 268110
rect 533894 267951 533896 267960
rect 533948 267951 533950 267960
rect 534034 267980 534086 267986
rect 533896 267922 533948 267928
rect 534034 267922 534086 267928
rect 533986 267744 534042 267753
rect 533986 267679 533988 267688
rect 534040 267679 534042 267688
rect 534172 267708 534224 267714
rect 533988 267650 534040 267656
rect 534172 267650 534224 267656
rect 534184 267345 534212 267650
rect 533894 267336 533950 267345
rect 534170 267336 534226 267345
rect 533894 267271 533896 267280
rect 533948 267271 533950 267280
rect 534034 267300 534086 267306
rect 533896 267242 533948 267248
rect 534170 267271 534226 267280
rect 534034 267242 534086 267248
rect 534046 267186 534074 267242
rect 533908 267158 534074 267186
rect 533908 266354 533936 267158
rect 534080 266620 534132 266626
rect 534080 266562 534132 266568
rect 534092 266354 534120 266562
rect 533896 266348 533948 266354
rect 533896 266290 533948 266296
rect 534080 266348 534132 266354
rect 534080 266290 534132 266296
rect 535104 264330 535132 275023
rect 535472 268025 535500 277766
rect 537588 275330 537616 277780
rect 538784 277394 538812 277780
rect 539612 277766 539902 277794
rect 538784 277366 538904 277394
rect 538034 275768 538090 275777
rect 538034 275703 538090 275712
rect 538048 275602 538076 275703
rect 538036 275596 538088 275602
rect 538036 275538 538088 275544
rect 538218 275496 538274 275505
rect 538218 275431 538220 275440
rect 538272 275431 538274 275440
rect 538220 275402 538272 275408
rect 537576 275324 537628 275330
rect 537576 275266 537628 275272
rect 537760 275324 537812 275330
rect 538588 275324 538640 275330
rect 537760 275266 537812 275272
rect 538416 275284 538588 275312
rect 536746 273864 536802 273873
rect 536746 273799 536802 273808
rect 536564 269952 536616 269958
rect 536564 269894 536616 269900
rect 535918 269512 535974 269521
rect 535918 269447 535974 269456
rect 535458 268016 535514 268025
rect 535458 267951 535514 267960
rect 535932 264330 535960 269447
rect 536576 265130 536604 269894
rect 536564 265124 536616 265130
rect 536564 265066 536616 265072
rect 536760 264330 536788 273799
rect 537772 273254 537800 275266
rect 538416 275097 538444 275284
rect 538588 275266 538640 275272
rect 538402 275088 538458 275097
rect 538402 275023 538458 275032
rect 538678 275088 538734 275097
rect 538678 275023 538734 275032
rect 538218 274816 538274 274825
rect 538692 274786 538720 275023
rect 538218 274751 538274 274760
rect 538680 274780 538732 274786
rect 538232 274666 538260 274751
rect 538680 274722 538732 274728
rect 538140 274650 538260 274666
rect 538128 274644 538260 274650
rect 538180 274638 538260 274644
rect 538128 274586 538180 274592
rect 538876 273254 538904 277366
rect 539046 275496 539102 275505
rect 539046 275431 539102 275440
rect 539060 274786 539088 275431
rect 539048 274780 539100 274786
rect 539048 274722 539100 274728
rect 539048 274644 539100 274650
rect 539048 274586 539100 274592
rect 539060 274281 539088 274586
rect 539046 274272 539102 274281
rect 539046 274207 539102 274216
rect 537680 273226 537800 273254
rect 538692 273226 538904 273254
rect 537484 269816 537536 269822
rect 537484 269758 537536 269764
rect 537496 269550 537524 269758
rect 537484 269544 537536 269550
rect 537484 269486 537536 269492
rect 537024 269272 537076 269278
rect 537022 269240 537024 269249
rect 537076 269240 537078 269249
rect 537022 269175 537078 269184
rect 537680 267866 537708 273226
rect 538310 270600 538366 270609
rect 538310 270535 538366 270544
rect 538034 269784 538090 269793
rect 538034 269719 538090 269728
rect 537036 267838 537708 267866
rect 537036 267714 537064 267838
rect 537024 267708 537076 267714
rect 537024 267650 537076 267656
rect 537208 267708 537260 267714
rect 537208 267650 537260 267656
rect 533724 264302 533922 264330
rect 534750 264302 535132 264330
rect 535578 264302 535960 264330
rect 536406 264302 536788 264330
rect 537220 264316 537248 267650
rect 538048 264316 538076 269719
rect 538324 267753 538352 270535
rect 538692 269249 538720 273226
rect 538864 270632 538916 270638
rect 539612 270586 539640 277766
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 541820 277766 542294 277794
rect 543200 277766 543490 277794
rect 544304 277766 544686 277794
rect 540992 275466 541020 277366
rect 540980 275460 541032 275466
rect 540980 275402 541032 275408
rect 541164 275460 541216 275466
rect 541164 275402 541216 275408
rect 541176 275097 541204 275402
rect 541162 275088 541218 275097
rect 541162 275023 541218 275032
rect 540520 270768 540572 270774
rect 540520 270710 540572 270716
rect 538916 270580 539640 270586
rect 538864 270574 539640 270580
rect 538876 270558 539640 270574
rect 538864 270088 538916 270094
rect 538864 270030 538916 270036
rect 538876 269822 538904 270030
rect 538864 269816 538916 269822
rect 538864 269758 538916 269764
rect 538678 269240 538734 269249
rect 538678 269175 538734 269184
rect 539230 268152 539286 268161
rect 539230 268087 539286 268096
rect 538310 267744 538366 267753
rect 538310 267679 538366 267688
rect 539048 267708 539100 267714
rect 539048 267650 539100 267656
rect 539060 267306 539088 267650
rect 538864 267300 538916 267306
rect 538864 267242 538916 267248
rect 539048 267300 539100 267306
rect 539048 267242 539100 267248
rect 538678 266656 538734 266665
rect 538876 266626 538904 267242
rect 538678 266591 538680 266600
rect 538732 266591 538734 266600
rect 538864 266620 538916 266626
rect 538680 266562 538732 266568
rect 538864 266562 538916 266568
rect 539244 264330 539272 268087
rect 539692 267708 539744 267714
rect 539692 267650 539744 267656
rect 538890 264302 539272 264330
rect 539704 264316 539732 267650
rect 540532 264316 540560 270710
rect 541820 270094 541848 277766
rect 543200 274825 543228 277766
rect 544304 275466 544332 277766
rect 544292 275460 544344 275466
rect 544292 275402 544344 275408
rect 544476 275460 544528 275466
rect 544476 275402 544528 275408
rect 543186 274816 543242 274825
rect 543186 274751 543242 274760
rect 544488 272785 544516 275402
rect 545868 274786 545896 277780
rect 546512 277766 547078 277794
rect 547892 277766 548182 277794
rect 546040 275460 546092 275466
rect 546040 275402 546092 275408
rect 546224 275460 546276 275466
rect 546224 275402 546276 275408
rect 546052 274786 546080 275402
rect 545856 274780 545908 274786
rect 545856 274722 545908 274728
rect 546040 274780 546092 274786
rect 546040 274722 546092 274728
rect 544474 272776 544530 272785
rect 544474 272711 544530 272720
rect 543002 272504 543058 272513
rect 543002 272439 543058 272448
rect 540980 270088 541032 270094
rect 540980 270030 541032 270036
rect 541808 270088 541860 270094
rect 541808 270030 541860 270036
rect 541992 270088 542044 270094
rect 541992 270030 542044 270036
rect 540992 269550 541020 270030
rect 540980 269544 541032 269550
rect 540980 269486 541032 269492
rect 541348 269544 541400 269550
rect 542004 269521 542032 270030
rect 541348 269486 541400 269492
rect 541990 269512 542046 269521
rect 541360 264316 541388 269486
rect 541990 269447 542046 269456
rect 542174 267336 542230 267345
rect 542174 267271 542230 267280
rect 542188 264316 542216 267271
rect 543016 264316 543044 272439
rect 546236 271561 546264 275402
rect 543554 271552 543610 271561
rect 543554 271487 543610 271496
rect 546222 271552 546278 271561
rect 546222 271487 546278 271496
rect 543568 270774 543596 271487
rect 543556 270768 543608 270774
rect 543556 270710 543608 270716
rect 543694 270768 543746 270774
rect 543694 270710 543746 270716
rect 543554 270600 543610 270609
rect 543706 270586 543734 270710
rect 543610 270558 543734 270586
rect 543554 270535 543610 270544
rect 546512 269498 546540 277766
rect 546236 269470 546540 269498
rect 546236 269414 546264 269470
rect 546224 269408 546276 269414
rect 546224 269350 546276 269356
rect 546408 269408 546460 269414
rect 546408 269350 546460 269356
rect 543554 267744 543610 267753
rect 546420 267714 546448 269350
rect 547510 268424 547566 268433
rect 547510 268359 547512 268368
rect 547564 268359 547566 268368
rect 547696 268388 547748 268394
rect 547512 268330 547564 268336
rect 547696 268330 547748 268336
rect 547708 268161 547736 268330
rect 547694 268152 547750 268161
rect 547694 268087 547750 268096
rect 546590 267744 546646 267753
rect 543554 267679 543556 267688
rect 543608 267679 543610 267688
rect 543694 267708 543746 267714
rect 543556 267650 543608 267656
rect 543694 267650 543746 267656
rect 546408 267708 546460 267714
rect 546590 267679 546592 267688
rect 546408 267650 546460 267656
rect 546644 267679 546646 267688
rect 546592 267650 546644 267656
rect 543706 267594 543734 267650
rect 543568 267566 543734 267594
rect 543568 266665 543596 267566
rect 543554 266656 543610 266665
rect 543554 266591 543610 266600
rect 547892 266082 547920 277766
rect 549364 277394 549392 277780
rect 549640 277766 550574 277794
rect 549640 277394 549668 277766
rect 549272 277366 549392 277394
rect 549456 277366 549668 277394
rect 549272 268433 549300 277366
rect 549456 269278 549484 277366
rect 551756 271046 551784 277780
rect 552492 277766 552966 277794
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552492 271998 552520 277766
rect 552480 271992 552532 271998
rect 552480 271934 552532 271940
rect 552848 271992 552900 271998
rect 552848 271934 552900 271940
rect 551744 271040 551796 271046
rect 551744 270982 551796 270988
rect 552664 271040 552716 271046
rect 552664 270982 552716 270988
rect 552202 270736 552258 270745
rect 552202 270671 552258 270680
rect 552216 270502 552244 270671
rect 552676 270638 552704 270982
rect 552664 270632 552716 270638
rect 552664 270574 552716 270580
rect 552204 270496 552256 270502
rect 552204 270438 552256 270444
rect 552388 270496 552440 270502
rect 552388 270438 552440 270444
rect 552400 269906 552428 270438
rect 552308 269878 552428 269906
rect 552308 269822 552336 269878
rect 552296 269816 552348 269822
rect 552296 269758 552348 269764
rect 552480 269816 552532 269822
rect 552480 269758 552532 269764
rect 552492 269634 552520 269758
rect 552400 269606 552520 269634
rect 552400 269550 552428 269606
rect 552388 269544 552440 269550
rect 552388 269486 552440 269492
rect 551928 269408 551980 269414
rect 551980 269356 552336 269362
rect 551928 269350 552336 269356
rect 551940 269334 552336 269350
rect 552308 269278 552336 269334
rect 549444 269272 549496 269278
rect 549444 269214 549496 269220
rect 549628 269272 549680 269278
rect 549628 269214 549680 269220
rect 552296 269272 552348 269278
rect 552296 269214 552348 269220
rect 549258 268424 549314 268433
rect 549258 268359 549314 268368
rect 549640 266422 549668 269214
rect 552860 267442 552888 271934
rect 553412 270745 553440 277766
rect 553398 270736 553454 270745
rect 553398 270671 553454 270680
rect 553032 269680 553084 269686
rect 553032 269622 553084 269628
rect 553044 269414 553072 269622
rect 553032 269408 553084 269414
rect 553032 269350 553084 269356
rect 552848 267436 552900 267442
rect 552848 267378 552900 267384
rect 552848 266756 552900 266762
rect 552848 266698 552900 266704
rect 552860 266490 552888 266698
rect 552848 266484 552900 266490
rect 552848 266426 552900 266432
rect 549628 266416 549680 266422
rect 549628 266358 549680 266364
rect 547880 266076 547932 266082
rect 547880 266018 547932 266024
rect 554792 265674 554820 277766
rect 556448 273426 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 273420 556488 273426
rect 556436 273362 556488 273368
rect 557552 269414 557580 277366
rect 558840 274786 558868 277780
rect 558828 274780 558880 274786
rect 558828 274722 558880 274728
rect 560036 272134 560064 277780
rect 560312 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 272128 560076 272134
rect 560024 272070 560076 272076
rect 560312 270366 560340 277766
rect 560300 270360 560352 270366
rect 560300 270302 560352 270308
rect 558920 269680 558972 269686
rect 558920 269622 558972 269628
rect 557540 269408 557592 269414
rect 557540 269350 557592 269356
rect 558932 266626 558960 269622
rect 558920 266620 558972 266626
rect 558920 266562 558972 266568
rect 561692 265946 561720 277766
rect 563532 273562 563560 277780
rect 564452 277766 564742 277794
rect 563520 273556 563572 273562
rect 563520 273498 563572 273504
rect 564452 270502 564480 277766
rect 565924 273698 565952 277780
rect 565912 273692 565964 273698
rect 565912 273634 565964 273640
rect 567120 272270 567148 277780
rect 567672 277766 568330 277794
rect 568592 277766 569526 277794
rect 567108 272264 567160 272270
rect 567108 272206 567160 272212
rect 564440 270496 564492 270502
rect 564440 270438 564492 270444
rect 567672 267850 567700 277766
rect 568592 269550 568620 277766
rect 570708 277394 570736 277780
rect 570616 277366 570736 277394
rect 570616 273834 570644 277366
rect 570788 274780 570840 274786
rect 570788 274722 570840 274728
rect 570800 274378 570828 274722
rect 571812 274650 571840 277780
rect 572732 277766 573022 277794
rect 570972 274644 571024 274650
rect 570972 274586 571024 274592
rect 571800 274644 571852 274650
rect 571800 274586 571852 274592
rect 570984 274378 571012 274586
rect 570788 274372 570840 274378
rect 570788 274314 570840 274320
rect 570972 274372 571024 274378
rect 570972 274314 571024 274320
rect 570604 273828 570656 273834
rect 570604 273770 570656 273776
rect 570604 273692 570656 273698
rect 570604 273634 570656 273640
rect 568580 269544 568632 269550
rect 568580 269486 568632 269492
rect 567660 267844 567712 267850
rect 567660 267786 567712 267792
rect 570616 266898 570644 273634
rect 572732 269686 572760 277766
rect 574204 273222 574232 277780
rect 574940 277766 575414 277794
rect 575860 277766 576610 277794
rect 574192 273216 574244 273222
rect 574192 273158 574244 273164
rect 574940 270337 574968 277766
rect 574926 270328 574982 270337
rect 574926 270263 574982 270272
rect 572720 269680 572772 269686
rect 572720 269622 572772 269628
rect 570604 266892 570656 266898
rect 570604 266834 570656 266840
rect 561680 265940 561732 265946
rect 561680 265882 561732 265888
rect 575860 265810 575888 277766
rect 577792 274650 577820 277780
rect 578528 277766 578910 277794
rect 577780 274644 577832 274650
rect 577780 274586 577832 274592
rect 578528 273086 578556 277766
rect 578884 273216 578936 273222
rect 578884 273158 578936 273164
rect 578516 273080 578568 273086
rect 578516 273022 578568 273028
rect 578896 267578 578924 273158
rect 580092 271998 580120 277780
rect 580264 273080 580316 273086
rect 580264 273022 580316 273028
rect 580080 271992 580132 271998
rect 580080 271934 580132 271940
rect 579620 268116 579672 268122
rect 579620 268058 579672 268064
rect 579632 267850 579660 268058
rect 579620 267844 579672 267850
rect 579620 267786 579672 267792
rect 580276 267714 580304 273022
rect 581288 272406 581316 277780
rect 582484 277394 582512 277780
rect 582392 277366 582512 277394
rect 581276 272400 581328 272406
rect 581276 272342 581328 272348
rect 581288 269198 581684 269226
rect 581288 268802 581316 269198
rect 581656 269074 581684 269198
rect 581460 269068 581512 269074
rect 581460 269010 581512 269016
rect 581644 269068 581696 269074
rect 581644 269010 581696 269016
rect 581276 268796 581328 268802
rect 581276 268738 581328 268744
rect 581472 268122 581500 269010
rect 581644 268796 581696 268802
rect 581644 268738 581696 268744
rect 581460 268116 581512 268122
rect 581460 268058 581512 268064
rect 581656 267986 581684 268738
rect 581644 267980 581696 267986
rect 581644 267922 581696 267928
rect 582392 267850 582420 277366
rect 583680 275058 583708 277780
rect 584140 277766 584890 277794
rect 583668 275052 583720 275058
rect 583668 274994 583720 275000
rect 584140 269074 584168 277766
rect 585784 274508 585836 274514
rect 585784 274450 585836 274456
rect 584128 269068 584180 269074
rect 584128 269010 584180 269016
rect 582380 267844 582432 267850
rect 582380 267786 582432 267792
rect 580264 267708 580316 267714
rect 580264 267650 580316 267656
rect 578884 267572 578936 267578
rect 578884 267514 578936 267520
rect 585796 267170 585824 274450
rect 586072 274378 586100 277780
rect 586060 274372 586112 274378
rect 586060 274314 586112 274320
rect 587176 273834 587204 277780
rect 587912 277766 588386 277794
rect 587164 273828 587216 273834
rect 587164 273770 587216 273776
rect 587912 268122 587940 277766
rect 589568 271862 589596 277780
rect 590764 275194 590792 277780
rect 591040 277766 591974 277794
rect 590752 275188 590804 275194
rect 590752 275130 590804 275136
rect 589556 271856 589608 271862
rect 589556 271798 589608 271804
rect 590660 269068 590712 269074
rect 590660 269010 590712 269016
rect 590672 268666 590700 269010
rect 590660 268660 590712 268666
rect 590660 268602 590712 268608
rect 591040 268258 591068 277766
rect 591488 271720 591540 271726
rect 591488 271662 591540 271668
rect 591500 271046 591528 271662
rect 591488 271040 591540 271046
rect 591488 270982 591540 270988
rect 593156 270910 593184 277780
rect 594352 273222 594380 277780
rect 594812 277766 595470 277794
rect 594340 273216 594392 273222
rect 594340 273158 594392 273164
rect 593144 270904 593196 270910
rect 593144 270846 593196 270852
rect 594812 268938 594840 277766
rect 596652 271862 596680 277780
rect 597848 274922 597876 277780
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597836 274916 597888 274922
rect 597836 274858 597888 274864
rect 598952 274666 598980 277366
rect 598860 274638 598980 274666
rect 596640 271856 596692 271862
rect 596640 271798 596692 271804
rect 594800 268932 594852 268938
rect 594800 268874 594852 268880
rect 598860 268802 598888 274638
rect 600240 271590 600268 277780
rect 601436 274378 601464 277780
rect 601424 274372 601476 274378
rect 601424 274314 601476 274320
rect 602540 274242 602568 277780
rect 602528 274236 602580 274242
rect 602528 274178 602580 274184
rect 603736 271726 603764 277780
rect 604932 276010 604960 277780
rect 604920 276004 604972 276010
rect 604920 275946 604972 275952
rect 606128 272814 606156 277780
rect 606116 272808 606168 272814
rect 606116 272750 606168 272756
rect 603724 271720 603776 271726
rect 603724 271662 603776 271668
rect 600228 271584 600280 271590
rect 600228 271526 600280 271532
rect 607324 270774 607352 277780
rect 607600 277766 608534 277794
rect 608704 277766 609730 277794
rect 607312 270768 607364 270774
rect 607312 270710 607364 270716
rect 607600 269278 607628 277766
rect 607864 271584 607916 271590
rect 607864 271526 607916 271532
rect 607588 269272 607640 269278
rect 607588 269214 607640 269220
rect 598848 268796 598900 268802
rect 598848 268738 598900 268744
rect 591028 268252 591080 268258
rect 591028 268194 591080 268200
rect 587900 268116 587952 268122
rect 587900 268058 587952 268064
rect 607876 267345 607904 271526
rect 608704 268666 608732 277766
rect 610820 271454 610848 277780
rect 612016 275874 612044 277780
rect 612004 275868 612056 275874
rect 612004 275810 612056 275816
rect 611360 275188 611412 275194
rect 611360 275130 611412 275136
rect 611372 272950 611400 275130
rect 613212 273970 613240 277780
rect 613384 274236 613436 274242
rect 613384 274178 613436 274184
rect 613200 273964 613252 273970
rect 613200 273906 613252 273912
rect 611360 272944 611412 272950
rect 611360 272886 611412 272892
rect 610808 271448 610860 271454
rect 610808 271390 610860 271396
rect 608692 268660 608744 268666
rect 608692 268602 608744 268608
rect 607862 267336 607918 267345
rect 607862 267271 607918 267280
rect 585784 267164 585836 267170
rect 585784 267106 585836 267112
rect 613396 267034 613424 274178
rect 614408 272678 614436 277780
rect 615604 274242 615632 277780
rect 616800 275194 616828 277780
rect 616788 275188 616840 275194
rect 616788 275130 616840 275136
rect 615592 274236 615644 274242
rect 615592 274178 615644 274184
rect 614396 272672 614448 272678
rect 614396 272614 614448 272620
rect 617996 271318 618024 277780
rect 619100 275738 619128 277780
rect 619652 277766 620310 277794
rect 619088 275732 619140 275738
rect 619088 275674 619140 275680
rect 619180 275188 619232 275194
rect 619180 275130 619232 275136
rect 619192 274106 619220 275130
rect 619180 274100 619232 274106
rect 619180 274042 619232 274048
rect 617984 271312 618036 271318
rect 617984 271254 618036 271260
rect 619652 268530 619680 277766
rect 621492 271182 621520 277780
rect 622412 277766 622702 277794
rect 621480 271176 621532 271182
rect 621480 271118 621532 271124
rect 621664 271176 621716 271182
rect 621664 271118 621716 271124
rect 619640 268524 619692 268530
rect 619640 268466 619692 268472
rect 621676 267306 621704 271118
rect 621664 267300 621716 267306
rect 621664 267242 621716 267248
rect 622412 267034 622440 277766
rect 623884 275194 623912 277780
rect 623872 275188 623924 275194
rect 623872 275130 623924 275136
rect 625080 271153 625108 277780
rect 626184 275602 626212 277780
rect 626552 277766 627394 277794
rect 627932 277766 628590 277794
rect 629312 277766 629786 277794
rect 630692 277766 630982 277794
rect 626172 275596 626224 275602
rect 626172 275538 626224 275544
rect 625066 271144 625122 271153
rect 625066 271079 625122 271088
rect 626552 270230 626580 277766
rect 626540 270224 626592 270230
rect 626540 270166 626592 270172
rect 627932 270065 627960 277766
rect 627918 270056 627974 270065
rect 627918 269991 627974 270000
rect 629312 267073 629340 277766
rect 630692 269958 630720 277766
rect 632164 272542 632192 277780
rect 633360 275330 633388 277780
rect 633636 277766 634478 277794
rect 633348 275324 633400 275330
rect 633348 275266 633400 275272
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 633636 270094 633664 277766
rect 635660 273873 635688 277780
rect 635646 273864 635702 273873
rect 635646 273799 635702 273808
rect 636856 271182 636884 277780
rect 637592 277766 638066 277794
rect 638972 277766 639262 277794
rect 636844 271176 636896 271182
rect 636844 271118 636896 271124
rect 633624 270088 633676 270094
rect 633624 270030 633676 270036
rect 630680 269952 630732 269958
rect 630680 269894 630732 269900
rect 637592 269793 637620 277766
rect 637578 269784 637634 269793
rect 637578 269719 637634 269728
rect 638972 268394 639000 277766
rect 640444 273086 640472 277780
rect 641640 275466 641668 277780
rect 641916 277766 642758 277794
rect 641628 275460 641680 275466
rect 641628 275402 641680 275408
rect 640432 273080 640484 273086
rect 640432 273022 640484 273028
rect 641916 269822 641944 277766
rect 643940 271590 643968 277780
rect 645136 272513 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645122 272504 645178 272513
rect 645122 272439 645178 272448
rect 643928 271584 643980 271590
rect 643928 271526 643980 271532
rect 641904 269816 641956 269822
rect 641904 269758 641956 269764
rect 638960 268388 639012 268394
rect 638960 268330 639012 268336
rect 629298 267064 629354 267073
rect 613384 267028 613436 267034
rect 613384 266970 613436 266976
rect 622400 267028 622452 267034
rect 629298 266999 629354 267008
rect 622400 266970 622452 266976
rect 575848 265804 575900 265810
rect 575848 265746 575900 265752
rect 554780 265668 554832 265674
rect 554780 265610 554832 265616
rect 558184 265668 558236 265674
rect 558184 265610 558236 265616
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553674 255640 553730 255649
rect 553674 255575 553730 255584
rect 553490 251288 553546 251297
rect 553490 251223 553492 251232
rect 553544 251223 553546 251232
rect 553492 251194 553544 251200
rect 553688 249082 553716 255575
rect 554502 253464 554558 253473
rect 554502 253399 554504 253408
rect 554556 253399 554558 253408
rect 554504 253370 554556 253376
rect 555424 251252 555476 251258
rect 555424 251194 555476 251200
rect 553858 249112 553914 249121
rect 553676 249076 553728 249082
rect 553858 249047 553914 249056
rect 553676 249018 553728 249024
rect 553872 246362 553900 249047
rect 554410 246936 554466 246945
rect 554410 246871 554466 246880
rect 553860 246356 553912 246362
rect 553860 246298 553912 246304
rect 554424 245682 554452 246871
rect 554412 245676 554464 245682
rect 554412 245618 554464 245624
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 553950 242584 554006 242593
rect 553950 242519 554006 242528
rect 553964 241534 553992 242519
rect 553952 241528 554004 241534
rect 553952 241470 554004 241476
rect 553858 240408 553914 240417
rect 553858 240343 553914 240352
rect 553872 240174 553900 240343
rect 553860 240168 553912 240174
rect 553860 240110 553912 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 186898 231798 187096 231826
rect 140792 231662 141174 231690
rect 141528 231662 141818 231690
rect 90364 230444 90416 230450
rect 90364 230386 90416 230392
rect 88248 230036 88300 230042
rect 88248 229978 88300 229984
rect 74448 229900 74500 229906
rect 74448 229842 74500 229848
rect 67548 229764 67600 229770
rect 67548 229706 67600 229712
rect 66168 228404 66220 228410
rect 66168 228346 66220 228352
rect 64788 225752 64840 225758
rect 64788 225694 64840 225700
rect 62946 222864 63002 222873
rect 62946 222799 63002 222808
rect 64604 221468 64656 221474
rect 64604 221410 64656 221416
rect 63132 220108 63184 220114
rect 63132 220050 63184 220056
rect 62764 218204 62816 218210
rect 62764 218146 62816 218152
rect 63144 217274 63172 220050
rect 64616 219434 64644 221410
rect 64800 219434 64828 225694
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 62270 217110 62344 217138
rect 63098 217246 63172 217274
rect 62270 216988 62298 217110
rect 63098 216988 63126 217246
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 228346
rect 66444 220244 66496 220250
rect 66444 220186 66496 220192
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64708 217246 64782 217274
rect 63926 217110 64000 217138
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217274 66484 220186
rect 67560 219434 67588 229706
rect 73066 226944 73122 226953
rect 73066 226879 73122 226888
rect 69572 226160 69624 226166
rect 69572 226102 69624 226108
rect 68926 224224 68982 224233
rect 68926 224159 68982 224168
rect 68100 221740 68152 221746
rect 68100 221682 68152 221688
rect 67284 219406 67588 219434
rect 67284 217274 67312 219406
rect 68112 217274 68140 221682
rect 68940 217274 68968 224159
rect 69584 218618 69612 226102
rect 71412 221876 71464 221882
rect 71412 221818 71464 221824
rect 69754 220144 69810 220153
rect 69754 220079 69810 220088
rect 69572 218612 69624 218618
rect 69572 218554 69624 218560
rect 69768 217274 69796 220079
rect 70584 219020 70636 219026
rect 70584 218962 70636 218968
rect 65582 217110 65656 217138
rect 66410 217246 66484 217274
rect 67238 217246 67312 217274
rect 68066 217246 68140 217274
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217246
rect 67238 216988 67266 217246
rect 68066 216988 68094 217246
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 218962
rect 71424 217274 71452 221818
rect 72882 220416 72938 220425
rect 72882 220351 72938 220360
rect 72896 219434 72924 220351
rect 73080 219434 73108 226879
rect 72240 219428 72292 219434
rect 72896 219406 73016 219434
rect 73080 219428 73212 219434
rect 73080 219406 73160 219428
rect 72240 219370 72292 219376
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 219370
rect 72988 217274 73016 219406
rect 73160 219370 73212 219376
rect 74460 218074 74488 229842
rect 82084 228676 82136 228682
rect 82084 228618 82136 228624
rect 79966 228304 80022 228313
rect 79966 228239 80022 228248
rect 75828 227180 75880 227186
rect 75828 227122 75880 227128
rect 75552 218340 75604 218346
rect 75552 218282 75604 218288
rect 73896 218068 73948 218074
rect 73896 218010 73948 218016
rect 74448 218068 74500 218074
rect 74448 218010 74500 218016
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72988 217246 73062 217274
rect 72206 217110 72280 217138
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73908 217138 73936 218010
rect 74736 217138 74764 218010
rect 75564 217138 75592 218282
rect 75840 218074 75868 227122
rect 76564 223984 76616 223990
rect 76564 223926 76616 223932
rect 76380 220380 76432 220386
rect 76380 220322 76432 220328
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220322
rect 76576 218890 76604 223926
rect 78588 223168 78640 223174
rect 78588 223110 78640 223116
rect 76564 218884 76616 218890
rect 76564 218826 76616 218832
rect 77208 218748 77260 218754
rect 77208 218690 77260 218696
rect 73862 217110 73936 217138
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 73862 216988 73890 217110
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218690
rect 78600 218074 78628 223110
rect 79692 218204 79744 218210
rect 79692 218146 79744 218152
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217138 79732 218146
rect 79980 218074 80008 228239
rect 81348 223440 81400 223446
rect 81348 223382 81400 223388
rect 80520 219428 80572 219434
rect 80520 219370 80572 219376
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217138 80560 219370
rect 81360 217274 81388 223382
rect 82096 218210 82124 228618
rect 86868 227316 86920 227322
rect 86868 227258 86920 227264
rect 83464 226296 83516 226302
rect 83464 226238 83516 226244
rect 82728 224392 82780 224398
rect 82728 224334 82780 224340
rect 82084 218204 82136 218210
rect 82084 218146 82136 218152
rect 82740 218074 82768 224334
rect 83004 220516 83056 220522
rect 83004 220458 83056 220464
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 82728 218068 82780 218074
rect 82728 218010 82780 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217110 79732 217138
rect 80486 217110 80560 217138
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217110
rect 80486 216988 80514 217110
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220458
rect 83476 218346 83504 226238
rect 85488 222760 85540 222766
rect 85488 222702 85540 222708
rect 85304 219156 85356 219162
rect 85304 219098 85356 219104
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218340 83516 218346
rect 83464 218282 83516 218288
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 84672 217138 84700 218010
rect 85316 217274 85344 219098
rect 85500 218074 85528 222702
rect 86880 218074 86908 227258
rect 87972 223576 88024 223582
rect 87972 223518 88024 223524
rect 85488 218068 85540 218074
rect 85488 218010 85540 218016
rect 86316 218068 86368 218074
rect 86316 218010 86368 218016
rect 86868 218068 86920 218074
rect 86868 218010 86920 218016
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 85316 217246 85482 217274
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86328 217138 86356 218010
rect 87156 217138 87184 218010
rect 87984 217274 88012 223518
rect 88260 218074 88288 229978
rect 90376 229094 90404 230386
rect 118424 230308 118476 230314
rect 118424 230250 118476 230256
rect 111064 230172 111116 230178
rect 111064 230114 111116 230120
rect 103610 229800 103666 229809
rect 103610 229735 103666 229744
rect 92480 229356 92532 229362
rect 92480 229298 92532 229304
rect 90284 229066 90404 229094
rect 89628 227452 89680 227458
rect 89628 227394 89680 227400
rect 89444 223032 89496 223038
rect 89444 222974 89496 222980
rect 89456 218074 89484 222974
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 86282 217110 86356 217138
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 86282 216988 86310 217110
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227394
rect 90284 219434 90312 229066
rect 92492 225758 92520 229298
rect 97908 228948 97960 228954
rect 97908 228890 97960 228896
rect 96252 228676 96304 228682
rect 96252 228618 96304 228624
rect 93768 226024 93820 226030
rect 93768 225966 93820 225972
rect 92480 225752 92532 225758
rect 92480 225694 92532 225700
rect 92112 223304 92164 223310
rect 92112 223246 92164 223252
rect 91284 220652 91336 220658
rect 91284 220594 91336 220600
rect 90272 219428 90324 219434
rect 90272 219370 90324 219376
rect 90456 219428 90508 219434
rect 90456 219370 90508 219376
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 219370
rect 91296 217274 91324 220594
rect 92124 217274 92152 223246
rect 93780 218618 93808 225966
rect 95148 225888 95200 225894
rect 95148 225830 95200 225836
rect 92940 218612 92992 218618
rect 92940 218554 92992 218560
rect 93768 218612 93820 218618
rect 93768 218554 93820 218560
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218554
rect 93768 218476 93820 218482
rect 93768 218418 93820 218424
rect 93780 217138 93808 218418
rect 95160 218074 95188 225830
rect 95424 222012 95476 222018
rect 95424 221954 95476 221960
rect 94596 218068 94648 218074
rect 94596 218010 94648 218016
rect 95148 218068 95200 218074
rect 95148 218010 95200 218016
rect 94608 217138 94636 218010
rect 95436 217274 95464 221954
rect 96264 217274 96292 228618
rect 97724 220788 97776 220794
rect 97724 220730 97776 220736
rect 97736 219434 97764 220730
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217110 94636 217138
rect 95390 217246 95464 217274
rect 96218 217246 96292 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217110
rect 95390 216988 95418 217246
rect 96218 216988 96246 217246
rect 97092 217138 97120 218010
rect 97828 217274 97856 219406
rect 97920 218090 97948 228890
rect 102048 228268 102100 228274
rect 102048 228210 102100 228216
rect 100668 227588 100720 227594
rect 100668 227530 100720 227536
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97920 218074 98040 218090
rect 99300 218074 99328 222566
rect 100392 218340 100444 218346
rect 100392 218282 100444 218288
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218282
rect 100680 218074 100708 227530
rect 101862 221504 101918 221513
rect 101862 221439 101918 221448
rect 101876 219434 101904 221439
rect 101876 219406 101996 219434
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101220 218068 101272 218074
rect 101220 218010 101272 218016
rect 101232 217138 101260 218010
rect 101968 217274 101996 219406
rect 102060 218090 102088 228210
rect 103428 225480 103480 225486
rect 103428 225422 103480 225428
rect 102060 218074 102180 218090
rect 103440 218074 103468 225422
rect 103624 224534 103652 229735
rect 106188 229084 106240 229090
rect 106188 229026 106240 229032
rect 106004 225344 106056 225350
rect 106004 225286 106056 225292
rect 103612 224528 103664 224534
rect 103612 224470 103664 224476
rect 104808 224120 104860 224126
rect 104808 224062 104860 224068
rect 104532 222012 104584 222018
rect 104532 221954 104584 221960
rect 102060 218068 102192 218074
rect 102060 218062 102140 218068
rect 102140 218010 102192 218016
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 103704 218068 103756 218074
rect 103704 218010 103756 218016
rect 101968 217246 102042 217274
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217110 101260 217138
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217110
rect 102014 216988 102042 217246
rect 102888 217138 102916 218010
rect 103716 217138 103744 218010
rect 104544 217274 104572 221954
rect 104820 218074 104848 224062
rect 105820 219496 105872 219502
rect 105820 219438 105872 219444
rect 105832 218346 105860 219438
rect 105820 218340 105872 218346
rect 105820 218282 105872 218288
rect 106016 218074 106044 225286
rect 104808 218068 104860 218074
rect 104808 218010 104860 218016
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 229026
rect 107016 228948 107068 228954
rect 107016 228890 107068 228896
rect 107028 228834 107056 228890
rect 106660 228818 107056 228834
rect 106648 228812 107056 228818
rect 106700 228806 107056 228812
rect 106648 228754 106700 228760
rect 110144 227724 110196 227730
rect 110144 227666 110196 227672
rect 106924 226908 106976 226914
rect 106924 226850 106976 226856
rect 106936 219298 106964 226850
rect 108304 225752 108356 225758
rect 108304 225694 108356 225700
rect 108316 225486 108344 225694
rect 108304 225480 108356 225486
rect 108304 225422 108356 225428
rect 108672 224528 108724 224534
rect 108672 224470 108724 224476
rect 107844 221196 107896 221202
rect 107844 221138 107896 221144
rect 106924 219292 106976 219298
rect 106924 219234 106976 219240
rect 107016 218340 107068 218346
rect 107016 218282 107068 218288
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218282
rect 107856 217274 107884 221138
rect 108028 220924 108080 220930
rect 108028 220866 108080 220872
rect 108040 220658 108068 220866
rect 108028 220652 108080 220658
rect 108028 220594 108080 220600
rect 108684 217274 108712 224470
rect 110156 218074 110184 227666
rect 111076 219434 111104 230114
rect 115756 229220 115808 229226
rect 115756 229162 115808 229168
rect 115572 228948 115624 228954
rect 115572 228890 115624 228896
rect 112996 228132 113048 228138
rect 112996 228074 113048 228080
rect 112812 222896 112864 222902
rect 112812 222838 112864 222844
rect 111248 219972 111300 219978
rect 111248 219914 111300 219920
rect 111260 219434 111288 219914
rect 110984 219406 111104 219434
rect 111168 219406 111288 219434
rect 110984 218074 111012 219406
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 110328 218068 110380 218074
rect 110328 218010 110380 218016
rect 110972 218068 111024 218074
rect 110972 218010 111024 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217138 110368 218010
rect 111168 217274 111196 219406
rect 112824 218074 112852 222838
rect 111984 218068 112036 218074
rect 111984 218010 112036 218016
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 109466 217110 109540 217138
rect 110294 217110 110368 217138
rect 111122 217246 111196 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217110
rect 111122 216988 111150 217246
rect 111996 217138 112024 218010
rect 113008 217274 113036 228074
rect 115584 228002 115612 228890
rect 115768 228138 115796 229162
rect 116032 229084 116084 229090
rect 116032 229026 116084 229032
rect 116044 228970 116072 229026
rect 116044 228954 116440 228970
rect 116044 228948 116452 228954
rect 116044 228942 116400 228948
rect 116400 228890 116452 228896
rect 115756 228132 115808 228138
rect 115756 228074 115808 228080
rect 115572 227996 115624 228002
rect 115572 227938 115624 227944
rect 117228 225344 117280 225350
rect 117228 225286 117280 225292
rect 116768 224936 116820 224942
rect 116768 224878 116820 224884
rect 115756 224664 115808 224670
rect 115756 224606 115808 224612
rect 114468 220924 114520 220930
rect 114468 220866 114520 220872
rect 113640 218476 113692 218482
rect 113640 218418 113692 218424
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 218418
rect 114480 217274 114508 220866
rect 115768 218074 115796 224606
rect 116780 224126 116808 224878
rect 116768 224120 116820 224126
rect 116768 224062 116820 224068
rect 116952 224120 117004 224126
rect 116952 224062 117004 224068
rect 115296 218068 115348 218074
rect 115296 218010 115348 218016
rect 115756 218068 115808 218074
rect 115756 218010 115808 218016
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 218010
rect 116136 217138 116164 218010
rect 116964 217274 116992 224062
rect 117240 218074 117268 225286
rect 118436 224126 118464 230250
rect 140044 229628 140096 229634
rect 140044 229570 140096 229576
rect 131120 229492 131172 229498
rect 131120 229434 131172 229440
rect 122932 229220 122984 229226
rect 122932 229162 122984 229168
rect 122748 227996 122800 228002
rect 122748 227938 122800 227944
rect 121092 226772 121144 226778
rect 121092 226714 121144 226720
rect 119988 226636 120040 226642
rect 119988 226578 120040 226584
rect 118608 224800 118660 224806
rect 118608 224742 118660 224748
rect 118424 224120 118476 224126
rect 118424 224062 118476 224068
rect 117780 222148 117832 222154
rect 117780 222090 117832 222096
rect 117964 222148 118016 222154
rect 117964 222090 118016 222096
rect 117792 221338 117820 222090
rect 117780 221332 117832 221338
rect 117780 221274 117832 221280
rect 117976 221202 118004 222090
rect 118424 221332 118476 221338
rect 118424 221274 118476 221280
rect 117964 221196 118016 221202
rect 117964 221138 118016 221144
rect 117780 221060 117832 221066
rect 117780 221002 117832 221008
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117792 217274 117820 221002
rect 118436 220930 118464 221274
rect 118424 220924 118476 220930
rect 118424 220866 118476 220872
rect 117964 219428 118016 219434
rect 117964 219370 118016 219376
rect 117976 219162 118004 219370
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 118620 217274 118648 224742
rect 120000 219434 120028 226578
rect 119252 219428 119304 219434
rect 119252 219370 119304 219376
rect 119436 219428 119488 219434
rect 119436 219370 119488 219376
rect 119988 219428 120040 219434
rect 119988 219370 120040 219376
rect 119264 219162 119292 219370
rect 119252 219156 119304 219162
rect 119252 219098 119304 219104
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217246 116992 217274
rect 117746 217246 117820 217274
rect 118574 217246 118648 217274
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217246
rect 117746 216988 117774 217246
rect 118574 216988 118602 217246
rect 119448 217138 119476 219370
rect 119988 218476 120040 218482
rect 119988 218418 120040 218424
rect 120000 218210 120028 218418
rect 119988 218204 120040 218210
rect 119988 218146 120040 218152
rect 120264 218068 120316 218074
rect 120264 218010 120316 218016
rect 120276 217138 120304 218010
rect 121104 217274 121132 226714
rect 121920 224120 121972 224126
rect 121920 224062 121972 224068
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 224062
rect 122760 217274 122788 227938
rect 122944 224942 122972 229162
rect 125784 226908 125836 226914
rect 125784 226850 125836 226856
rect 125796 226506 125824 226850
rect 125784 226500 125836 226506
rect 125784 226442 125836 226448
rect 129372 226500 129424 226506
rect 129372 226442 129424 226448
rect 127440 225480 127492 225486
rect 127440 225422 127492 225428
rect 127452 225214 127480 225422
rect 127440 225208 127492 225214
rect 127440 225150 127492 225156
rect 128268 225208 128320 225214
rect 128268 225150 128320 225156
rect 126888 225072 126940 225078
rect 126888 225014 126940 225020
rect 122932 224936 122984 224942
rect 122932 224878 122984 224884
rect 123484 224936 123536 224942
rect 123484 224878 123536 224884
rect 123496 224398 123524 224878
rect 123484 224392 123536 224398
rect 123484 224334 123536 224340
rect 125232 223848 125284 223854
rect 125232 223790 125284 223796
rect 123390 222864 123446 222873
rect 123390 222799 123446 222808
rect 123404 219162 123432 222799
rect 124404 219836 124456 219842
rect 124404 219778 124456 219784
rect 123392 219156 123444 219162
rect 123392 219098 123444 219104
rect 123576 219156 123628 219162
rect 123576 219098 123628 219104
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 219098
rect 124416 217138 124444 219778
rect 125244 217138 125272 223790
rect 126704 223712 126756 223718
rect 126704 223654 126756 223660
rect 126060 219428 126112 219434
rect 126060 219370 126112 219376
rect 126072 217138 126100 219370
rect 126716 217274 126744 223654
rect 126900 219434 126928 225014
rect 128280 219434 128308 225150
rect 128544 220924 128596 220930
rect 128544 220866 128596 220872
rect 126888 219428 126940 219434
rect 126888 219370 126940 219376
rect 127716 219428 127768 219434
rect 127716 219370 127768 219376
rect 128268 219428 128320 219434
rect 128268 219370 128320 219376
rect 126716 217246 126882 217274
rect 123542 217110 123616 217138
rect 124370 217110 124444 217138
rect 125198 217110 125272 217138
rect 126026 217110 126100 217138
rect 123542 216988 123570 217110
rect 124370 216988 124398 217110
rect 125198 216988 125226 217110
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 219370
rect 128556 217274 128584 220866
rect 128728 219156 128780 219162
rect 128728 219098 128780 219104
rect 128740 218482 128768 219098
rect 128728 218476 128780 218482
rect 128728 218418 128780 218424
rect 129384 217274 129412 226442
rect 131132 223718 131160 229434
rect 140056 229094 140084 229570
rect 139964 229066 140084 229094
rect 133786 227896 133842 227905
rect 133786 227831 133842 227840
rect 134616 227860 134668 227866
rect 131304 224392 131356 224398
rect 131304 224334 131356 224340
rect 131316 224126 131344 224334
rect 131304 224120 131356 224126
rect 131304 224062 131356 224068
rect 131488 224120 131540 224126
rect 131488 224062 131540 224068
rect 131500 223854 131528 224062
rect 131488 223848 131540 223854
rect 131488 223790 131540 223796
rect 131120 223712 131172 223718
rect 131120 223654 131172 223660
rect 132408 223712 132460 223718
rect 132408 223654 132460 223660
rect 131028 219700 131080 219706
rect 131028 219642 131080 219648
rect 130200 219428 130252 219434
rect 130200 219370 130252 219376
rect 127682 217110 127756 217138
rect 128510 217246 128584 217274
rect 129338 217246 129412 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217246
rect 129338 216988 129366 217246
rect 130212 217138 130240 219370
rect 131040 217274 131068 219642
rect 132420 219162 132448 223654
rect 133512 222488 133564 222494
rect 133512 222430 133564 222436
rect 132684 219428 132736 219434
rect 132684 219370 132736 219376
rect 131856 219156 131908 219162
rect 131856 219098 131908 219104
rect 132408 219156 132460 219162
rect 132408 219098 132460 219104
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219098
rect 132696 217138 132724 219370
rect 133524 217274 133552 222430
rect 133800 219434 133828 227831
rect 134616 227802 134668 227808
rect 134432 223848 134484 223854
rect 134432 223790 134484 223796
rect 133788 219428 133840 219434
rect 133788 219370 133840 219376
rect 134444 219026 134472 223790
rect 134432 219020 134484 219026
rect 134432 218962 134484 218968
rect 134628 217274 134656 227802
rect 135260 227044 135312 227050
rect 135260 226986 135312 226992
rect 135444 227044 135496 227050
rect 135444 226986 135496 226992
rect 135272 226522 135300 226986
rect 135456 226642 135484 226986
rect 135444 226636 135496 226642
rect 135444 226578 135496 226584
rect 135628 226636 135680 226642
rect 135628 226578 135680 226584
rect 137560 226636 137612 226642
rect 137560 226578 137612 226584
rect 135640 226522 135668 226578
rect 137572 226522 137600 226578
rect 135272 226494 135668 226522
rect 137204 226506 137600 226522
rect 137192 226500 137600 226506
rect 137244 226494 137600 226500
rect 139306 226536 139362 226545
rect 139306 226471 139362 226480
rect 137192 226442 137244 226448
rect 136824 225616 136876 225622
rect 136824 225558 136876 225564
rect 137008 225616 137060 225622
rect 137008 225558 137060 225564
rect 136546 225312 136602 225321
rect 136546 225247 136602 225256
rect 136560 219026 136588 225247
rect 136836 225162 136864 225558
rect 137020 225350 137048 225558
rect 137008 225344 137060 225350
rect 137008 225286 137060 225292
rect 136836 225134 137508 225162
rect 137480 225078 137508 225134
rect 137468 225072 137520 225078
rect 137468 225014 137520 225020
rect 138294 221776 138350 221785
rect 138294 221711 138350 221720
rect 137284 221604 137336 221610
rect 137284 221546 137336 221552
rect 137468 221604 137520 221610
rect 137468 221546 137520 221552
rect 137296 221202 137324 221546
rect 137100 221196 137152 221202
rect 137100 221138 137152 221144
rect 137284 221196 137336 221202
rect 137284 221138 137336 221144
rect 137112 221082 137140 221138
rect 137480 221082 137508 221546
rect 138308 221474 138336 221711
rect 138296 221468 138348 221474
rect 138296 221410 138348 221416
rect 138480 221468 138532 221474
rect 138480 221410 138532 221416
rect 137112 221054 137508 221082
rect 137284 220788 137336 220794
rect 137284 220730 137336 220736
rect 137468 220788 137520 220794
rect 137468 220730 137520 220736
rect 137296 219706 137324 220730
rect 137284 219700 137336 219706
rect 137284 219642 137336 219648
rect 137480 219570 137508 220730
rect 137468 219564 137520 219570
rect 137468 219506 137520 219512
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 135076 219020 135128 219026
rect 135076 218962 135128 218968
rect 135996 219020 136048 219026
rect 135996 218962 136048 218968
rect 136548 219020 136600 219026
rect 136548 218962 136600 218968
rect 136824 219020 136876 219026
rect 136824 218962 136876 218968
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133552 217274
rect 134306 217246 134656 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135088 217138 135116 218962
rect 136008 217138 136036 218962
rect 136836 217138 136864 218962
rect 137664 217274 137692 219506
rect 137834 219192 137890 219201
rect 137834 219127 137890 219136
rect 138110 219192 138166 219201
rect 138110 219127 138112 219136
rect 137848 219026 137876 219127
rect 138164 219127 138166 219136
rect 138112 219098 138164 219104
rect 137836 219020 137888 219026
rect 137836 218962 137888 218968
rect 135088 217110 135162 217138
rect 135134 216988 135162 217110
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 221410
rect 139320 217274 139348 226471
rect 139964 219026 139992 229066
rect 140792 228546 140820 231662
rect 140780 228540 140832 228546
rect 140780 228482 140832 228488
rect 140964 228540 141016 228546
rect 140964 228482 141016 228488
rect 140976 228138 141004 228482
rect 140964 228132 141016 228138
rect 140964 228074 141016 228080
rect 141148 228132 141200 228138
rect 141148 228074 141200 228080
rect 141160 227866 141188 228074
rect 141330 227896 141386 227905
rect 141148 227860 141200 227866
rect 141330 227831 141332 227840
rect 141148 227802 141200 227808
rect 141384 227831 141386 227840
rect 141332 227802 141384 227808
rect 141528 225078 141556 231662
rect 142158 227216 142214 227225
rect 142158 227151 142214 227160
rect 142172 226658 142200 227151
rect 142126 226630 142200 226658
rect 142126 226506 142154 226630
rect 142250 226536 142306 226545
rect 142114 226500 142166 226506
rect 142250 226471 142252 226480
rect 142114 226442 142166 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 142114 225344 142166 225350
rect 142252 225344 142304 225350
rect 142114 225286 142166 225292
rect 142250 225312 142252 225321
rect 142304 225312 142306 225321
rect 142126 225162 142154 225286
rect 142250 225247 142306 225256
rect 142448 225162 142476 231676
rect 143092 227225 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 145038 231662 145236 231690
rect 143078 227216 143134 227225
rect 143078 227151 143134 227160
rect 143552 226166 143580 231662
rect 143540 226160 143592 226166
rect 143540 226102 143592 226108
rect 143170 225584 143226 225593
rect 143170 225519 143226 225528
rect 142126 225134 142200 225162
rect 142448 225134 142660 225162
rect 141516 225072 141568 225078
rect 141516 225014 141568 225020
rect 141792 225072 141844 225078
rect 142172 225060 142200 225134
rect 142436 225072 142488 225078
rect 142172 225032 142436 225060
rect 141792 225014 141844 225020
rect 142436 225014 142488 225020
rect 140964 223984 141016 223990
rect 140962 223952 140964 223961
rect 141016 223952 141018 223961
rect 140962 223887 141018 223896
rect 140778 220144 140834 220153
rect 140778 220079 140780 220088
rect 140832 220079 140834 220088
rect 140964 220108 141016 220114
rect 140780 220050 140832 220056
rect 140964 220050 141016 220056
rect 139952 219020 140004 219026
rect 139952 218962 140004 218968
rect 140136 219020 140188 219026
rect 140136 218962 140188 218968
rect 140148 218770 140176 218962
rect 139964 218742 140176 218770
rect 139964 218618 139992 218742
rect 139952 218612 140004 218618
rect 139952 218554 140004 218560
rect 140136 218612 140188 218618
rect 140136 218554 140188 218560
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218554
rect 140976 217138 141004 220050
rect 141804 217274 141832 225014
rect 142068 224936 142120 224942
rect 142068 224878 142120 224884
rect 142080 223990 142108 224878
rect 142068 223984 142120 223990
rect 142068 223926 142120 223932
rect 142632 222358 142660 225134
rect 142620 222352 142672 222358
rect 142620 222294 142672 222300
rect 142804 221876 142856 221882
rect 142804 221818 142856 221824
rect 142988 221876 143040 221882
rect 142988 221818 143040 221824
rect 142816 221610 142844 221818
rect 142804 221604 142856 221610
rect 142804 221546 142856 221552
rect 143000 221474 143028 221818
rect 142436 221468 142488 221474
rect 142436 221410 142488 221416
rect 142988 221468 143040 221474
rect 142988 221410 143040 221416
rect 142448 221241 142476 221410
rect 142434 221232 142490 221241
rect 142434 221167 142490 221176
rect 143184 219434 143212 225519
rect 143448 222284 143500 222290
rect 143448 222226 143500 222232
rect 142436 219428 142488 219434
rect 142436 219370 142488 219376
rect 142620 219428 142672 219434
rect 142620 219370 142672 219376
rect 143172 219428 143224 219434
rect 143172 219370 143224 219376
rect 142250 219056 142306 219065
rect 142448 219026 142476 219370
rect 142250 218991 142252 219000
rect 142304 218991 142306 219000
rect 142436 219020 142488 219026
rect 142252 218962 142304 218968
rect 142436 218962 142488 218968
rect 140102 217110 140176 217138
rect 140930 217110 141004 217138
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217110
rect 141758 216988 141786 217246
rect 142632 217138 142660 219370
rect 143460 217138 143488 222226
rect 144012 221202 144040 231662
rect 144644 230580 144696 230586
rect 144644 230522 144696 230528
rect 144656 229770 144684 230522
rect 144644 229764 144696 229770
rect 144644 229706 144696 229712
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 222290 144868 229706
rect 145208 224262 145236 231662
rect 145668 229809 145696 231676
rect 146326 231662 146524 231690
rect 145654 229800 145710 229809
rect 145654 229735 145710 229744
rect 146298 229392 146354 229401
rect 146298 229327 146300 229336
rect 146352 229327 146354 229336
rect 146300 229298 146352 229304
rect 145930 225312 145986 225321
rect 145930 225247 145986 225256
rect 145196 224256 145248 224262
rect 145196 224198 145248 224204
rect 145380 224256 145432 224262
rect 145380 224198 145432 224204
rect 145392 223961 145420 224198
rect 145654 224088 145710 224097
rect 145654 224023 145710 224032
rect 145378 223952 145434 223961
rect 145378 223887 145434 223896
rect 145012 222352 145064 222358
rect 145012 222294 145064 222300
rect 144828 222284 144880 222290
rect 144828 222226 144880 222232
rect 145024 222170 145052 222294
rect 144840 222142 145052 222170
rect 144182 221232 144238 221241
rect 144000 221196 144052 221202
rect 144182 221167 144184 221176
rect 144000 221138 144052 221144
rect 144236 221167 144238 221176
rect 144184 221138 144236 221144
rect 143632 219428 143684 219434
rect 143632 219370 143684 219376
rect 143644 219162 143672 219370
rect 143632 219156 143684 219162
rect 143632 219098 143684 219104
rect 143816 219156 143868 219162
rect 143816 219098 143868 219104
rect 143828 218618 143856 219098
rect 144840 218618 144868 222142
rect 145668 219065 145696 224023
rect 145654 219056 145710 219065
rect 145654 218991 145710 219000
rect 143816 218612 143868 218618
rect 143816 218554 143868 218560
rect 144276 218612 144328 218618
rect 144276 218554 144328 218560
rect 144828 218612 144880 218618
rect 144828 218554 144880 218560
rect 144288 217138 144316 218554
rect 145944 217274 145972 225247
rect 146496 224954 146524 231662
rect 146680 231662 146970 231690
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 148428 231662 148902 231690
rect 149072 231662 149546 231690
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 151096 231662 151478 231690
rect 151740 231662 152122 231690
rect 152476 231662 152766 231690
rect 146680 229094 146708 231662
rect 146944 229628 146996 229634
rect 146944 229570 146996 229576
rect 146956 229362 146984 229570
rect 146944 229356 146996 229362
rect 146944 229298 146996 229304
rect 146404 224926 146524 224954
rect 146588 229066 146708 229094
rect 146404 220153 146432 224926
rect 146588 221785 146616 229066
rect 147034 225992 147090 226001
rect 147034 225927 147090 225936
rect 147048 225622 147076 225927
rect 147036 225616 147088 225622
rect 147036 225558 147088 225564
rect 147232 224262 147260 231662
rect 147968 229401 147996 231662
rect 147954 229392 148010 229401
rect 147954 229327 148010 229336
rect 147678 228576 147734 228585
rect 147678 228511 147734 228520
rect 147692 228426 147720 228511
rect 147646 228410 147720 228426
rect 147634 228404 147720 228410
rect 147686 228398 147720 228404
rect 147634 228346 147686 228352
rect 147404 225616 147456 225622
rect 147402 225584 147404 225593
rect 147456 225584 147458 225593
rect 147402 225519 147458 225528
rect 148428 224954 148456 231662
rect 148600 229764 148652 229770
rect 148600 229706 148652 229712
rect 148244 224926 148456 224954
rect 147220 224256 147272 224262
rect 147220 224198 147272 224204
rect 147772 224256 147824 224262
rect 147772 224198 147824 224204
rect 147784 224097 147812 224198
rect 147770 224088 147826 224097
rect 147770 224023 147826 224032
rect 147310 222184 147366 222193
rect 147310 222119 147366 222128
rect 146574 221776 146630 221785
rect 146574 221711 146630 221720
rect 147324 221610 147352 222119
rect 147494 221912 147550 221921
rect 147494 221847 147550 221856
rect 147508 221746 147536 221847
rect 147496 221740 147548 221746
rect 147496 221682 147548 221688
rect 147772 221740 147824 221746
rect 147772 221682 147824 221688
rect 147312 221604 147364 221610
rect 147312 221546 147364 221552
rect 147494 220280 147550 220289
rect 147494 220215 147496 220224
rect 147548 220215 147550 220224
rect 147634 220244 147686 220250
rect 147496 220186 147548 220192
rect 147634 220186 147686 220192
rect 146390 220144 146446 220153
rect 147646 220130 147674 220186
rect 146390 220079 146446 220088
rect 147036 220108 147088 220114
rect 147036 220050 147088 220056
rect 147508 220102 147674 220130
rect 147048 219473 147076 220050
rect 147508 219706 147536 220102
rect 147496 219700 147548 219706
rect 147496 219642 147548 219648
rect 147034 219464 147090 219473
rect 147034 219399 147090 219408
rect 147494 218784 147550 218793
rect 147494 218719 147496 218728
rect 147548 218719 147550 218728
rect 147496 218690 147548 218696
rect 146760 218612 146812 218618
rect 146760 218554 146812 218560
rect 145058 217252 145110 217258
rect 145058 217194 145110 217200
rect 145898 217246 145972 217274
rect 142586 217110 142660 217138
rect 143414 217110 143488 217138
rect 144242 217110 144316 217138
rect 142586 216988 142614 217110
rect 143414 216988 143442 217110
rect 144242 216988 144270 217110
rect 145070 216988 145098 217194
rect 145898 216988 145926 217246
rect 146772 217138 146800 218554
rect 147784 217258 147812 221682
rect 148244 220289 148272 224926
rect 148416 221468 148468 221474
rect 148416 221410 148468 221416
rect 148230 220280 148286 220289
rect 148230 220215 148286 220224
rect 148048 219700 148100 219706
rect 148048 219642 148100 219648
rect 148060 219473 148088 219642
rect 148046 219464 148102 219473
rect 148046 219399 148102 219408
rect 147772 217252 147824 217258
rect 147772 217194 147824 217200
rect 148428 217138 148456 221410
rect 148612 218793 148640 229706
rect 149072 221921 149100 231662
rect 149808 228585 149836 231662
rect 150544 230586 150572 231662
rect 150532 230580 150584 230586
rect 150532 230522 150584 230528
rect 150900 230580 150952 230586
rect 150900 230522 150952 230528
rect 150912 229770 150940 230522
rect 150900 229764 150952 229770
rect 150900 229706 150952 229712
rect 149794 228576 149850 228585
rect 149794 228511 149850 228520
rect 150162 227216 150218 227225
rect 150162 227151 150164 227160
rect 150216 227151 150218 227160
rect 150348 227180 150400 227186
rect 150164 227122 150216 227128
rect 150348 227122 150400 227128
rect 149058 221912 149114 221921
rect 149058 221847 149114 221856
rect 150070 220824 150126 220833
rect 150070 220759 150126 220768
rect 150084 220402 150112 220759
rect 150038 220386 150112 220402
rect 150026 220380 150112 220386
rect 150078 220374 150112 220380
rect 150026 220322 150078 220328
rect 148598 218784 148654 218793
rect 148598 218719 148654 218728
rect 149060 218612 149112 218618
rect 149060 218554 149112 218560
rect 149072 218346 149100 218554
rect 150360 218346 150388 227122
rect 150900 220380 150952 220386
rect 150900 220322 150952 220328
rect 150716 220108 150768 220114
rect 150716 220050 150768 220056
rect 149060 218340 149112 218346
rect 149060 218282 149112 218288
rect 149244 218340 149296 218346
rect 149244 218282 149296 218288
rect 150348 218340 150400 218346
rect 150348 218282 150400 218288
rect 150532 218340 150584 218346
rect 150532 218282 150584 218288
rect 149256 217138 149284 218282
rect 150544 218226 150572 218282
rect 150084 218198 150572 218226
rect 150084 217274 150112 218198
rect 146726 217110 146800 217138
rect 147542 217116 147594 217122
rect 146726 216988 146754 217110
rect 147542 217058 147594 217064
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150112 217274
rect 147554 216988 147582 217058
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150728 217122 150756 220050
rect 150912 217138 150940 220322
rect 151096 219881 151124 231662
rect 151360 229764 151412 229770
rect 151360 229706 151412 229712
rect 151372 222494 151400 229706
rect 151740 226930 151768 231662
rect 151910 227488 151966 227497
rect 151910 227423 151966 227432
rect 151924 227322 151952 227423
rect 151912 227316 151964 227322
rect 151912 227258 151964 227264
rect 152280 227180 152332 227186
rect 151924 227140 152280 227168
rect 151924 227050 151952 227140
rect 152280 227122 152332 227128
rect 151912 227044 151964 227050
rect 151912 226986 151964 226992
rect 151740 226902 152136 226930
rect 151726 223816 151782 223825
rect 151726 223751 151782 223760
rect 151360 222488 151412 222494
rect 151360 222430 151412 222436
rect 151082 219872 151138 219881
rect 151082 219807 151138 219816
rect 151740 217138 151768 223751
rect 152108 222193 152136 226902
rect 152476 224369 152504 231662
rect 153396 229362 153424 231676
rect 153672 231662 154054 231690
rect 154592 231662 154698 231690
rect 153384 229356 153436 229362
rect 153384 229298 153436 229304
rect 153292 228540 153344 228546
rect 153292 228482 153344 228488
rect 152922 227488 152978 227497
rect 152922 227423 152978 227432
rect 152936 227322 152964 227423
rect 152924 227316 152976 227322
rect 152924 227258 152976 227264
rect 152832 226296 152884 226302
rect 152832 226238 152884 226244
rect 152844 226001 152872 226238
rect 153106 226128 153162 226137
rect 153106 226063 153162 226072
rect 152830 225992 152886 226001
rect 152830 225927 152886 225936
rect 152462 224360 152518 224369
rect 152462 224295 152518 224304
rect 152094 222184 152150 222193
rect 152094 222119 152150 222128
rect 152648 220516 152700 220522
rect 152648 220458 152700 220464
rect 152280 220380 152332 220386
rect 152280 220322 152332 220328
rect 152292 220130 152320 220322
rect 152660 220250 152688 220458
rect 152648 220244 152700 220250
rect 152648 220186 152700 220192
rect 152832 220244 152884 220250
rect 152832 220186 152884 220192
rect 152844 220130 152872 220186
rect 152292 220102 152872 220130
rect 152384 219422 152780 219450
rect 152384 219298 152412 219422
rect 152752 219314 152780 219422
rect 152372 219292 152424 219298
rect 152372 219234 152424 219240
rect 152556 219292 152608 219298
rect 152752 219286 152964 219314
rect 153120 219298 153148 226063
rect 153304 225321 153332 228482
rect 153290 225312 153346 225321
rect 153290 225247 153346 225256
rect 153672 220561 153700 231662
rect 153844 229356 153896 229362
rect 153844 229298 153896 229304
rect 153658 220552 153714 220561
rect 153658 220487 153714 220496
rect 152556 219234 152608 219240
rect 152280 219156 152332 219162
rect 152280 219098 152332 219104
rect 152094 218920 152150 218929
rect 152292 218890 152320 219098
rect 152094 218855 152096 218864
rect 152148 218855 152150 218864
rect 152280 218884 152332 218890
rect 152096 218826 152148 218832
rect 152280 218826 152332 218832
rect 152568 217138 152596 219234
rect 152740 219020 152792 219026
rect 152740 218962 152792 218968
rect 152752 218754 152780 218962
rect 152936 218754 152964 219286
rect 153108 219292 153160 219298
rect 153108 219234 153160 219240
rect 153384 219292 153436 219298
rect 153384 219234 153436 219240
rect 152740 218748 152792 218754
rect 152740 218690 152792 218696
rect 152924 218748 152976 218754
rect 152924 218690 152976 218696
rect 153396 217138 153424 219234
rect 153856 218929 153884 229298
rect 154592 227225 154620 231662
rect 154578 227216 154634 227225
rect 154578 227151 154634 227160
rect 155328 226953 155356 231676
rect 155972 229906 156000 231676
rect 156156 231662 156630 231690
rect 155960 229900 156012 229906
rect 155960 229842 156012 229848
rect 155866 228032 155922 228041
rect 155866 227967 155922 227976
rect 155314 226944 155370 226953
rect 155314 226879 155370 226888
rect 155038 223136 155094 223145
rect 155038 223071 155094 223080
rect 154212 222488 154264 222494
rect 154212 222430 154264 222436
rect 153842 218920 153898 218929
rect 153842 218855 153898 218864
rect 154224 217138 154252 222430
rect 155052 217138 155080 223071
rect 155880 217274 155908 227967
rect 156156 220833 156184 231662
rect 156328 229900 156380 229906
rect 156328 229842 156380 229848
rect 156142 220824 156198 220833
rect 156142 220759 156198 220768
rect 156340 218754 156368 229842
rect 157260 224954 157288 231676
rect 157628 231662 157918 231690
rect 158272 231662 158562 231690
rect 158824 231662 159206 231690
rect 157430 228576 157486 228585
rect 157430 228511 157486 228520
rect 157444 228410 157472 228511
rect 157432 228404 157484 228410
rect 157432 228346 157484 228352
rect 157628 226250 157656 231662
rect 158272 230722 158300 231662
rect 158260 230716 158312 230722
rect 158260 230658 158312 230664
rect 157982 229392 158038 229401
rect 157982 229327 158038 229336
rect 157800 228404 157852 228410
rect 157800 228346 157852 228352
rect 157812 228041 157840 228346
rect 157798 228032 157854 228041
rect 157798 227967 157854 227976
rect 157444 226222 157656 226250
rect 157444 226166 157472 226222
rect 157432 226160 157484 226166
rect 157616 226160 157668 226166
rect 157432 226102 157484 226108
rect 157614 226128 157616 226137
rect 157668 226128 157670 226137
rect 157614 226063 157670 226072
rect 156892 224926 157288 224954
rect 156696 224256 156748 224262
rect 156696 224198 156748 224204
rect 156708 224097 156736 224198
rect 156694 224088 156750 224097
rect 156694 224023 156750 224032
rect 156892 223174 156920 224926
rect 157062 224360 157118 224369
rect 157062 224295 157118 224304
rect 157076 223990 157104 224295
rect 157432 224256 157484 224262
rect 157432 224198 157484 224204
rect 157444 224097 157472 224198
rect 157430 224088 157486 224097
rect 157430 224023 157486 224032
rect 157064 223984 157116 223990
rect 157064 223926 157116 223932
rect 157248 223984 157300 223990
rect 157248 223926 157300 223932
rect 157260 223825 157288 223926
rect 157246 223816 157302 223825
rect 157246 223751 157302 223760
rect 157248 223440 157300 223446
rect 157246 223408 157248 223417
rect 157432 223440 157484 223446
rect 157300 223408 157302 223417
rect 157246 223343 157302 223352
rect 157430 223408 157432 223417
rect 157484 223408 157486 223417
rect 157430 223343 157486 223352
rect 156880 223168 156932 223174
rect 157064 223168 157116 223174
rect 156880 223110 156932 223116
rect 157062 223136 157064 223145
rect 157116 223136 157118 223145
rect 157062 223071 157118 223080
rect 157338 220416 157394 220425
rect 157338 220351 157340 220360
rect 157392 220351 157394 220360
rect 157524 220380 157576 220386
rect 157340 220322 157392 220328
rect 157524 220322 157576 220328
rect 156328 218748 156380 218754
rect 156328 218690 156380 218696
rect 156696 218748 156748 218754
rect 156696 218690 156748 218696
rect 150716 217116 150768 217122
rect 150716 217058 150768 217064
rect 150866 217110 150940 217138
rect 151694 217110 151768 217138
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217110 154252 217138
rect 155006 217110 155080 217138
rect 155834 217246 155908 217274
rect 150866 216988 150894 217110
rect 151694 216988 151722 217110
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217110
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218690
rect 157246 218648 157302 218657
rect 157246 218583 157302 218592
rect 157260 218346 157288 218583
rect 157248 218340 157300 218346
rect 157248 218282 157300 218288
rect 157536 217138 157564 220322
rect 157706 218648 157762 218657
rect 157996 218618 158024 229327
rect 158824 228585 158852 231662
rect 158810 228576 158866 228585
rect 158810 228511 158866 228520
rect 159638 227488 159694 227497
rect 159638 227423 159640 227432
rect 159692 227423 159694 227432
rect 159640 227394 159692 227400
rect 159836 223446 159864 231676
rect 160480 228313 160508 231676
rect 161124 230450 161152 231676
rect 161112 230444 161164 230450
rect 161112 230386 161164 230392
rect 161296 230444 161348 230450
rect 161296 230386 161348 230392
rect 160466 228304 160522 228313
rect 160466 228239 160522 228248
rect 160008 227452 160060 227458
rect 160008 227394 160060 227400
rect 159824 223440 159876 223446
rect 159824 223382 159876 223388
rect 158350 223136 158406 223145
rect 158350 223071 158406 223080
rect 157706 218583 157762 218592
rect 157984 218612 158036 218618
rect 157720 218210 157748 218583
rect 157984 218554 158036 218560
rect 157708 218204 157760 218210
rect 157708 218146 157760 218152
rect 158364 217138 158392 223071
rect 160020 219298 160048 227394
rect 160834 222592 160890 222601
rect 160834 222527 160890 222536
rect 158996 219292 159048 219298
rect 158996 219234 159048 219240
rect 159180 219292 159232 219298
rect 159180 219234 159232 219240
rect 160008 219292 160060 219298
rect 160008 219234 160060 219240
rect 160192 219292 160244 219298
rect 160192 219234 160244 219240
rect 159008 218618 159036 219234
rect 158996 218612 159048 218618
rect 158996 218554 159048 218560
rect 159192 217138 159220 219234
rect 160204 218770 160232 219234
rect 159836 218742 160232 218770
rect 159836 218346 159864 218742
rect 159824 218340 159876 218346
rect 159824 218282 159876 218288
rect 160008 218340 160060 218346
rect 160008 218282 160060 218288
rect 160020 217138 160048 218282
rect 160848 217138 160876 222527
rect 161308 218210 161336 230386
rect 161572 226024 161624 226030
rect 161572 225966 161624 225972
rect 161584 225593 161612 225966
rect 161570 225584 161626 225593
rect 161570 225519 161626 225528
rect 161768 224954 161796 231676
rect 162136 231662 162426 231690
rect 162964 231662 163070 231690
rect 161940 226296 161992 226302
rect 161940 226238 161992 226244
rect 161952 226030 161980 226238
rect 161940 226024 161992 226030
rect 161940 225966 161992 225972
rect 162136 224954 162164 231662
rect 162308 226296 162360 226302
rect 162308 226238 162360 226244
rect 162320 225078 162348 226238
rect 162308 225072 162360 225078
rect 162308 225014 162360 225020
rect 162492 225072 162544 225078
rect 162492 225014 162544 225020
rect 161492 224926 161796 224954
rect 161860 224926 162164 224954
rect 161492 220425 161520 224926
rect 161860 223666 161888 224926
rect 161768 223638 161888 223666
rect 161768 222766 161796 223638
rect 161940 223576 161992 223582
rect 161940 223518 161992 223524
rect 161952 223038 161980 223518
rect 162124 223168 162176 223174
rect 162124 223110 162176 223116
rect 161940 223032 161992 223038
rect 161940 222974 161992 222980
rect 162136 222766 162164 223110
rect 162308 222896 162360 222902
rect 162308 222838 162360 222844
rect 161756 222760 161808 222766
rect 161756 222702 161808 222708
rect 162124 222760 162176 222766
rect 162124 222702 162176 222708
rect 162320 222601 162348 222838
rect 162306 222592 162362 222601
rect 162306 222527 162362 222536
rect 161664 221740 161716 221746
rect 161664 221682 161716 221688
rect 161478 220416 161534 220425
rect 161478 220351 161534 220360
rect 161296 218204 161348 218210
rect 161296 218146 161348 218152
rect 161676 217138 161704 221682
rect 162124 218748 162176 218754
rect 162124 218690 162176 218696
rect 162136 218210 162164 218690
rect 162124 218204 162176 218210
rect 162124 218146 162176 218152
rect 162504 217274 162532 225014
rect 162964 224369 162992 231662
rect 163700 229362 163728 231676
rect 163870 229392 163926 229401
rect 163688 229356 163740 229362
rect 163870 229327 163872 229336
rect 163688 229298 163740 229304
rect 163924 229327 163926 229336
rect 163872 229298 163924 229304
rect 164344 227322 164372 231676
rect 164332 227316 164384 227322
rect 164332 227258 164384 227264
rect 162950 224360 163006 224369
rect 162950 224295 163006 224304
rect 163962 223952 164018 223961
rect 163962 223887 164018 223896
rect 163976 219298 164004 223887
rect 164988 223446 165016 231676
rect 165436 227316 165488 227322
rect 165436 227258 165488 227264
rect 164976 223440 165028 223446
rect 164976 223382 165028 223388
rect 165252 223440 165304 223446
rect 165252 223382 165304 223388
rect 165264 223174 165292 223382
rect 164148 223168 164200 223174
rect 164148 223110 164200 223116
rect 165252 223168 165304 223174
rect 165252 223110 165304 223116
rect 163964 219292 164016 219298
rect 163964 219234 164016 219240
rect 162676 218612 162728 218618
rect 162676 218554 162728 218560
rect 162688 218346 162716 218554
rect 162676 218340 162728 218346
rect 162676 218282 162728 218288
rect 162860 218340 162912 218346
rect 162860 218282 162912 218288
rect 162872 218074 162900 218282
rect 162860 218068 162912 218074
rect 162860 218010 162912 218016
rect 163320 218068 163372 218074
rect 163320 218010 163372 218016
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217110 158392 217138
rect 159146 217110 159220 217138
rect 159974 217110 160048 217138
rect 160802 217110 160876 217138
rect 161630 217110 161704 217138
rect 162458 217246 162532 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217110
rect 159146 216988 159174 217110
rect 159974 216988 160002 217110
rect 160802 216988 160830 217110
rect 161630 216988 161658 217110
rect 162458 216988 162486 217246
rect 163332 217138 163360 218010
rect 164160 217138 164188 223110
rect 165448 219298 165476 227258
rect 165632 222873 165660 231676
rect 166276 230042 166304 231676
rect 166460 231662 166934 231690
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 166264 230036 166316 230042
rect 166264 229978 166316 229984
rect 166460 227497 166488 231662
rect 166632 230036 166684 230042
rect 166632 229978 166684 229984
rect 166644 229362 166672 229978
rect 166632 229356 166684 229362
rect 166632 229298 166684 229304
rect 166630 228440 166686 228449
rect 166630 228375 166686 228384
rect 166446 227488 166502 227497
rect 166446 227423 166502 227432
rect 166644 225706 166672 228375
rect 166908 227452 166960 227458
rect 166908 227394 166960 227400
rect 166920 226386 166948 227394
rect 166920 226370 166994 226386
rect 166920 226364 167006 226370
rect 166920 226358 166954 226364
rect 166954 226306 167006 226312
rect 166816 226296 166868 226302
rect 166816 226238 166868 226244
rect 166828 225978 166856 226238
rect 166828 225950 166994 225978
rect 166966 225894 166994 225950
rect 166816 225888 166868 225894
rect 166814 225856 166816 225865
rect 166954 225888 167006 225894
rect 166868 225856 166870 225865
rect 166954 225830 167006 225836
rect 166814 225791 166870 225800
rect 166644 225678 166948 225706
rect 166722 225584 166778 225593
rect 166722 225519 166778 225528
rect 166736 225078 166764 225519
rect 166540 225072 166592 225078
rect 166538 225040 166540 225049
rect 166724 225072 166776 225078
rect 166592 225040 166594 225049
rect 166724 225014 166776 225020
rect 166538 224975 166594 224984
rect 166920 224954 166948 225678
rect 166736 224926 166948 224954
rect 166736 223394 166764 224926
rect 166552 223366 166764 223394
rect 165804 223168 165856 223174
rect 165802 223136 165804 223145
rect 165856 223136 165858 223145
rect 165802 223071 165858 223080
rect 165618 222864 165674 222873
rect 165618 222799 165674 222808
rect 166552 219298 166580 223366
rect 166816 223304 166868 223310
rect 166814 223272 166816 223281
rect 166954 223304 167006 223310
rect 166868 223272 166870 223281
rect 166954 223246 167006 223252
rect 166814 223207 166870 223216
rect 166966 223122 166994 223246
rect 166828 223094 166994 223122
rect 164976 219292 165028 219298
rect 164976 219234 165028 219240
rect 165436 219292 165488 219298
rect 165436 219234 165488 219240
rect 165804 219292 165856 219298
rect 165804 219234 165856 219240
rect 166540 219292 166592 219298
rect 166540 219234 166592 219240
rect 164988 217138 165016 219234
rect 165816 217138 165844 219234
rect 166262 219192 166318 219201
rect 166262 219127 166318 219136
rect 166276 219026 166304 219127
rect 166264 219020 166316 219026
rect 166264 218962 166316 218968
rect 166446 218920 166502 218929
rect 166446 218855 166448 218864
rect 166500 218855 166502 218864
rect 166448 218826 166500 218832
rect 166264 218748 166316 218754
rect 166264 218690 166316 218696
rect 166276 218385 166304 218690
rect 166538 218648 166594 218657
rect 166538 218583 166540 218592
rect 166592 218583 166594 218592
rect 166540 218554 166592 218560
rect 166828 218498 166856 223094
rect 167196 220522 167224 231662
rect 167644 229356 167696 229362
rect 167644 229298 167696 229304
rect 167184 220516 167236 220522
rect 167184 220458 167236 220464
rect 167182 219192 167238 219201
rect 167000 219156 167052 219162
rect 167182 219127 167238 219136
rect 167000 219098 167052 219104
rect 167012 218929 167040 219098
rect 167196 219026 167224 219127
rect 167184 219020 167236 219026
rect 167184 218962 167236 218968
rect 166998 218920 167054 218929
rect 166998 218855 167054 218864
rect 167184 218884 167236 218890
rect 167184 218826 167236 218832
rect 167196 218657 167224 218826
rect 167368 218748 167420 218754
rect 167368 218690 167420 218696
rect 167182 218648 167238 218657
rect 167182 218583 167238 218592
rect 166460 218470 166856 218498
rect 166262 218376 166318 218385
rect 166460 218346 166488 218470
rect 167380 218385 167408 218690
rect 167366 218376 167422 218385
rect 166262 218311 166318 218320
rect 166448 218340 166500 218346
rect 166448 218282 166500 218288
rect 166632 218340 166684 218346
rect 167366 218311 167422 218320
rect 166632 218282 166684 218288
rect 166644 217138 166672 218282
rect 167656 218210 167684 229298
rect 167840 223582 167868 231662
rect 168852 227186 168880 231676
rect 169036 231662 169510 231690
rect 169864 231662 170154 231690
rect 170416 231662 170798 231690
rect 171152 231662 171442 231690
rect 168840 227180 168892 227186
rect 168840 227122 168892 227128
rect 169036 225078 169064 231662
rect 169576 227180 169628 227186
rect 169576 227122 169628 227128
rect 169024 225072 169076 225078
rect 169024 225014 169076 225020
rect 169208 225072 169260 225078
rect 169208 225014 169260 225020
rect 167828 223576 167880 223582
rect 167828 223518 167880 223524
rect 168288 223576 168340 223582
rect 168288 223518 168340 223524
rect 167644 218204 167696 218210
rect 167644 218146 167696 218152
rect 168104 218204 168156 218210
rect 168104 218146 168156 218152
rect 167460 218068 167512 218074
rect 167460 218010 167512 218016
rect 167472 217138 167500 218010
rect 168116 217274 168144 218146
rect 168300 218074 168328 223518
rect 169220 219434 169248 225014
rect 168944 219406 169248 219434
rect 168944 219298 168972 219406
rect 168932 219292 168984 219298
rect 168932 219234 168984 219240
rect 169300 219292 169352 219298
rect 169300 219234 169352 219240
rect 168288 218068 168340 218074
rect 168288 218010 168340 218016
rect 169116 218068 169168 218074
rect 169116 218010 169168 218016
rect 168116 217246 168282 217274
rect 163286 217110 163360 217138
rect 164114 217110 164188 217138
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 163286 216988 163314 217110
rect 164114 216988 164142 217110
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 218010
rect 169312 217938 169340 219234
rect 169588 218074 169616 227122
rect 169864 225865 169892 231662
rect 169850 225856 169906 225865
rect 169850 225791 169906 225800
rect 170416 223281 170444 231662
rect 171152 229094 171180 231662
rect 171152 229066 171456 229094
rect 171138 228712 171194 228721
rect 171138 228647 171194 228656
rect 171152 228562 171180 228647
rect 171060 228534 171180 228562
rect 171060 228274 171088 228534
rect 171230 228440 171286 228449
rect 171230 228375 171286 228384
rect 171244 228274 171272 228375
rect 171048 228268 171100 228274
rect 171048 228210 171100 228216
rect 171232 228268 171284 228274
rect 171232 228210 171284 228216
rect 171048 226024 171100 226030
rect 170862 225992 170918 226001
rect 171232 226024 171284 226030
rect 171048 225966 171100 225972
rect 171230 225992 171232 226001
rect 171284 225992 171286 226001
rect 170862 225927 170918 225936
rect 170876 225078 170904 225927
rect 171060 225842 171088 225966
rect 171230 225927 171286 225936
rect 171060 225814 171272 225842
rect 171244 225758 171272 225814
rect 171048 225752 171100 225758
rect 171046 225720 171048 225729
rect 171232 225752 171284 225758
rect 171100 225720 171102 225729
rect 171232 225694 171284 225700
rect 171046 225655 171102 225664
rect 170864 225072 170916 225078
rect 171048 225072 171100 225078
rect 170864 225014 170916 225020
rect 171046 225040 171048 225049
rect 171100 225040 171102 225049
rect 171046 224975 171102 224984
rect 170956 224256 171008 224262
rect 170954 224224 170956 224233
rect 171094 224256 171146 224262
rect 171008 224224 171010 224233
rect 171428 224233 171456 229066
rect 172072 228682 172100 231676
rect 172426 228848 172482 228857
rect 172426 228783 172482 228792
rect 172242 228712 172298 228721
rect 172060 228676 172112 228682
rect 172242 228647 172244 228656
rect 172060 228618 172112 228624
rect 172296 228647 172298 228656
rect 172244 228618 172296 228624
rect 171094 224198 171146 224204
rect 171414 224224 171470 224233
rect 170954 224159 171010 224168
rect 171106 224074 171134 224198
rect 171414 224159 171470 224168
rect 170968 224046 171134 224074
rect 170968 223961 170996 224046
rect 170954 223952 171010 223961
rect 170954 223887 171010 223896
rect 170402 223272 170458 223281
rect 170402 223207 170458 223216
rect 171230 222320 171286 222329
rect 171230 222255 171286 222264
rect 171244 222170 171272 222255
rect 171060 222154 171272 222170
rect 171048 222148 171272 222154
rect 171100 222142 171272 222148
rect 171048 222090 171100 222096
rect 171046 221912 171102 221921
rect 171046 221847 171102 221856
rect 171506 221912 171562 221921
rect 171506 221847 171508 221856
rect 170772 220516 170824 220522
rect 170772 220458 170824 220464
rect 169944 218612 169996 218618
rect 169944 218554 169996 218560
rect 169576 218068 169628 218074
rect 169576 218010 169628 218016
rect 169300 217932 169352 217938
rect 169300 217874 169352 217880
rect 169956 217138 169984 218554
rect 170784 217274 170812 220458
rect 171060 218210 171088 221847
rect 171560 221847 171562 221856
rect 171508 221818 171560 221824
rect 172440 219434 172468 228783
rect 172716 220658 172744 231676
rect 172992 231662 173374 231690
rect 172992 222018 173020 231662
rect 174004 228818 174032 231676
rect 174174 228848 174230 228857
rect 173992 228812 174044 228818
rect 174174 228783 174176 228792
rect 173992 228754 174044 228760
rect 174228 228783 174230 228792
rect 174176 228754 174228 228760
rect 174648 227594 174676 231676
rect 174818 228848 174874 228857
rect 174818 228783 174874 228792
rect 174636 227588 174688 227594
rect 174636 227530 174688 227536
rect 174832 224210 174860 228783
rect 175292 228682 175320 231676
rect 175568 231662 175950 231690
rect 175280 228676 175332 228682
rect 175280 228618 175332 228624
rect 175188 227452 175240 227458
rect 175188 227394 175240 227400
rect 174556 224182 174860 224210
rect 172980 222012 173032 222018
rect 172980 221954 173032 221960
rect 172704 220652 172756 220658
rect 172704 220594 172756 220600
rect 172348 219406 172468 219434
rect 171048 218204 171100 218210
rect 171048 218146 171100 218152
rect 171600 218204 171652 218210
rect 171600 218146 171652 218152
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217246 170812 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217246
rect 171612 217138 171640 218146
rect 172348 217274 172376 219406
rect 174556 218482 174584 224182
rect 174912 222216 174964 222222
rect 174912 222158 174964 222164
rect 174544 218476 174596 218482
rect 174544 218418 174596 218424
rect 174728 218476 174780 218482
rect 174728 218418 174780 218424
rect 173256 218068 173308 218074
rect 173256 218010 173308 218016
rect 174084 218068 174136 218074
rect 174084 218010 174136 218016
rect 172348 217246 172422 217274
rect 171566 217110 171640 217138
rect 171566 216988 171594 217110
rect 172394 216988 172422 217246
rect 173268 217138 173296 218010
rect 174096 217138 174124 218010
rect 174740 217938 174768 218418
rect 174728 217932 174780 217938
rect 174728 217874 174780 217880
rect 174924 217274 174952 222158
rect 175200 218074 175228 227394
rect 175568 222630 175596 231662
rect 176580 229906 176608 231676
rect 176948 231662 177238 231690
rect 177408 231662 177882 231690
rect 178052 231662 178526 231690
rect 176568 229900 176620 229906
rect 176568 229842 176620 229848
rect 175738 228848 175794 228857
rect 175738 228783 175740 228792
rect 175792 228783 175794 228792
rect 175740 228754 175792 228760
rect 176658 226128 176714 226137
rect 176658 226063 176714 226072
rect 176672 225978 176700 226063
rect 176626 225950 176700 225978
rect 176626 225894 176654 225950
rect 176292 225888 176344 225894
rect 175936 225836 176292 225842
rect 175936 225830 176344 225836
rect 176614 225888 176666 225894
rect 176614 225830 176666 225836
rect 176752 225888 176804 225894
rect 176752 225830 176804 225836
rect 175936 225814 176332 225830
rect 175936 225758 175964 225814
rect 175924 225752 175976 225758
rect 175924 225694 175976 225700
rect 176764 225321 176792 225830
rect 176948 225729 176976 231662
rect 176934 225720 176990 225729
rect 176934 225655 176990 225664
rect 176474 225312 176530 225321
rect 176474 225247 176530 225256
rect 176750 225312 176806 225321
rect 176750 225247 176806 225256
rect 176108 223304 176160 223310
rect 176108 223246 176160 223252
rect 176292 223304 176344 223310
rect 176292 223246 176344 223252
rect 176120 222766 176148 223246
rect 176108 222760 176160 222766
rect 176108 222702 176160 222708
rect 175556 222624 175608 222630
rect 175556 222566 175608 222572
rect 176304 222222 176332 223246
rect 176292 222216 176344 222222
rect 176292 222158 176344 222164
rect 176108 222080 176160 222086
rect 176106 222048 176108 222057
rect 176160 222048 176162 222057
rect 176106 221983 176162 221992
rect 176292 222012 176344 222018
rect 176292 221954 176344 221960
rect 175740 218204 175792 218210
rect 175740 218146 175792 218152
rect 175188 218068 175240 218074
rect 175188 218010 175240 218016
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217246 174952 217274
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217246
rect 175752 217138 175780 218146
rect 176304 218074 176332 221954
rect 176488 218210 176516 225247
rect 177408 224954 177436 231662
rect 177580 229900 177632 229906
rect 177580 229842 177632 229848
rect 176856 224926 177436 224954
rect 176658 222320 176714 222329
rect 176658 222255 176714 222264
rect 176672 222154 176700 222255
rect 176660 222148 176712 222154
rect 176660 222090 176712 222096
rect 176856 222057 176884 224926
rect 177212 224800 177264 224806
rect 177212 224742 177264 224748
rect 177396 224800 177448 224806
rect 177396 224742 177448 224748
rect 177224 224534 177252 224742
rect 177028 224528 177080 224534
rect 177028 224470 177080 224476
rect 177212 224528 177264 224534
rect 177212 224470 177264 224476
rect 177040 224346 177068 224470
rect 177408 224346 177436 224742
rect 177040 224318 177436 224346
rect 176842 222048 176898 222057
rect 176842 221983 176898 221992
rect 177394 221776 177450 221785
rect 177394 221711 177450 221720
rect 177408 221338 177436 221711
rect 177396 221332 177448 221338
rect 177396 221274 177448 221280
rect 177212 220652 177264 220658
rect 177212 220594 177264 220600
rect 177224 219978 177252 220594
rect 177212 219972 177264 219978
rect 177212 219914 177264 219920
rect 177396 219972 177448 219978
rect 177396 219914 177448 219920
rect 176476 218204 176528 218210
rect 176476 218146 176528 218152
rect 176292 218068 176344 218074
rect 176292 218010 176344 218016
rect 176568 218068 176620 218074
rect 176568 218010 176620 218016
rect 176580 217138 176608 218010
rect 177408 217138 177436 219914
rect 177592 218074 177620 229842
rect 178052 221513 178080 231662
rect 179156 229226 179184 231676
rect 179144 229220 179196 229226
rect 179144 229162 179196 229168
rect 179800 229090 179828 231676
rect 179984 231662 180458 231690
rect 180812 231662 181102 231690
rect 179788 229084 179840 229090
rect 179788 229026 179840 229032
rect 179052 227588 179104 227594
rect 179052 227530 179104 227536
rect 178038 221504 178094 221513
rect 178038 221439 178094 221448
rect 178224 221332 178276 221338
rect 178224 221274 178276 221280
rect 177580 218068 177632 218074
rect 177580 218010 177632 218016
rect 178236 217138 178264 221274
rect 179064 217274 179092 227530
rect 179984 222154 180012 231662
rect 180616 229084 180668 229090
rect 180616 229026 180668 229032
rect 179972 222148 180024 222154
rect 179972 222090 180024 222096
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 175706 217110 175780 217138
rect 176534 217110 176608 217138
rect 177362 217110 177436 217138
rect 178190 217110 178264 217138
rect 179018 217246 179092 217274
rect 175706 216988 175734 217110
rect 176534 216988 176562 217110
rect 177362 216988 177390 217110
rect 178190 216988 178218 217110
rect 179018 216988 179046 217246
rect 179892 217138 179920 218146
rect 180628 217274 180656 229026
rect 180812 226137 180840 231662
rect 181732 230042 181760 231676
rect 181720 230036 181772 230042
rect 181720 229978 181772 229984
rect 181628 229220 181680 229226
rect 181628 229162 181680 229168
rect 180798 226128 180854 226137
rect 180798 226063 180854 226072
rect 181074 226128 181130 226137
rect 181074 226063 181130 226072
rect 181088 225894 181116 226063
rect 181076 225888 181128 225894
rect 181076 225830 181128 225836
rect 181444 225752 181496 225758
rect 181444 225694 181496 225700
rect 181456 225486 181484 225694
rect 181444 225480 181496 225486
rect 181444 225422 181496 225428
rect 181640 224954 181668 229162
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 181088 224926 181668 224954
rect 180892 223032 180944 223038
rect 180892 222974 180944 222980
rect 180904 222222 180932 222974
rect 180892 222216 180944 222222
rect 180892 222158 180944 222164
rect 181088 218618 181116 224926
rect 181260 224800 181312 224806
rect 181260 224742 181312 224748
rect 181272 224618 181300 224742
rect 181272 224590 181760 224618
rect 181732 224534 181760 224590
rect 181720 224528 181772 224534
rect 181720 224470 181772 224476
rect 181444 223304 181496 223310
rect 181444 223246 181496 223252
rect 181628 223304 181680 223310
rect 181628 223246 181680 223252
rect 181456 223038 181484 223246
rect 181444 223032 181496 223038
rect 181444 222974 181496 222980
rect 181640 222766 181668 223246
rect 181628 222760 181680 222766
rect 181628 222702 181680 222708
rect 181628 222080 181680 222086
rect 181628 222022 181680 222028
rect 181444 222012 181496 222018
rect 181444 221954 181496 221960
rect 181258 221504 181314 221513
rect 181258 221439 181314 221448
rect 181272 221338 181300 221439
rect 181456 221338 181484 221954
rect 181260 221332 181312 221338
rect 181260 221274 181312 221280
rect 181444 221332 181496 221338
rect 181444 221274 181496 221280
rect 181076 218612 181128 218618
rect 181076 218554 181128 218560
rect 181640 217274 181668 222022
rect 182652 220658 182680 231662
rect 183284 225480 183336 225486
rect 183284 225422 183336 225428
rect 182640 220652 182692 220658
rect 182640 220594 182692 220600
rect 183100 220652 183152 220658
rect 183100 220594 183152 220600
rect 182364 218612 182416 218618
rect 182364 218554 182416 218560
rect 180628 217246 180702 217274
rect 179846 217110 179920 217138
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181502 217246 181668 217274
rect 181502 216988 181530 217246
rect 182376 217138 182404 218554
rect 182330 217110 182404 217138
rect 183112 217138 183140 220594
rect 183296 218618 183324 225422
rect 183848 224534 183876 231662
rect 184308 230178 184336 231676
rect 184296 230172 184348 230178
rect 184296 230114 184348 230120
rect 184204 230036 184256 230042
rect 184204 229978 184256 229984
rect 183836 224528 183888 224534
rect 183836 224470 183888 224476
rect 184020 224528 184072 224534
rect 184020 224470 184072 224476
rect 183284 218612 183336 218618
rect 183284 218554 183336 218560
rect 184032 217138 184060 224470
rect 184216 220658 184244 229978
rect 184952 228954 184980 231676
rect 185136 231662 185610 231690
rect 185780 231662 186254 231690
rect 184940 228948 184992 228954
rect 184940 228890 184992 228896
rect 184846 225720 184902 225729
rect 184846 225655 184902 225664
rect 184204 220652 184256 220658
rect 184204 220594 184256 220600
rect 184388 220652 184440 220658
rect 184388 220594 184440 220600
rect 184400 219978 184428 220594
rect 184388 219972 184440 219978
rect 184388 219914 184440 219920
rect 184860 217274 184888 225655
rect 185136 224954 185164 231662
rect 185780 229242 185808 231662
rect 185044 224926 185164 224954
rect 185228 229214 185808 229242
rect 185044 221785 185072 224926
rect 185228 222222 185256 229214
rect 185676 229084 185728 229090
rect 185676 229026 185728 229032
rect 185688 225570 185716 229026
rect 186688 227724 186740 227730
rect 186688 227666 186740 227672
rect 186042 226128 186098 226137
rect 186042 226063 186098 226072
rect 186056 225978 186084 226063
rect 186272 226026 186328 226035
rect 186056 225950 186176 225978
rect 186272 225961 186328 225970
rect 186412 226024 186464 226030
rect 186412 225966 186464 225972
rect 186148 225894 186176 225950
rect 185952 225888 186004 225894
rect 185952 225830 186004 225836
rect 186136 225888 186188 225894
rect 186136 225830 186188 225836
rect 185964 225740 185992 225830
rect 185964 225712 186084 225740
rect 186424 225729 186452 225966
rect 186700 225758 186728 227666
rect 186688 225752 186740 225758
rect 185688 225542 185992 225570
rect 185676 225480 185728 225486
rect 185674 225448 185676 225457
rect 185728 225448 185730 225457
rect 185674 225383 185730 225392
rect 185964 224954 185992 225542
rect 186056 225434 186084 225712
rect 186410 225720 186466 225729
rect 186688 225694 186740 225700
rect 186872 225752 186924 225758
rect 186872 225694 186924 225700
rect 186410 225655 186466 225664
rect 186884 225570 186912 225694
rect 186608 225542 186912 225570
rect 186608 225457 186636 225542
rect 186594 225448 186650 225457
rect 186056 225406 186360 225434
rect 186332 225185 186360 225406
rect 186594 225383 186650 225392
rect 186870 225448 186926 225457
rect 186870 225383 186926 225392
rect 186884 225214 186912 225383
rect 186872 225208 186924 225214
rect 186318 225176 186374 225185
rect 186872 225150 186924 225156
rect 186318 225111 186374 225120
rect 187068 224954 187096 231798
rect 187252 231662 187542 231690
rect 187896 231662 188186 231690
rect 187252 227730 187280 231662
rect 187240 227724 187292 227730
rect 187240 227666 187292 227672
rect 187238 225992 187294 226001
rect 187238 225927 187294 225936
rect 187252 225214 187280 225927
rect 187240 225208 187292 225214
rect 187240 225150 187292 225156
rect 185688 224926 185992 224954
rect 186884 224926 187096 224954
rect 185216 222216 185268 222222
rect 185216 222158 185268 222164
rect 185030 221776 185086 221785
rect 185030 221711 185086 221720
rect 185688 217274 185716 224926
rect 186884 224262 186912 224926
rect 187056 224800 187108 224806
rect 187056 224742 187108 224748
rect 187332 224800 187384 224806
rect 187332 224742 187384 224748
rect 187068 224262 187096 224742
rect 186872 224256 186924 224262
rect 186872 224198 186924 224204
rect 187056 224256 187108 224262
rect 187056 224198 187108 224204
rect 185860 222012 185912 222018
rect 185860 221954 185912 221960
rect 185872 221513 185900 221954
rect 185858 221504 185914 221513
rect 185858 221439 185914 221448
rect 186504 218476 186556 218482
rect 186504 218418 186556 218424
rect 183112 217110 183186 217138
rect 182330 216988 182358 217110
rect 183158 216988 183186 217110
rect 183986 217110 184060 217138
rect 184814 217246 184888 217274
rect 185642 217246 185716 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185642 216988 185670 217246
rect 186516 217138 186544 218418
rect 187344 217274 187372 224742
rect 187896 221066 187924 231662
rect 188342 228848 188398 228857
rect 188342 228783 188344 228792
rect 188396 228783 188398 228792
rect 188344 228754 188396 228760
rect 188816 224262 188844 231676
rect 189460 230314 189488 231676
rect 189736 231662 190118 231690
rect 189448 230308 189500 230314
rect 189448 230250 189500 230256
rect 189736 226778 189764 231662
rect 190184 230036 190236 230042
rect 190184 229978 190236 229984
rect 189724 226772 189776 226778
rect 189724 226714 189776 226720
rect 188804 224256 188856 224262
rect 188804 224198 188856 224204
rect 188988 224256 189040 224262
rect 188988 224198 189040 224204
rect 187884 221060 187936 221066
rect 187884 221002 187936 221008
rect 188160 221060 188212 221066
rect 188160 221002 188212 221008
rect 188172 217274 188200 221002
rect 189000 217274 189028 224198
rect 190196 222194 190224 229978
rect 190368 229084 190420 229090
rect 190368 229026 190420 229032
rect 190380 228857 190408 229026
rect 190366 228848 190422 228857
rect 190366 228783 190422 228792
rect 190748 226914 190776 231676
rect 190920 230308 190972 230314
rect 190920 230250 190972 230256
rect 190932 229770 190960 230250
rect 190920 229764 190972 229770
rect 190920 229706 190972 229712
rect 190736 226908 190788 226914
rect 190736 226850 190788 226856
rect 190736 225480 190788 225486
rect 190736 225422 190788 225428
rect 190748 224806 190776 225422
rect 190736 224800 190788 224806
rect 190736 224742 190788 224748
rect 191392 224670 191420 231676
rect 191564 230172 191616 230178
rect 191564 230114 191616 230120
rect 191576 229906 191604 230114
rect 191564 229900 191616 229906
rect 191564 229842 191616 229848
rect 191564 227724 191616 227730
rect 191564 227666 191616 227672
rect 191380 224664 191432 224670
rect 191380 224606 191432 224612
rect 190196 222166 190316 222194
rect 190092 219156 190144 219162
rect 190092 219098 190144 219104
rect 189816 218068 189868 218074
rect 189816 218010 189868 218016
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 188126 217246 188200 217274
rect 188954 217246 189028 217274
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188126 216988 188154 217246
rect 188954 216988 188982 217246
rect 189828 217138 189856 218010
rect 190104 217938 190132 219098
rect 190288 218074 190316 222166
rect 190644 219972 190696 219978
rect 190644 219914 190696 219920
rect 190276 218068 190328 218074
rect 190276 218010 190328 218016
rect 190092 217932 190144 217938
rect 190092 217874 190144 217880
rect 190656 217274 190684 219914
rect 191576 219434 191604 227666
rect 192036 223310 192064 231676
rect 192680 228002 192708 231676
rect 193338 231662 193536 231690
rect 192668 227996 192720 228002
rect 192668 227938 192720 227944
rect 192760 224664 192812 224670
rect 192760 224606 192812 224612
rect 192772 224126 192800 224606
rect 192760 224120 192812 224126
rect 192760 224062 192812 224068
rect 192944 224120 192996 224126
rect 192944 224062 192996 224068
rect 192024 223304 192076 223310
rect 192024 223246 192076 223252
rect 192116 222760 192168 222766
rect 192116 222702 192168 222708
rect 191484 219406 191604 219434
rect 191484 217274 191512 219406
rect 192128 218074 192156 222702
rect 192956 218074 192984 224062
rect 193508 219842 193536 231662
rect 193968 224398 193996 231676
rect 194612 229090 194640 231676
rect 194888 231662 195270 231690
rect 195532 231662 195914 231690
rect 194600 229084 194652 229090
rect 194600 229026 194652 229032
rect 194888 225457 194916 231662
rect 194874 225448 194930 225457
rect 194874 225383 194930 225392
rect 195532 225185 195560 231662
rect 195704 229084 195756 229090
rect 195704 229026 195756 229032
rect 195518 225176 195574 225185
rect 195518 225111 195574 225120
rect 195716 224954 195744 229026
rect 195888 226772 195940 226778
rect 195888 226714 195940 226720
rect 195900 225214 195928 226714
rect 195888 225208 195940 225214
rect 195888 225150 195940 225156
rect 195716 224926 195928 224954
rect 194508 224800 194560 224806
rect 194508 224742 194560 224748
rect 194324 224664 194376 224670
rect 194324 224606 194376 224612
rect 193956 224392 194008 224398
rect 193956 224334 194008 224340
rect 194140 224392 194192 224398
rect 194140 224334 194192 224340
rect 194152 224126 194180 224334
rect 194336 224126 194364 224606
rect 194140 224120 194192 224126
rect 194140 224062 194192 224068
rect 194324 224120 194376 224126
rect 194324 224062 194376 224068
rect 193496 219836 193548 219842
rect 193496 219778 193548 219784
rect 193128 219292 193180 219298
rect 193128 219234 193180 219240
rect 192116 218068 192168 218074
rect 192116 218010 192168 218016
rect 192300 218068 192352 218074
rect 192300 218010 192352 218016
rect 192944 218068 192996 218074
rect 192944 218010 192996 218016
rect 189782 217110 189856 217138
rect 190610 217246 190684 217274
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217246
rect 191438 216988 191466 217246
rect 192312 217138 192340 218010
rect 193140 217138 193168 219234
rect 194520 218074 194548 224742
rect 195612 224664 195664 224670
rect 195612 224606 195664 224612
rect 195244 221332 195296 221338
rect 195244 221274 195296 221280
rect 195428 221332 195480 221338
rect 195428 221274 195480 221280
rect 195256 221066 195284 221274
rect 195060 221060 195112 221066
rect 195060 221002 195112 221008
rect 195244 221060 195296 221066
rect 195244 221002 195296 221008
rect 195072 220946 195100 221002
rect 195440 220946 195468 221274
rect 195072 220918 195468 220946
rect 195058 219328 195114 219337
rect 195058 219263 195114 219272
rect 195428 219292 195480 219298
rect 195072 219162 195100 219263
rect 195428 219234 195480 219240
rect 195060 219156 195112 219162
rect 195060 219098 195112 219104
rect 195244 219156 195296 219162
rect 195244 219098 195296 219104
rect 195256 218618 195284 219098
rect 195440 218618 195468 219234
rect 195244 218612 195296 218618
rect 195244 218554 195296 218560
rect 195428 218612 195480 218618
rect 195428 218554 195480 218560
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217274 195652 224606
rect 195900 218074 195928 224926
rect 196544 224126 196572 231676
rect 196992 230308 197044 230314
rect 196992 230250 197044 230256
rect 197004 229094 197032 230250
rect 197188 229498 197216 231676
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 198936 231662 199134 231690
rect 199304 231662 199778 231690
rect 197176 229492 197228 229498
rect 197176 229434 197228 229440
rect 197004 229066 197124 229094
rect 196532 224120 196584 224126
rect 196532 224062 196584 224068
rect 196070 219328 196126 219337
rect 196070 219263 196072 219272
rect 196124 219263 196126 219272
rect 196072 219234 196124 219240
rect 197096 218074 197124 229066
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197740 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 197740 220794 197768 229066
rect 197912 227996 197964 228002
rect 197912 227938 197964 227944
rect 197728 220788 197780 220794
rect 197728 220730 197780 220736
rect 197268 219836 197320 219842
rect 197268 219778 197320 219784
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196440 218068 196492 218074
rect 196440 218010 196492 218016
rect 197084 218068 197136 218074
rect 197084 218010 197136 218016
rect 192266 217110 192340 217138
rect 193094 217110 193168 217138
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217246 195652 217274
rect 192266 216988 192294 217110
rect 193094 216988 193122 217110
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217246
rect 196452 217138 196480 218010
rect 197280 217274 197308 219778
rect 197924 219434 197952 227938
rect 198936 220930 198964 231662
rect 199304 226778 199332 231662
rect 200408 227866 200436 231676
rect 201052 228138 201080 231676
rect 201040 228132 201092 228138
rect 201040 228074 201092 228080
rect 201408 228132 201460 228138
rect 201408 228074 201460 228080
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 226908 200080 226914
rect 200028 226850 200080 226856
rect 199292 226772 199344 226778
rect 199292 226714 199344 226720
rect 199384 225208 199436 225214
rect 199384 225150 199436 225156
rect 198924 220924 198976 220930
rect 198924 220866 198976 220872
rect 198096 220788 198148 220794
rect 198096 220730 198148 220736
rect 197912 219428 197964 219434
rect 197912 219370 197964 219376
rect 198108 217274 198136 220730
rect 199396 219298 199424 225150
rect 199752 219428 199804 219434
rect 199752 219370 199804 219376
rect 199384 219292 199436 219298
rect 199384 219234 199436 219240
rect 198924 218068 198976 218074
rect 198924 218010 198976 218016
rect 196406 217110 196480 217138
rect 197234 217246 197308 217274
rect 198062 217246 198136 217274
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198062 216988 198090 217246
rect 198936 217138 198964 218010
rect 199764 217138 199792 219370
rect 200040 218074 200068 226850
rect 201224 224120 201276 224126
rect 201224 224062 201276 224068
rect 201236 219434 201264 224062
rect 201236 219406 201356 219434
rect 200580 219020 200632 219026
rect 200580 218962 200632 218968
rect 200028 218068 200080 218074
rect 200028 218010 200080 218016
rect 200592 217138 200620 218962
rect 201328 217274 201356 219406
rect 201420 219042 201448 228074
rect 201696 223718 201724 231676
rect 202340 230178 202368 231676
rect 202998 231662 203196 231690
rect 202328 230172 202380 230178
rect 202328 230114 202380 230120
rect 203168 225350 203196 231662
rect 203260 231662 203642 231690
rect 203260 229094 203288 231662
rect 203892 229492 203944 229498
rect 203892 229434 203944 229440
rect 203904 229094 203932 229434
rect 203260 229066 203472 229094
rect 203156 225344 203208 225350
rect 203156 225286 203208 225292
rect 202694 225176 202750 225185
rect 202694 225111 202750 225120
rect 201684 223712 201736 223718
rect 201684 223654 201736 223660
rect 201420 219026 201540 219042
rect 201420 219020 201552 219026
rect 201420 219014 201500 219020
rect 201500 218962 201552 218968
rect 202708 218074 202736 225111
rect 203248 221196 203300 221202
rect 203248 221138 203300 221144
rect 203260 220930 203288 221138
rect 203248 220924 203300 220930
rect 203248 220866 203300 220872
rect 203444 219570 203472 229066
rect 203720 229066 203932 229094
rect 203432 219564 203484 219570
rect 203432 219506 203484 219512
rect 203720 218074 203748 229066
rect 203892 225616 203944 225622
rect 203892 225558 203944 225564
rect 203904 225350 203932 225558
rect 203892 225344 203944 225350
rect 203892 225286 203944 225292
rect 204272 223854 204300 231676
rect 204916 229094 204944 231676
rect 204548 229066 204944 229094
rect 205192 231662 205574 231690
rect 205836 231662 206218 231690
rect 206480 231662 206862 231690
rect 205192 229094 205220 231662
rect 205364 230308 205416 230314
rect 205364 230250 205416 230256
rect 205376 229498 205404 230250
rect 205364 229492 205416 229498
rect 205364 229434 205416 229440
rect 205192 229066 205312 229094
rect 204548 228002 204576 229066
rect 204720 228812 204772 228818
rect 204720 228754 204772 228760
rect 204904 228812 204956 228818
rect 204904 228754 204956 228760
rect 204732 228426 204760 228754
rect 204916 228546 204944 228754
rect 204904 228540 204956 228546
rect 204904 228482 204956 228488
rect 205088 228540 205140 228546
rect 205088 228482 205140 228488
rect 205100 228426 205128 228482
rect 204732 228398 205128 228426
rect 204536 227996 204588 228002
rect 204536 227938 204588 227944
rect 205284 226506 205312 229066
rect 205456 227996 205508 228002
rect 205456 227938 205508 227944
rect 205272 226500 205324 226506
rect 205272 226442 205324 226448
rect 204904 225616 204956 225622
rect 204904 225558 204956 225564
rect 204916 225214 204944 225558
rect 204904 225208 204956 225214
rect 205088 225208 205140 225214
rect 204904 225150 204956 225156
rect 205086 225176 205088 225185
rect 205140 225176 205142 225185
rect 205086 225111 205142 225120
rect 204732 224454 205128 224482
rect 204732 224126 204760 224454
rect 205100 224398 205128 224454
rect 204904 224392 204956 224398
rect 204904 224334 204956 224340
rect 205088 224392 205140 224398
rect 205088 224334 205140 224340
rect 204916 224126 204944 224334
rect 204720 224120 204772 224126
rect 204720 224062 204772 224068
rect 204904 224120 204956 224126
rect 204904 224062 204956 224068
rect 204260 223848 204312 223854
rect 204260 223790 204312 223796
rect 205272 223848 205324 223854
rect 205272 223790 205324 223796
rect 203892 223304 203944 223310
rect 203892 223246 203944 223252
rect 202236 218068 202288 218074
rect 202236 218010 202288 218016
rect 202696 218068 202748 218074
rect 202696 218010 202748 218016
rect 203064 218068 203116 218074
rect 203064 218010 203116 218016
rect 203708 218068 203760 218074
rect 203708 218010 203760 218016
rect 201328 217246 201402 217274
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217110 200620 217138
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202248 217138 202276 218010
rect 203076 217138 203104 218010
rect 203904 217274 203932 223246
rect 204904 221604 204956 221610
rect 204904 221546 204956 221552
rect 205088 221604 205140 221610
rect 205088 221546 205140 221552
rect 204916 221066 204944 221546
rect 205100 221202 205128 221546
rect 205088 221196 205140 221202
rect 205088 221138 205140 221144
rect 204904 221060 204956 221066
rect 204904 221002 204956 221008
rect 205284 219434 205312 223790
rect 204720 219428 204772 219434
rect 204720 219370 204772 219376
rect 204916 219406 205312 219434
rect 204732 219162 204760 219370
rect 204720 219156 204772 219162
rect 204720 219098 204772 219104
rect 204916 219026 204944 219406
rect 204904 219020 204956 219026
rect 204904 218962 204956 218968
rect 204720 218068 204772 218074
rect 204720 218010 204772 218016
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218010
rect 205468 217274 205496 227938
rect 205836 219706 205864 231662
rect 206008 221196 206060 221202
rect 206008 221138 206060 221144
rect 205824 219700 205876 219706
rect 205824 219642 205876 219648
rect 206020 218074 206048 221138
rect 206480 220930 206508 231662
rect 207492 222766 207520 231676
rect 207768 231662 208150 231690
rect 207768 225350 207796 231662
rect 207756 225344 207808 225350
rect 207756 225286 207808 225292
rect 208032 225344 208084 225350
rect 208032 225286 208084 225292
rect 207480 222760 207532 222766
rect 207480 222702 207532 222708
rect 206468 220924 206520 220930
rect 206468 220866 206520 220872
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206376 219020 206428 219026
rect 206376 218962 206428 218968
rect 206008 218068 206060 218074
rect 206008 218010 206060 218016
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218962
rect 207216 217274 207244 219642
rect 208044 217274 208072 225286
rect 208780 222358 208808 231676
rect 209424 224942 209452 231676
rect 210068 229634 210096 231676
rect 210056 229628 210108 229634
rect 210056 229570 210108 229576
rect 210240 229628 210292 229634
rect 210240 229570 210292 229576
rect 209412 224936 209464 224942
rect 209412 224878 209464 224884
rect 209688 224936 209740 224942
rect 209688 224878 209740 224884
rect 209504 222760 209556 222766
rect 209504 222702 209556 222708
rect 208768 222352 208820 222358
rect 208768 222294 208820 222300
rect 209516 219434 209544 222702
rect 209700 219450 209728 224878
rect 210252 222766 210280 229570
rect 210712 228818 210740 231676
rect 210700 228812 210752 228818
rect 210700 228754 210752 228760
rect 210240 222760 210292 222766
rect 210240 222702 210292 222708
rect 210976 222352 211028 222358
rect 210976 222294 211028 222300
rect 210240 220380 210292 220386
rect 210240 220322 210292 220328
rect 210252 219570 210280 220322
rect 210240 219564 210292 219570
rect 210240 219506 210292 219512
rect 209700 219434 209820 219450
rect 208860 219428 208912 219434
rect 209516 219406 209636 219434
rect 209700 219428 209832 219434
rect 209700 219422 209780 219428
rect 208860 219370 208912 219376
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 207998 217246 208072 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 207998 216988 208026 217246
rect 208872 217138 208900 219370
rect 209608 217274 209636 219406
rect 209780 219370 209832 219376
rect 209792 219339 209820 219370
rect 210988 218074 211016 222294
rect 211356 220250 211384 231676
rect 211632 231662 212014 231690
rect 211632 221066 211660 231662
rect 212172 226772 212224 226778
rect 212172 226714 212224 226720
rect 211988 221468 212040 221474
rect 211988 221410 212040 221416
rect 212000 221066 212028 221410
rect 211620 221060 211672 221066
rect 211620 221002 211672 221008
rect 211988 221060 212040 221066
rect 211988 221002 212040 221008
rect 211344 220244 211396 220250
rect 211344 220186 211396 220192
rect 211344 220108 211396 220114
rect 211344 220050 211396 220056
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 209608 217246 209682 217274
rect 208826 217110 208900 217138
rect 208826 216988 208854 217110
rect 209654 216988 209682 217246
rect 210528 217138 210556 218010
rect 211356 217274 211384 220050
rect 212184 217274 212212 226714
rect 212644 223854 212672 231676
rect 213288 227050 213316 231676
rect 213946 231662 214144 231690
rect 214116 229094 214144 231662
rect 213932 229066 214144 229094
rect 214300 231662 214590 231690
rect 213276 227044 213328 227050
rect 213276 226986 213328 226992
rect 213184 226500 213236 226506
rect 213184 226442 213236 226448
rect 212632 223848 212684 223854
rect 212632 223790 212684 223796
rect 213196 218754 213224 226442
rect 213932 222850 213960 229066
rect 214104 228812 214156 228818
rect 214104 228754 214156 228760
rect 214116 228410 214144 228754
rect 214104 228404 214156 228410
rect 214104 228346 214156 228352
rect 213932 222822 214052 222850
rect 213828 222760 213880 222766
rect 213828 222702 213880 222708
rect 213184 218748 213236 218754
rect 213184 218690 213236 218696
rect 213552 218748 213604 218754
rect 213552 218690 213604 218696
rect 213564 218346 213592 218690
rect 213552 218340 213604 218346
rect 213552 218282 213604 218288
rect 213000 218068 213052 218074
rect 213000 218010 213052 218016
rect 210482 217110 210556 217138
rect 211310 217246 211384 217274
rect 212138 217246 212212 217274
rect 210482 216988 210510 217110
rect 211310 216988 211338 217246
rect 212138 216988 212166 217246
rect 213012 217138 213040 218010
rect 213840 217274 213868 222702
rect 214024 220386 214052 222822
rect 214300 222748 214328 231662
rect 215220 230450 215248 231676
rect 215208 230444 215260 230450
rect 215208 230386 215260 230392
rect 214748 228268 214800 228274
rect 214748 228210 214800 228216
rect 214760 228002 214788 228210
rect 214748 227996 214800 228002
rect 214748 227938 214800 227944
rect 215864 226166 215892 231676
rect 216232 231662 216522 231690
rect 215852 226160 215904 226166
rect 215852 226102 215904 226108
rect 215944 223848 215996 223854
rect 215944 223790 215996 223796
rect 214208 222720 214328 222748
rect 214208 221066 214236 222720
rect 214748 222624 214800 222630
rect 214748 222566 214800 222572
rect 214380 222488 214432 222494
rect 214380 222430 214432 222436
rect 214392 222170 214420 222430
rect 214760 222358 214788 222566
rect 214748 222352 214800 222358
rect 214748 222294 214800 222300
rect 214932 222284 214984 222290
rect 214932 222226 214984 222232
rect 214944 222170 214972 222226
rect 214392 222142 214972 222170
rect 214656 221604 214708 221610
rect 214656 221546 214708 221552
rect 214196 221060 214248 221066
rect 214196 221002 214248 221008
rect 214012 220380 214064 220386
rect 214012 220322 214064 220328
rect 214668 217274 214696 221546
rect 215956 218890 215984 223790
rect 216232 222290 216260 231662
rect 216496 226160 216548 226166
rect 216496 226102 216548 226108
rect 216220 222284 216272 222290
rect 216220 222226 216272 222232
rect 215944 218884 215996 218890
rect 215944 218826 215996 218832
rect 216312 218340 216364 218346
rect 216312 218282 216364 218288
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 214622 217246 214696 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214622 216988 214650 217246
rect 215496 217138 215524 218010
rect 216324 217138 216352 218282
rect 216508 218074 216536 226102
rect 217152 223990 217180 231676
rect 217796 226506 217824 231676
rect 218440 228818 218468 231676
rect 218624 231662 219098 231690
rect 218428 228812 218480 228818
rect 218428 228754 218480 228760
rect 217784 226500 217836 226506
rect 217784 226442 217836 226448
rect 217140 223984 217192 223990
rect 217140 223926 217192 223932
rect 217324 223984 217376 223990
rect 217324 223926 217376 223932
rect 217140 220244 217192 220250
rect 217140 220186 217192 220192
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 217152 217274 217180 220186
rect 217336 218754 217364 223926
rect 218624 219570 218652 231662
rect 219348 228812 219400 228818
rect 219348 228754 219400 228760
rect 218612 219564 218664 219570
rect 218612 219506 218664 219512
rect 217968 218884 218020 218890
rect 217968 218826 218020 218832
rect 217324 218748 217376 218754
rect 217324 218690 217376 218696
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218826
rect 219360 218754 219388 228754
rect 219728 222494 219756 231676
rect 220372 229362 220400 231676
rect 220360 229356 220412 229362
rect 220360 229298 220412 229304
rect 221016 226370 221044 231676
rect 221004 226364 221056 226370
rect 221004 226306 221056 226312
rect 221660 222902 221688 231676
rect 222016 226636 222068 226642
rect 222016 226578 222068 226584
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221648 222896 221700 222902
rect 221648 222838 221700 222844
rect 219716 222488 219768 222494
rect 219716 222430 219768 222436
rect 220084 222488 220136 222494
rect 220084 222430 220136 222436
rect 220096 218890 220124 222430
rect 220452 222352 220504 222358
rect 220452 222294 220504 222300
rect 220084 218884 220136 218890
rect 220084 218826 220136 218832
rect 218796 218748 218848 218754
rect 218796 218690 218848 218696
rect 219348 218748 219400 218754
rect 219348 218690 219400 218696
rect 219624 218748 219676 218754
rect 219624 218690 219676 218696
rect 218808 217138 218836 218690
rect 219636 217138 219664 218690
rect 220464 217274 220492 222294
rect 221648 219496 221700 219502
rect 221648 219438 221700 219444
rect 221096 218748 221148 218754
rect 221096 218690 221148 218696
rect 221108 218210 221136 218690
rect 221660 218346 221688 219438
rect 221648 218340 221700 218346
rect 221648 218282 221700 218288
rect 221844 218210 221872 226442
rect 221096 218204 221148 218210
rect 221096 218146 221148 218152
rect 221280 218204 221332 218210
rect 221280 218146 221332 218152
rect 221832 218204 221884 218210
rect 221832 218146 221884 218152
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218146
rect 222028 217274 222056 226578
rect 222304 223174 222332 231676
rect 222752 228404 222804 228410
rect 222752 228346 222804 228352
rect 222764 228002 222792 228346
rect 222752 227996 222804 228002
rect 222752 227938 222804 227944
rect 222476 226296 222528 226302
rect 222476 226238 222528 226244
rect 222488 225622 222516 226238
rect 222476 225616 222528 225622
rect 222476 225558 222528 225564
rect 222948 223854 222976 231676
rect 223396 230444 223448 230450
rect 223396 230386 223448 230392
rect 222936 223848 222988 223854
rect 222936 223790 222988 223796
rect 222292 223168 222344 223174
rect 222292 223110 222344 223116
rect 223408 218210 223436 230386
rect 223592 225078 223620 231676
rect 224040 228812 224092 228818
rect 224040 228754 224092 228760
rect 224052 228410 224080 228754
rect 224040 228404 224092 228410
rect 224040 228346 224092 228352
rect 224236 226114 224264 231676
rect 224052 226086 224264 226114
rect 224420 231662 224894 231690
rect 223580 225072 223632 225078
rect 223580 225014 223632 225020
rect 224052 223446 224080 226086
rect 224224 226024 224276 226030
rect 224224 225966 224276 225972
rect 224236 225622 224264 225966
rect 224224 225616 224276 225622
rect 224224 225558 224276 225564
rect 224040 223440 224092 223446
rect 224040 223382 224092 223388
rect 224224 223168 224276 223174
rect 224224 223110 224276 223116
rect 224236 218754 224264 223110
rect 224420 221746 224448 231662
rect 225524 226302 225552 231676
rect 225696 228404 225748 228410
rect 225696 228346 225748 228352
rect 225512 226296 225564 226302
rect 225512 226238 225564 226244
rect 224868 225072 224920 225078
rect 224868 225014 224920 225020
rect 224408 221740 224460 221746
rect 224408 221682 224460 221688
rect 224224 218748 224276 218754
rect 224224 218690 224276 218696
rect 224592 218340 224644 218346
rect 224592 218282 224644 218288
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 223396 218204 223448 218210
rect 223396 218146 223448 218152
rect 223764 218204 223816 218210
rect 223764 218146 223816 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 223776 217138 223804 218146
rect 224604 217138 224632 218282
rect 224880 218210 224908 225014
rect 225708 219434 225736 228346
rect 226168 228002 226196 231676
rect 226812 229094 226840 231676
rect 226720 229066 226840 229094
rect 226156 227996 226208 228002
rect 226156 227938 226208 227944
rect 226156 227860 226208 227866
rect 226156 227802 226208 227808
rect 225616 219406 225736 219434
rect 225616 218346 225644 219406
rect 225972 218884 226024 218890
rect 225972 218826 226024 218832
rect 225604 218340 225656 218346
rect 225604 218282 225656 218288
rect 224868 218204 224920 218210
rect 224868 218146 224920 218152
rect 225420 218204 225472 218210
rect 225420 218146 225472 218152
rect 225432 217138 225460 218146
rect 225984 217274 226012 218826
rect 226168 218210 226196 227802
rect 226720 223582 226748 229066
rect 227456 227322 227484 231676
rect 227444 227316 227496 227322
rect 227444 227258 227496 227264
rect 226892 227044 226944 227050
rect 226892 226986 226944 226992
rect 226708 223576 226760 223582
rect 226708 223518 226760 223524
rect 226904 219298 226932 226986
rect 228100 223990 228128 231676
rect 228744 227186 228772 231676
rect 229296 231662 229402 231690
rect 229664 231662 230046 231690
rect 228732 227180 228784 227186
rect 228732 227122 228784 227128
rect 229054 227044 229106 227050
rect 229054 226986 229106 226992
rect 229066 226930 229094 226986
rect 229020 226902 229094 226930
rect 229020 226506 229048 226902
rect 229008 226500 229060 226506
rect 229008 226442 229060 226448
rect 228732 226296 228784 226302
rect 228732 226238 228784 226244
rect 228088 223984 228140 223990
rect 228088 223926 228140 223932
rect 227076 221740 227128 221746
rect 227076 221682 227128 221688
rect 226892 219292 226944 219298
rect 226892 219234 226944 219240
rect 226156 218204 226208 218210
rect 226156 218146 226208 218152
rect 227088 217274 227116 221682
rect 227904 218340 227956 218346
rect 227904 218282 227956 218288
rect 225984 217246 226242 217274
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217110 224632 217138
rect 225386 217110 225460 217138
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217110
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 217246 227116 217274
rect 227042 216988 227070 217246
rect 227916 217138 227944 218282
rect 228744 217274 228772 226238
rect 229296 220522 229324 231662
rect 229664 221882 229692 231662
rect 230676 229226 230704 231676
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230664 229220 230716 229226
rect 230664 229162 230716 229168
rect 229652 221876 229704 221882
rect 229652 221818 229704 221824
rect 230388 221876 230440 221882
rect 230388 221818 230440 221824
rect 229284 220516 229336 220522
rect 229284 220458 229336 220464
rect 229192 220380 229244 220386
rect 229192 220322 229244 220328
rect 229204 218346 229232 220322
rect 229192 218340 229244 218346
rect 229192 218282 229244 218288
rect 229560 218204 229612 218210
rect 229560 218146 229612 218152
rect 227870 217110 227944 217138
rect 228698 217246 228772 217274
rect 227870 216988 227898 217110
rect 228698 216988 228726 217246
rect 229572 217138 229600 218146
rect 230400 217274 230428 221818
rect 231136 219434 231164 229434
rect 231320 228818 231348 231676
rect 231308 228812 231360 228818
rect 231308 228754 231360 228760
rect 231964 227458 231992 231676
rect 232148 231662 232622 231690
rect 231952 227452 232004 227458
rect 231952 227394 232004 227400
rect 231676 223984 231728 223990
rect 231676 223926 231728 223932
rect 231044 219406 231164 219434
rect 231044 218210 231072 219406
rect 231688 218210 231716 223926
rect 232148 221474 232176 231662
rect 233252 227322 233280 231676
rect 233240 227316 233292 227322
rect 233240 227258 233292 227264
rect 232504 226500 232556 226506
rect 232504 226442 232556 226448
rect 232136 221468 232188 221474
rect 232136 221410 232188 221416
rect 232516 219434 232544 226442
rect 233896 226030 233924 231676
rect 234080 231662 234554 231690
rect 234816 231662 235198 231690
rect 233884 226024 233936 226030
rect 233884 225966 233936 225972
rect 233700 224528 233752 224534
rect 233700 224470 233752 224476
rect 233884 224528 233936 224534
rect 233884 224470 233936 224476
rect 233712 223854 233740 224470
rect 233896 224126 233924 224470
rect 233884 224120 233936 224126
rect 233884 224062 233936 224068
rect 233700 223848 233752 223854
rect 233700 223790 233752 223796
rect 233148 222896 233200 222902
rect 233148 222838 233200 222844
rect 232504 219428 232556 219434
rect 232504 219370 232556 219376
rect 232872 219292 232924 219298
rect 232872 219234 232924 219240
rect 231032 218204 231084 218210
rect 231032 218146 231084 218152
rect 231216 218204 231268 218210
rect 231216 218146 231268 218152
rect 231676 218204 231728 218210
rect 231676 218146 231728 218152
rect 232044 218204 232096 218210
rect 232044 218146 232096 218152
rect 229526 217110 229600 217138
rect 230354 217246 230428 217274
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218146
rect 232056 217138 232084 218146
rect 232884 217138 232912 219234
rect 233160 218210 233188 222838
rect 234080 220658 234108 231662
rect 234528 227316 234580 227322
rect 234528 227258 234580 227264
rect 234344 225616 234396 225622
rect 234344 225558 234396 225564
rect 234068 220652 234120 220658
rect 234068 220594 234120 220600
rect 234356 219434 234384 225558
rect 234540 219434 234568 227258
rect 234816 223038 234844 231662
rect 235828 229770 235856 231676
rect 235816 229764 235868 229770
rect 235816 229706 235868 229712
rect 236472 227594 236500 231676
rect 236920 229764 236972 229770
rect 236920 229706 236972 229712
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 235908 227180 235960 227186
rect 235908 227122 235960 227128
rect 234804 223032 234856 223038
rect 234804 222974 234856 222980
rect 235172 223032 235224 223038
rect 235172 222974 235224 222980
rect 233700 219428 233752 219434
rect 234356 219406 234476 219434
rect 234540 219428 234672 219434
rect 234540 219406 234620 219428
rect 233700 219370 233752 219376
rect 233148 218204 233200 218210
rect 233148 218146 233200 218152
rect 233712 217138 233740 219370
rect 234448 217274 234476 219406
rect 234620 219370 234672 219376
rect 235184 218482 235212 222974
rect 235172 218476 235224 218482
rect 235172 218418 235224 218424
rect 235920 218210 235948 227122
rect 236932 218210 236960 229706
rect 237116 228682 237144 231676
rect 237576 231662 237774 231690
rect 237104 228676 237156 228682
rect 237104 228618 237156 228624
rect 237576 222018 237604 231662
rect 238404 223174 238432 231676
rect 239048 225894 239076 231676
rect 239404 228676 239456 228682
rect 239404 228618 239456 228624
rect 239036 225888 239088 225894
rect 239036 225830 239088 225836
rect 238668 223984 238720 223990
rect 238668 223926 238720 223932
rect 238392 223168 238444 223174
rect 238392 223110 238444 223116
rect 237564 222012 237616 222018
rect 237564 221954 237616 221960
rect 237104 221060 237156 221066
rect 237104 221002 237156 221008
rect 235356 218204 235408 218210
rect 235356 218146 235408 218152
rect 235908 218204 235960 218210
rect 235908 218146 235960 218152
rect 236184 218204 236236 218210
rect 236184 218146 236236 218152
rect 236920 218204 236972 218210
rect 236920 218146 236972 218152
rect 234448 217246 234522 217274
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217110 233740 217138
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217110
rect 234494 216988 234522 217246
rect 235368 217138 235396 218146
rect 236196 217138 236224 218146
rect 237116 217274 237144 221002
rect 237840 219292 237892 219298
rect 237840 219234 237892 219240
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237144 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219234
rect 238680 217274 238708 223926
rect 239416 219298 239444 228618
rect 239692 223854 239720 231676
rect 240152 231662 240350 231690
rect 239680 223848 239732 223854
rect 239680 223790 239732 223796
rect 240152 222154 240180 231662
rect 240980 229906 241008 231676
rect 240968 229900 241020 229906
rect 240968 229842 241020 229848
rect 241624 228954 241652 231676
rect 241612 228948 241664 228954
rect 241612 228890 241664 228896
rect 242268 225486 242296 231676
rect 242716 227792 242768 227798
rect 242716 227734 242768 227740
rect 242256 225480 242308 225486
rect 242256 225422 242308 225428
rect 241980 223848 242032 223854
rect 241980 223790 242032 223796
rect 240140 222148 240192 222154
rect 240140 222090 240192 222096
rect 241152 221468 241204 221474
rect 241152 221410 241204 221416
rect 240324 220652 240376 220658
rect 240324 220594 240376 220600
rect 239404 219292 239456 219298
rect 239404 219234 239456 219240
rect 239496 218476 239548 218482
rect 239496 218418 239548 218424
rect 237806 217110 237880 217138
rect 238634 217246 238708 217274
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 218418
rect 240336 217274 240364 220594
rect 241164 217274 241192 221410
rect 241992 217274 242020 223790
rect 239462 217110 239536 217138
rect 240290 217246 240364 217274
rect 241118 217246 241192 217274
rect 241946 217246 242020 217274
rect 242728 217274 242756 227734
rect 242912 225758 242940 231676
rect 243280 231662 243570 231690
rect 243832 231662 244214 231690
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 242900 225752 242952 225758
rect 242900 225694 242952 225700
rect 243280 223038 243308 231662
rect 243452 226024 243504 226030
rect 243452 225966 243504 225972
rect 243268 223032 243320 223038
rect 243268 222974 243320 222980
rect 243464 218618 243492 225966
rect 243832 224262 243860 231662
rect 243820 224256 243872 224262
rect 243820 224198 243872 224204
rect 243636 222012 243688 222018
rect 243636 221954 243688 221960
rect 243452 218612 243504 218618
rect 243452 218554 243504 218560
rect 243648 217274 243676 221954
rect 244476 219978 244504 231662
rect 245120 221338 245148 231662
rect 246132 230042 246160 231676
rect 246120 230036 246172 230042
rect 246120 229978 246172 229984
rect 245660 229900 245712 229906
rect 245660 229842 245712 229848
rect 245672 227798 245700 229842
rect 246304 228812 246356 228818
rect 246304 228754 246356 228760
rect 245660 227792 245712 227798
rect 245660 227734 245712 227740
rect 245292 223168 245344 223174
rect 245292 223110 245344 223116
rect 245108 221332 245160 221338
rect 245108 221274 245160 221280
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 244464 218340 244516 218346
rect 244464 218282 244516 218288
rect 242728 217246 242802 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217246
rect 241118 216988 241146 217246
rect 241946 216988 241974 217246
rect 242774 216988 242802 217246
rect 243602 217246 243676 217274
rect 243602 216988 243630 217246
rect 244476 217138 244504 218282
rect 245304 217274 245332 223110
rect 246120 219428 246172 219434
rect 246120 219370 246172 219376
rect 244430 217110 244504 217138
rect 245258 217246 245332 217274
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 219370
rect 246316 219162 246344 228754
rect 246776 224534 246804 231676
rect 247420 224806 247448 231676
rect 248064 227662 248092 231676
rect 248052 227656 248104 227662
rect 248052 227598 248104 227604
rect 248236 227452 248288 227458
rect 248236 227394 248288 227400
rect 247408 224800 247460 224806
rect 247408 224742 247460 224748
rect 246764 224528 246816 224534
rect 246764 224470 246816 224476
rect 247684 224528 247736 224534
rect 247684 224470 247736 224476
rect 246948 224256 247000 224262
rect 246948 224198 247000 224204
rect 246304 219156 246356 219162
rect 246304 219098 246356 219104
rect 246960 217274 246988 224198
rect 247696 218346 247724 224470
rect 247684 218340 247736 218346
rect 247684 218282 247736 218288
rect 248248 218074 248276 227394
rect 248708 226030 248736 231676
rect 248892 231662 249366 231690
rect 249904 231662 250010 231690
rect 248696 226024 248748 226030
rect 248696 225966 248748 225972
rect 248892 224670 248920 231662
rect 249708 225888 249760 225894
rect 249708 225830 249760 225836
rect 248880 224664 248932 224670
rect 248880 224606 248932 224612
rect 249064 224664 249116 224670
rect 249064 224606 249116 224612
rect 249076 218210 249104 224606
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218146
rect 249720 218074 249748 225830
rect 249904 219842 249932 231662
rect 250640 229090 250668 231676
rect 251284 230178 251312 231676
rect 251272 230172 251324 230178
rect 251272 230114 251324 230120
rect 251732 230036 251784 230042
rect 251732 229978 251784 229984
rect 250628 229084 250680 229090
rect 250628 229026 250680 229032
rect 251088 228948 251140 228954
rect 251088 228890 251140 228896
rect 250904 223032 250956 223038
rect 250904 222974 250956 222980
rect 249892 219836 249944 219842
rect 249892 219778 249944 219784
rect 250916 219434 250944 222974
rect 250916 219406 251036 219434
rect 249708 218068 249760 218074
rect 249708 218010 249760 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250272 217138 250300 218010
rect 251008 217274 251036 219406
rect 251100 218090 251128 228890
rect 251744 218210 251772 229978
rect 251928 226914 251956 231676
rect 252572 228138 252600 231676
rect 252756 231662 253230 231690
rect 252560 228132 252612 228138
rect 252560 228074 252612 228080
rect 252468 227588 252520 227594
rect 252468 227530 252520 227536
rect 251916 226908 251968 226914
rect 251916 226850 251968 226856
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 251100 218074 251220 218090
rect 252480 218074 252508 227530
rect 252756 220794 252784 231662
rect 253860 228818 253888 231676
rect 253848 228812 253900 228818
rect 253848 228754 253900 228760
rect 254504 225214 254532 231676
rect 254872 231662 255162 231690
rect 254492 225208 254544 225214
rect 254492 225150 254544 225156
rect 254872 223310 254900 231662
rect 255136 228812 255188 228818
rect 255136 228754 255188 228760
rect 254860 223304 254912 223310
rect 254860 223246 254912 223252
rect 252744 220788 252796 220794
rect 252744 220730 252796 220736
rect 253572 220788 253624 220794
rect 253572 220730 253624 220736
rect 252744 218612 252796 218618
rect 252744 218554 252796 218560
rect 251100 218068 251232 218074
rect 251100 218062 251180 218068
rect 251180 218010 251232 218016
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 251008 217246 251082 217274
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218554
rect 253584 217274 253612 220730
rect 254400 220516 254452 220522
rect 254400 220458 254452 220464
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 220458
rect 255148 217274 255176 228754
rect 255792 224398 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 257080 228274 257108 231676
rect 257264 231662 257738 231690
rect 258184 231662 258382 231690
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 255964 227792 256016 227798
rect 255964 227734 256016 227740
rect 255780 224392 255832 224398
rect 255780 224334 255832 224340
rect 255976 221082 256004 227734
rect 255884 221054 256004 221082
rect 255884 219026 255912 221054
rect 256056 220924 256108 220930
rect 256056 220866 256108 220872
rect 255872 219020 255924 219026
rect 255872 218962 255924 218968
rect 255148 217246 255222 217274
rect 254366 217110 254440 217138
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 220866
rect 256884 219972 256936 219978
rect 256884 219914 256936 219920
rect 256896 217274 256924 219914
rect 257264 219706 257292 231662
rect 258184 229094 258212 231662
rect 258184 229066 258396 229094
rect 257712 225752 257764 225758
rect 257712 225694 257764 225700
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 257724 217274 257752 225694
rect 258368 221202 258396 229066
rect 259012 227798 259040 231676
rect 259276 229084 259328 229090
rect 259276 229026 259328 229032
rect 259000 227792 259052 227798
rect 259000 227734 259052 227740
rect 258724 221876 258776 221882
rect 258724 221818 258776 221824
rect 258736 221610 258764 221818
rect 258540 221604 258592 221610
rect 258540 221546 258592 221552
rect 258724 221604 258776 221610
rect 258724 221546 258776 221552
rect 258552 221338 258580 221546
rect 258540 221332 258592 221338
rect 258540 221274 258592 221280
rect 258356 221196 258408 221202
rect 258356 221138 258408 221144
rect 259288 219162 259316 229026
rect 259656 224942 259684 231676
rect 259644 224936 259696 224942
rect 259644 224878 259696 224884
rect 260104 223440 260156 223446
rect 260104 223382 260156 223388
rect 258540 219156 258592 219162
rect 258540 219098 258592 219104
rect 259276 219156 259328 219162
rect 259276 219098 259328 219104
rect 259460 219156 259512 219162
rect 259460 219098 259512 219104
rect 256022 217110 256096 217138
rect 256850 217246 256924 217274
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217246
rect 257678 216988 257706 217246
rect 258552 217138 258580 219098
rect 259276 219020 259328 219026
rect 259276 218962 259328 218968
rect 258506 217110 258580 217138
rect 259288 217138 259316 218962
rect 259472 218618 259500 219098
rect 259460 218612 259512 218618
rect 259460 218554 259512 218560
rect 260116 217138 260144 223382
rect 260300 222630 260328 231676
rect 260944 225350 260972 231676
rect 261392 230172 261444 230178
rect 261392 230114 261444 230120
rect 260932 225344 260984 225350
rect 260932 225286 260984 225292
rect 260288 222624 260340 222630
rect 260288 222566 260340 222572
rect 261024 222148 261076 222154
rect 261024 222090 261076 222096
rect 261036 217138 261064 222090
rect 261404 220930 261432 230114
rect 261588 229634 261616 231676
rect 261576 229628 261628 229634
rect 261576 229570 261628 229576
rect 262232 226778 262260 231676
rect 262220 226772 262272 226778
rect 262220 226714 262272 226720
rect 261852 224392 261904 224398
rect 261852 224334 261904 224340
rect 261392 220924 261444 220930
rect 261392 220866 261444 220872
rect 261864 217138 261892 224334
rect 262876 222766 262904 231676
rect 263060 231662 263534 231690
rect 263888 231662 264178 231690
rect 262864 222760 262916 222766
rect 262864 222702 262916 222708
rect 263060 220114 263088 231662
rect 263888 224670 263916 231662
rect 264808 226166 264836 231676
rect 265176 231662 265466 231690
rect 265728 231662 266110 231690
rect 264796 226160 264848 226166
rect 264796 226102 264848 226108
rect 264152 224936 264204 224942
rect 264152 224878 264204 224884
rect 263876 224664 263928 224670
rect 263876 224606 263928 224612
rect 263508 222760 263560 222766
rect 263508 222702 263560 222708
rect 263048 220108 263100 220114
rect 263048 220050 263100 220056
rect 263324 220108 263376 220114
rect 263324 220050 263376 220056
rect 262680 218068 262732 218074
rect 262680 218010 262732 218016
rect 262692 217138 262720 218010
rect 263336 217274 263364 220050
rect 263520 218090 263548 222702
rect 264164 218754 264192 224878
rect 264796 223304 264848 223310
rect 264796 223246 264848 223252
rect 264152 218748 264204 218754
rect 264152 218690 264204 218696
rect 263520 218074 263640 218090
rect 264808 218074 264836 223246
rect 265176 220250 265204 231662
rect 265728 221338 265756 231662
rect 266740 226506 266768 231676
rect 267384 228546 267412 231676
rect 267372 228540 267424 228546
rect 267372 228482 267424 228488
rect 267556 228540 267608 228546
rect 267556 228482 267608 228488
rect 266728 226500 266780 226506
rect 266728 226442 266780 226448
rect 266268 226160 266320 226166
rect 266268 226102 266320 226108
rect 265716 221332 265768 221338
rect 265716 221274 265768 221280
rect 265164 220244 265216 220250
rect 265164 220186 265216 220192
rect 265992 218748 266044 218754
rect 265992 218690 266044 218696
rect 263520 218068 263652 218074
rect 263520 218062 263600 218068
rect 263600 218010 263652 218016
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263336 217246 263502 217274
rect 259288 217110 259362 217138
rect 260116 217110 260190 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217110
rect 260162 216988 260190 217110
rect 260990 217110 261064 217138
rect 261818 217110 261892 217138
rect 262646 217110 262720 217138
rect 260990 216988 261018 217110
rect 261818 216988 261846 217110
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217274 266032 218690
rect 266280 218074 266308 226102
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266820 218068 266872 218074
rect 266820 218010 266872 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217246 266032 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217246
rect 266832 217138 266860 218010
rect 267568 217274 267596 228482
rect 267694 226024 267746 226030
rect 267660 225972 267694 225978
rect 267660 225966 267746 225972
rect 267660 225950 267734 225966
rect 267660 218090 267688 225950
rect 268028 222358 268056 231676
rect 268672 222494 268700 231676
rect 269316 224942 269344 231676
rect 269960 226642 269988 231676
rect 270132 227724 270184 227730
rect 270132 227666 270184 227672
rect 269948 226636 270000 226642
rect 269948 226578 270000 226584
rect 269304 224936 269356 224942
rect 269304 224878 269356 224884
rect 269028 223576 269080 223582
rect 269028 223518 269080 223524
rect 268660 222488 268712 222494
rect 268660 222430 268712 222436
rect 268016 222352 268068 222358
rect 268016 222294 268068 222300
rect 267832 221876 267884 221882
rect 267832 221818 267884 221824
rect 267844 218618 267872 221818
rect 267832 218612 267884 218618
rect 267832 218554 267884 218560
rect 267660 218074 267734 218090
rect 269040 218074 269068 223518
rect 269304 218204 269356 218210
rect 269304 218146 269356 218152
rect 267660 218068 267746 218074
rect 267660 218062 267694 218068
rect 267694 218010 267746 218016
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 269028 218068 269080 218074
rect 269028 218010 269080 218016
rect 267568 217246 267642 217274
rect 266786 217110 266860 217138
rect 266786 216988 266814 217110
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218146
rect 270144 217274 270172 227666
rect 270604 225078 270632 231676
rect 271248 227050 271276 231676
rect 271892 230450 271920 231676
rect 271880 230444 271932 230450
rect 271880 230386 271932 230392
rect 272536 228002 272564 231676
rect 272720 231662 273194 231690
rect 272524 227996 272576 228002
rect 272524 227938 272576 227944
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 225072 270644 225078
rect 270592 225014 270644 225020
rect 271604 224664 271656 224670
rect 271604 224606 271656 224612
rect 270776 219564 270828 219570
rect 270776 219506 270828 219512
rect 270788 219298 270816 219506
rect 270776 219292 270828 219298
rect 270776 219234 270828 219240
rect 271616 218074 271644 224606
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 271604 218068 271656 218074
rect 271604 218010 271656 218016
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 270098 217246 270172 217274
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272432 226908 272484 226914
rect 272432 226850 272484 226856
rect 272444 218482 272472 226850
rect 272720 221746 272748 231662
rect 273824 228410 273852 231676
rect 274008 231662 274482 231690
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274008 221882 274036 231662
rect 274180 230444 274232 230450
rect 274180 230386 274232 230392
rect 273996 221876 274048 221882
rect 273996 221818 274048 221824
rect 272708 221740 272760 221746
rect 272708 221682 272760 221688
rect 273444 221332 273496 221338
rect 273444 221274 273496 221280
rect 272616 218612 272668 218618
rect 272616 218554 272668 218560
rect 272432 218476 272484 218482
rect 272432 218418 272484 218424
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272628 217138 272656 218554
rect 273456 217274 273484 221274
rect 274192 219434 274220 230386
rect 275112 226302 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 226296 275152 226302
rect 275100 226238 275152 226244
rect 275296 221746 275324 231662
rect 275836 225004 275888 225010
rect 275836 224946 275888 224952
rect 275284 221740 275336 221746
rect 275284 221682 275336 221688
rect 275100 221604 275152 221610
rect 275100 221546 275152 221552
rect 273916 219406 274220 219434
rect 273916 218210 273944 219406
rect 274272 218884 274324 218890
rect 274272 218826 274324 218832
rect 273904 218204 273956 218210
rect 273904 218146 273956 218152
rect 272582 217110 272656 217138
rect 273410 217246 273484 217274
rect 272582 216988 272610 217110
rect 273410 216988 273438 217246
rect 274284 217138 274312 218826
rect 275112 217274 275140 221546
rect 274238 217110 274312 217138
rect 275066 217246 275140 217274
rect 275848 217274 275876 224946
rect 276124 220386 276152 231662
rect 276296 230308 276348 230314
rect 276296 230250 276348 230256
rect 276308 225010 276336 230250
rect 277044 229498 277072 231676
rect 277032 229492 277084 229498
rect 277032 229434 277084 229440
rect 277216 228268 277268 228274
rect 277216 228210 277268 228216
rect 276296 225004 276348 225010
rect 276296 224946 276348 224952
rect 276112 220380 276164 220386
rect 276112 220322 276164 220328
rect 277228 218074 277256 228210
rect 277688 222902 277716 231676
rect 278332 227322 278360 231676
rect 278320 227316 278372 227322
rect 278320 227258 278372 227264
rect 278504 226296 278556 226302
rect 278504 226238 278556 226244
rect 277676 222896 277728 222902
rect 277676 222838 277728 222844
rect 278320 221740 278372 221746
rect 278320 221682 278372 221688
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 274238 216988 274266 217110
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278332 217274 278360 221682
rect 278516 218074 278544 226238
rect 278976 224126 279004 231676
rect 279252 231662 279634 231690
rect 278964 224120 279016 224126
rect 278964 224062 279016 224068
rect 279252 219570 279280 231662
rect 280264 227186 280292 231676
rect 280448 231662 280922 231690
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 280448 221066 280476 231662
rect 280712 227316 280764 227322
rect 280712 227258 280764 227264
rect 280436 221060 280488 221066
rect 280436 221002 280488 221008
rect 280068 220380 280120 220386
rect 280068 220322 280120 220328
rect 279240 219564 279292 219570
rect 279240 219506 279292 219512
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278504 218068 278556 218074
rect 278504 218010 278556 218016
rect 278332 217246 278406 217274
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 220322
rect 280724 218890 280752 227258
rect 281552 225622 281580 231676
rect 282196 229770 282224 231676
rect 282184 229764 282236 229770
rect 282184 229706 282236 229712
rect 282840 229094 282868 231676
rect 282380 229066 282868 229094
rect 283024 231662 283498 231690
rect 281540 225616 281592 225622
rect 281540 225558 281592 225564
rect 282380 223990 282408 229066
rect 282736 225004 282788 225010
rect 282736 224946 282788 224952
rect 282552 224800 282604 224806
rect 282552 224742 282604 224748
rect 282368 223984 282420 223990
rect 282368 223926 282420 223932
rect 280896 220244 280948 220250
rect 280896 220186 280948 220192
rect 280712 218884 280764 218890
rect 280712 218826 280764 218832
rect 280908 217274 280936 220186
rect 281080 218884 281132 218890
rect 281080 218826 281132 218832
rect 281092 218482 281120 218826
rect 281080 218476 281132 218482
rect 281080 218418 281132 218424
rect 282564 218074 282592 224742
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282552 218068 282604 218074
rect 282552 218010 282604 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 280862 217246 280936 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280862 216988 280890 217246
rect 281736 217138 281764 218010
rect 282748 217274 282776 224946
rect 283024 220658 283052 231662
rect 284128 228682 284156 231676
rect 284116 228676 284168 228682
rect 284116 228618 284168 228624
rect 284116 228404 284168 228410
rect 284116 228346 284168 228352
rect 283380 222896 283432 222902
rect 283380 222838 283432 222844
rect 283012 220652 283064 220658
rect 283012 220594 283064 220600
rect 283392 217274 283420 222838
rect 281690 217110 281764 217138
rect 282518 217246 282776 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 228346
rect 284772 226914 284800 231676
rect 285048 231662 285430 231690
rect 285968 231662 286074 231690
rect 286336 231662 286718 231690
rect 284760 226908 284812 226914
rect 284760 226850 284812 226856
rect 285048 223854 285076 231662
rect 285312 229764 285364 229770
rect 285312 229706 285364 229712
rect 285324 225010 285352 229706
rect 285496 225616 285548 225622
rect 285496 225558 285548 225564
rect 285312 225004 285364 225010
rect 285312 224946 285364 224952
rect 285036 223848 285088 223854
rect 285036 223790 285088 223796
rect 285508 218074 285536 225558
rect 285968 222018 285996 231662
rect 285956 222012 286008 222018
rect 285956 221954 286008 221960
rect 286336 221882 286364 231662
rect 287348 229906 287376 231676
rect 287624 231662 288006 231690
rect 287336 229900 287388 229906
rect 287336 229842 287388 229848
rect 286692 224120 286744 224126
rect 286692 224062 286744 224068
rect 285680 221876 285732 221882
rect 285680 221818 285732 221824
rect 286324 221876 286376 221882
rect 286324 221818 286376 221824
rect 285692 221474 285720 221818
rect 285680 221468 285732 221474
rect 285680 221410 285732 221416
rect 285956 221468 286008 221474
rect 285956 221410 286008 221416
rect 285968 219434 285996 221410
rect 285956 219428 286008 219434
rect 285956 219370 286008 219376
rect 285864 218476 285916 218482
rect 285864 218418 285916 218424
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 218418
rect 286704 217274 286732 224062
rect 287624 223174 287652 231662
rect 288164 228132 288216 228138
rect 288164 228074 288216 228080
rect 287612 223168 287664 223174
rect 287612 223110 287664 223116
rect 288176 219434 288204 228074
rect 288348 224936 288400 224942
rect 288348 224878 288400 224884
rect 288360 219434 288388 224878
rect 288636 224262 288664 231676
rect 289280 224534 289308 231676
rect 289924 229094 289952 231676
rect 289832 229066 289952 229094
rect 289268 224528 289320 224534
rect 289268 224470 289320 224476
rect 288624 224256 288676 224262
rect 288624 224198 288676 224204
rect 289636 224256 289688 224262
rect 289636 224198 289688 224204
rect 287520 219428 287572 219434
rect 288176 219406 288296 219434
rect 288360 219428 288492 219434
rect 288360 219406 288440 219428
rect 287520 219370 287572 219376
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 219370
rect 288268 217274 288296 219406
rect 288440 219370 288492 219376
rect 289648 218074 289676 224198
rect 289832 221474 289860 229066
rect 290568 225894 290596 231676
rect 291212 228954 291240 231676
rect 291200 228948 291252 228954
rect 291200 228890 291252 228896
rect 291856 227458 291884 231676
rect 292500 230042 292528 231676
rect 292488 230036 292540 230042
rect 292488 229978 292540 229984
rect 292396 228676 292448 228682
rect 292396 228618 292448 228624
rect 291844 227452 291896 227458
rect 291844 227394 291896 227400
rect 291844 226432 291896 226438
rect 291844 226374 291896 226380
rect 290556 225888 290608 225894
rect 290556 225830 290608 225836
rect 290832 223168 290884 223174
rect 290832 223110 290884 223116
rect 289820 221468 289872 221474
rect 289820 221410 289872 221416
rect 290004 221468 290056 221474
rect 290004 221410 290056 221416
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289636 218068 289688 218074
rect 289636 218010 289688 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217274 290044 221410
rect 290844 217274 290872 223110
rect 291660 219428 291712 219434
rect 291660 219370 291712 219376
rect 289142 217110 289216 217138
rect 289970 217246 290044 217274
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217246
rect 290798 216988 290826 217246
rect 291672 217138 291700 219370
rect 291856 219162 291884 226374
rect 291844 219156 291896 219162
rect 291844 219098 291896 219104
rect 292408 217274 292436 228618
rect 293144 227594 293172 231676
rect 293328 231662 293802 231690
rect 293132 227588 293184 227594
rect 293132 227530 293184 227536
rect 293328 220794 293356 231662
rect 293776 227452 293828 227458
rect 293776 227394 293828 227400
rect 293316 220788 293368 220794
rect 293316 220730 293368 220736
rect 293592 219836 293644 219842
rect 293592 219778 293644 219784
rect 293604 219026 293632 219778
rect 293592 219020 293644 219026
rect 293592 218962 293644 218968
rect 293788 218074 293816 227394
rect 294432 223038 294460 231676
rect 295076 226438 295104 231676
rect 295720 228818 295748 231676
rect 295904 231662 296378 231690
rect 296824 231662 297022 231690
rect 295708 228812 295760 228818
rect 295708 228754 295760 228760
rect 295064 226432 295116 226438
rect 295064 226374 295116 226380
rect 294972 225888 295024 225894
rect 294972 225830 295024 225836
rect 294420 223032 294472 223038
rect 294420 222974 294472 222980
rect 294144 219156 294196 219162
rect 294144 219098 294196 219104
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 292408 217246 292482 217274
rect 291626 217110 291700 217138
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 219098
rect 294984 217274 295012 225830
rect 295904 219978 295932 231662
rect 296444 227180 296496 227186
rect 296444 227122 296496 227128
rect 295892 219972 295944 219978
rect 295892 219914 295944 219920
rect 296456 218074 296484 227122
rect 296628 220652 296680 220658
rect 296628 220594 296680 220600
rect 295800 218068 295852 218074
rect 295800 218010 295852 218016
rect 296444 218068 296496 218074
rect 296444 218010 296496 218016
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 218010
rect 296640 217274 296668 220594
rect 296824 220522 296852 231662
rect 297652 230178 297680 231676
rect 297640 230172 297692 230178
rect 297640 230114 297692 230120
rect 296996 230036 297048 230042
rect 296996 229978 297048 229984
rect 297008 222766 297036 229978
rect 298296 229090 298324 231676
rect 298284 229084 298336 229090
rect 298284 229026 298336 229032
rect 298008 223576 298060 223582
rect 298008 223518 298060 223524
rect 296996 222760 297048 222766
rect 296996 222702 297048 222708
rect 296996 220788 297048 220794
rect 296996 220730 297048 220736
rect 296812 220516 296864 220522
rect 296812 220458 296864 220464
rect 297008 218618 297036 220730
rect 296996 218612 297048 218618
rect 296996 218554 297048 218560
rect 298020 218074 298048 223518
rect 298940 223446 298968 231676
rect 299296 227588 299348 227594
rect 299296 227530 299348 227536
rect 298928 223440 298980 223446
rect 298928 223382 298980 223388
rect 299112 218204 299164 218210
rect 299112 218146 299164 218152
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 298008 218068 298060 218074
rect 298008 218010 298060 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 295766 217110 295840 217138
rect 296594 217246 296668 217274
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299124 217138 299152 218146
rect 299308 218074 299336 227530
rect 299584 225758 299612 231676
rect 299952 231662 300242 231690
rect 299952 229094 299980 231662
rect 300124 229900 300176 229906
rect 300124 229842 300176 229848
rect 299768 229066 299980 229094
rect 299572 225752 299624 225758
rect 299572 225694 299624 225700
rect 299768 219842 299796 229066
rect 300136 223582 300164 229842
rect 300872 224398 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 302528 231662 302818 231690
rect 300860 224392 300912 224398
rect 300860 224334 300912 224340
rect 300124 223576 300176 223582
rect 300124 223518 300176 223524
rect 300308 223032 300360 223038
rect 300308 222974 300360 222980
rect 299940 220516 299992 220522
rect 299940 220458 299992 220464
rect 299756 219836 299808 219842
rect 299756 219778 299808 219784
rect 299296 218068 299348 218074
rect 299296 218010 299348 218016
rect 299952 217274 299980 220458
rect 300320 218210 300348 222974
rect 301056 220114 301084 231662
rect 301700 222154 301728 231662
rect 302528 230042 302556 231662
rect 302884 230104 302936 230110
rect 302884 230046 302936 230052
rect 302516 230036 302568 230042
rect 302516 229978 302568 229984
rect 302148 223440 302200 223446
rect 302148 223382 302200 223388
rect 301688 222148 301740 222154
rect 301688 222090 301740 222096
rect 301044 220108 301096 220114
rect 301044 220050 301096 220056
rect 300768 219020 300820 219026
rect 300768 218962 300820 218968
rect 300308 218204 300360 218210
rect 300308 218146 300360 218152
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217110 299152 217138
rect 299906 217246 299980 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217110
rect 299906 216988 299934 217246
rect 300780 217138 300808 218962
rect 302160 218074 302188 223382
rect 302896 218754 302924 230046
rect 303448 226166 303476 231676
rect 303436 226160 303488 226166
rect 303436 226102 303488 226108
rect 304092 226030 304120 231676
rect 304080 226024 304132 226030
rect 304080 225966 304132 225972
rect 303252 224392 303304 224398
rect 303252 224334 303304 224340
rect 302884 218748 302936 218754
rect 302884 218690 302936 218696
rect 302424 218204 302476 218210
rect 302424 218146 302476 218152
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 301608 217138 301636 218010
rect 302436 217138 302464 218146
rect 303264 217274 303292 224334
rect 304736 223310 304764 231676
rect 305380 230110 305408 231676
rect 305368 230104 305420 230110
rect 305368 230046 305420 230052
rect 305644 230036 305696 230042
rect 305644 229978 305696 229984
rect 304908 225752 304960 225758
rect 304908 225694 304960 225700
rect 304724 223304 304776 223310
rect 304724 223246 304776 223252
rect 304632 221876 304684 221882
rect 304632 221818 304684 221824
rect 304644 218210 304672 221818
rect 304632 218204 304684 218210
rect 304632 218146 304684 218152
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 300734 217110 300808 217138
rect 301562 217110 301636 217138
rect 302390 217110 302464 217138
rect 303218 217246 303292 217274
rect 300734 216988 300762 217110
rect 301562 216988 301590 217110
rect 302390 216988 302418 217110
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 225694
rect 305656 219434 305684 229978
rect 306024 223582 306052 231676
rect 306668 227730 306696 231676
rect 307312 228546 307340 231676
rect 307956 230450 307984 231676
rect 307944 230444 307996 230450
rect 307944 230386 307996 230392
rect 308128 230172 308180 230178
rect 308128 230114 308180 230120
rect 307300 228540 307352 228546
rect 307300 228482 307352 228488
rect 307668 228540 307720 228546
rect 307668 228482 307720 228488
rect 306656 227724 306708 227730
rect 306656 227666 306708 227672
rect 306012 223576 306064 223582
rect 306012 223518 306064 223524
rect 306288 223304 306340 223310
rect 306288 223246 306340 223252
rect 305564 219406 305684 219434
rect 305564 218074 305592 219406
rect 306300 218074 306328 223246
rect 306748 219972 306800 219978
rect 306748 219914 306800 219920
rect 306760 218482 306788 219914
rect 307392 218748 307444 218754
rect 307392 218690 307444 218696
rect 306748 218476 306800 218482
rect 306748 218418 306800 218424
rect 305552 218068 305604 218074
rect 305552 218010 305604 218016
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306288 218068 306340 218074
rect 306288 218010 306340 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218690
rect 307680 218074 307708 228482
rect 308140 224262 308168 230114
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308772 227044 308824 227050
rect 308772 226986 308824 226992
rect 308128 224256 308180 224262
rect 308128 224198 308180 224204
rect 308784 218074 308812 226986
rect 308956 224256 309008 224262
rect 308956 224198 309008 224204
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308772 218068 308824 218074
rect 308772 218010 308824 218016
rect 308232 217138 308260 218010
rect 308968 217274 308996 224198
rect 309244 221338 309272 231676
rect 309888 224670 309916 231676
rect 310546 231662 310744 231690
rect 309876 224664 309928 224670
rect 309876 224606 309928 224612
rect 309876 222012 309928 222018
rect 309876 221954 309928 221960
rect 309232 221332 309284 221338
rect 309232 221274 309284 221280
rect 309888 217274 309916 221954
rect 310716 220794 310744 231662
rect 310900 231662 311190 231690
rect 310900 221610 310928 231662
rect 311820 228274 311848 231676
rect 312096 231662 312478 231690
rect 311808 228268 311860 228274
rect 311808 228210 311860 228216
rect 312096 227322 312124 231662
rect 312544 230444 312596 230450
rect 312544 230386 312596 230392
rect 312084 227316 312136 227322
rect 312084 227258 312136 227264
rect 311532 222148 311584 222154
rect 311532 222090 311584 222096
rect 310888 221604 310940 221610
rect 310888 221546 310940 221552
rect 310704 220788 310756 220794
rect 310704 220730 310756 220736
rect 310704 218204 310756 218210
rect 310704 218146 310756 218152
rect 308968 217246 309042 217274
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309842 217246 309916 217274
rect 309842 216988 309870 217246
rect 310716 217138 310744 218146
rect 311544 217274 311572 222090
rect 311808 220788 311860 220794
rect 311808 220730 311860 220736
rect 311820 219162 311848 220730
rect 311808 219156 311860 219162
rect 311808 219098 311860 219104
rect 312556 218890 312584 230386
rect 313108 230314 313136 231676
rect 313476 231662 313766 231690
rect 314120 231662 314410 231690
rect 313096 230308 313148 230314
rect 313096 230250 313148 230256
rect 313096 226024 313148 226030
rect 313096 225966 313148 225972
rect 312544 218884 312596 218890
rect 312544 218826 312596 218832
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 310670 217110 310744 217138
rect 311498 217246 311572 217274
rect 310670 216988 310698 217110
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313108 217274 313136 225966
rect 313476 221746 313504 231662
rect 313464 221740 313516 221746
rect 313464 221682 313516 221688
rect 314120 220386 314148 231662
rect 315040 226302 315068 231676
rect 315684 230450 315712 231676
rect 315672 230444 315724 230450
rect 315672 230386 315724 230392
rect 315304 230172 315356 230178
rect 315304 230114 315356 230120
rect 315028 226296 315080 226302
rect 315028 226238 315080 226244
rect 314568 221604 314620 221610
rect 314568 221546 314620 221552
rect 314108 220380 314160 220386
rect 314108 220322 314160 220328
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 313108 217246 313182 217274
rect 312326 217110 312400 217138
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 314580 218074 314608 221546
rect 315316 218210 315344 230114
rect 316328 224806 316356 231676
rect 316316 224800 316368 224806
rect 316316 224742 316368 224748
rect 315856 224664 315908 224670
rect 315856 224606 315908 224612
rect 315672 219156 315724 219162
rect 315672 219098 315724 219104
rect 315304 218204 315356 218210
rect 315304 218146 315356 218152
rect 314568 218068 314620 218074
rect 314568 218010 314620 218016
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 314856 217138 314884 218010
rect 315684 217138 315712 219098
rect 315868 218074 315896 224606
rect 316972 222902 317000 231676
rect 317524 231662 317630 231690
rect 317328 226296 317380 226302
rect 317328 226238 317380 226244
rect 316960 222896 317012 222902
rect 316960 222838 317012 222844
rect 317144 222896 317196 222902
rect 317144 222838 317196 222844
rect 317156 218074 317184 222838
rect 315856 218068 315908 218074
rect 315856 218010 315908 218016
rect 316500 218068 316552 218074
rect 316500 218010 316552 218016
rect 317144 218068 317196 218074
rect 317144 218010 317196 218016
rect 316512 217138 316540 218010
rect 317340 217274 317368 226238
rect 317524 220250 317552 231662
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 317972 228812 318024 228818
rect 317972 228754 318024 228760
rect 317512 220244 317564 220250
rect 317512 220186 317564 220192
rect 317984 219162 318012 228754
rect 318904 225622 318932 231676
rect 318892 225616 318944 225622
rect 318892 225558 318944 225564
rect 319548 224126 319576 231676
rect 319812 228948 319864 228954
rect 319812 228890 319864 228896
rect 319536 224120 319588 224126
rect 319536 224062 319588 224068
rect 318156 220108 318208 220114
rect 318156 220050 318208 220056
rect 317972 219156 318024 219162
rect 317972 219098 318024 219104
rect 318168 217274 318196 220050
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217110 315712 217138
rect 316466 217110 316540 217138
rect 317294 217246 317368 217274
rect 318122 217246 318196 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217110
rect 316466 216988 316494 217110
rect 317294 216988 317322 217246
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 228890
rect 320192 228410 320220 231676
rect 320376 231662 320850 231690
rect 320180 228404 320232 228410
rect 320180 228346 320232 228352
rect 319996 224528 320048 224534
rect 319996 224470 320048 224476
rect 320008 218074 320036 224470
rect 320376 219978 320404 231662
rect 321480 228138 321508 231676
rect 321756 231662 322138 231690
rect 322400 231662 322782 231690
rect 321468 228132 321520 228138
rect 321468 228074 321520 228080
rect 321376 227724 321428 227730
rect 321376 227666 321428 227672
rect 320364 219972 320416 219978
rect 320364 219914 320416 219920
rect 320640 219156 320692 219162
rect 320640 219098 320692 219104
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219098
rect 321388 217274 321416 227666
rect 321756 221474 321784 231662
rect 322400 224942 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 225616 322900 225622
rect 322848 225558 322900 225564
rect 322388 224936 322440 224942
rect 322388 224878 322440 224884
rect 321744 221468 321796 221474
rect 321744 221410 321796 221416
rect 322860 218074 322888 225558
rect 323688 223174 323716 231662
rect 324044 229764 324096 229770
rect 324044 229706 324096 229712
rect 323676 223168 323728 223174
rect 323676 223110 323728 223116
rect 323124 220380 323176 220386
rect 323124 220322 323176 220328
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217274 323164 220322
rect 324056 219434 324084 229706
rect 324700 219434 324728 231676
rect 325344 227458 325372 231676
rect 325332 227452 325384 227458
rect 325332 227394 325384 227400
rect 325424 226160 325476 226166
rect 325424 226102 325476 226108
rect 323964 219406 324084 219434
rect 324688 219428 324740 219434
rect 323964 217274 323992 219406
rect 324688 219370 324740 219376
rect 325436 218074 325464 226102
rect 325988 225894 326016 231676
rect 326632 228682 326660 231676
rect 327092 231662 327290 231690
rect 327460 231662 327934 231690
rect 326620 228676 326672 228682
rect 326620 228618 326672 228624
rect 326896 228404 326948 228410
rect 326896 228346 326948 228352
rect 326344 227316 326396 227322
rect 326344 227258 326396 227264
rect 325976 225888 326028 225894
rect 325976 225830 326028 225836
rect 326356 219434 326384 227258
rect 325608 219428 325660 219434
rect 325608 219370 325660 219376
rect 326344 219428 326396 219434
rect 326344 219370 326396 219376
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217246 323164 217274
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217246
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217138 325648 219370
rect 326908 218074 326936 228346
rect 327092 220794 327120 231662
rect 327080 220788 327132 220794
rect 327080 220730 327132 220736
rect 327460 220658 327488 231662
rect 328564 227594 328592 231676
rect 328552 227588 328604 227594
rect 328552 227530 328604 227536
rect 329208 227186 329236 231676
rect 329852 229906 329880 231676
rect 330036 231662 330510 231690
rect 329840 229900 329892 229906
rect 329840 229842 329892 229848
rect 329196 227180 329248 227186
rect 329196 227122 329248 227128
rect 329748 227180 329800 227186
rect 329748 227122 329800 227128
rect 329104 223576 329156 223582
rect 329104 223518 329156 223524
rect 327448 220652 327500 220658
rect 327448 220594 327500 220600
rect 328092 220652 328144 220658
rect 328092 220594 328144 220600
rect 327264 219292 327316 219298
rect 327264 219234 327316 219240
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 326448 217138 326476 218010
rect 327276 217274 327304 219234
rect 328104 217274 328132 220594
rect 329116 218890 329144 223518
rect 329288 220788 329340 220794
rect 329288 220730 329340 220736
rect 329300 219026 329328 220730
rect 329288 219020 329340 219026
rect 329288 218962 329340 218968
rect 329104 218884 329156 218890
rect 329104 218826 329156 218832
rect 328920 218068 328972 218074
rect 328920 218010 328972 218016
rect 324746 217110 324820 217138
rect 325574 217110 325648 217138
rect 326402 217110 326476 217138
rect 327230 217246 327304 217274
rect 328058 217246 328132 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217110
rect 326402 216988 326430 217110
rect 327230 216988 327258 217246
rect 328058 216988 328086 217246
rect 328932 217138 328960 218010
rect 329760 217274 329788 227122
rect 330036 220522 330064 231662
rect 331140 223446 331168 231676
rect 331128 223440 331180 223446
rect 331128 223382 331180 223388
rect 330484 223168 330536 223174
rect 330484 223110 330536 223116
rect 330024 220516 330076 220522
rect 330024 220458 330076 220464
rect 330496 218074 330524 223110
rect 331784 223038 331812 231676
rect 331968 231662 332442 231690
rect 331772 223032 331824 223038
rect 331772 222974 331824 222980
rect 331404 221740 331456 221746
rect 331404 221682 331456 221688
rect 330668 218204 330720 218210
rect 330668 218146 330720 218152
rect 330484 218068 330536 218074
rect 330484 218010 330536 218016
rect 330680 217274 330708 218146
rect 331416 217274 331444 221682
rect 331968 220794 331996 231662
rect 333072 224398 333100 231676
rect 333244 228676 333296 228682
rect 333244 228618 333296 228624
rect 333060 224392 333112 224398
rect 333060 224334 333112 224340
rect 331956 220788 332008 220794
rect 331956 220730 332008 220736
rect 332232 220244 332284 220250
rect 332232 220186 332284 220192
rect 332244 217274 332272 220186
rect 333256 218210 333284 228618
rect 333716 225758 333744 231676
rect 334084 231662 334374 231690
rect 333704 225752 333756 225758
rect 333704 225694 333756 225700
rect 333888 224392 333940 224398
rect 333888 224334 333940 224340
rect 333704 219020 333756 219026
rect 333704 218962 333756 218968
rect 333244 218204 333296 218210
rect 333244 218146 333296 218152
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 330542 217246 330708 217274
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330542 216988 330570 217246
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 218962
rect 333900 218074 333928 224334
rect 334084 221882 334112 231662
rect 335004 230042 335032 231676
rect 334992 230036 335044 230042
rect 334992 229978 335044 229984
rect 334256 229900 334308 229906
rect 334256 229842 334308 229848
rect 334268 226302 334296 229842
rect 335648 228546 335676 231676
rect 335636 228540 335688 228546
rect 335636 228482 335688 228488
rect 336292 227050 336320 231676
rect 336648 228540 336700 228546
rect 336648 228482 336700 228488
rect 336280 227044 336332 227050
rect 336280 226986 336332 226992
rect 336464 227044 336516 227050
rect 336464 226986 336516 226992
rect 334256 226296 334308 226302
rect 334256 226238 334308 226244
rect 335268 225752 335320 225758
rect 335268 225694 335320 225700
rect 334072 221876 334124 221882
rect 334072 221818 334124 221824
rect 335280 218074 335308 225694
rect 336476 219434 336504 226986
rect 336660 219434 336688 228482
rect 336936 223310 336964 231676
rect 337120 231662 337594 231690
rect 336924 223304 336976 223310
rect 336924 223246 336976 223252
rect 337120 219434 337148 231662
rect 337936 223032 337988 223038
rect 337936 222974 337988 222980
rect 336384 219406 336504 219434
rect 336568 219406 336688 219434
rect 337028 219406 337148 219434
rect 336384 218074 336412 219406
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335268 218068 335320 218074
rect 335268 218010 335320 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 336372 218068 336424 218074
rect 336372 218010 336424 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336568 217274 336596 219406
rect 337028 218754 337056 219406
rect 337200 218884 337252 218890
rect 337200 218826 337252 218832
rect 337016 218748 337068 218754
rect 337016 218690 337068 218696
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336596 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218826
rect 337948 217274 337976 222974
rect 338224 222018 338252 231676
rect 338408 231662 338882 231690
rect 338408 222154 338436 231662
rect 339512 224262 339540 231676
rect 340156 230178 340184 231676
rect 340144 230172 340196 230178
rect 340144 230114 340196 230120
rect 340604 227452 340656 227458
rect 340604 227394 340656 227400
rect 340144 225888 340196 225894
rect 340144 225830 340196 225836
rect 339500 224256 339552 224262
rect 339500 224198 339552 224204
rect 338396 222148 338448 222154
rect 338396 222090 338448 222096
rect 338212 222012 338264 222018
rect 338212 221954 338264 221960
rect 338856 221468 338908 221474
rect 338856 221410 338908 221416
rect 338868 217274 338896 221410
rect 340156 219162 340184 225830
rect 340616 219434 340644 227394
rect 340800 226030 340828 231676
rect 340788 226024 340840 226030
rect 340788 225966 340840 225972
rect 341444 224670 341472 231676
rect 341628 231662 342102 231690
rect 341432 224664 341484 224670
rect 341432 224606 341484 224612
rect 341628 221950 341656 231662
rect 342076 224256 342128 224262
rect 342076 224198 342128 224204
rect 340880 221944 340932 221950
rect 340880 221886 340932 221892
rect 341616 221944 341668 221950
rect 341616 221886 341668 221892
rect 340892 221610 340920 221886
rect 340880 221604 340932 221610
rect 340880 221546 340932 221552
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 340616 219406 340736 219434
rect 340144 219156 340196 219162
rect 340144 219098 340196 219104
rect 340512 218748 340564 218754
rect 340512 218690 340564 218696
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338822 217246 338896 217274
rect 338822 216988 338850 217246
rect 339696 217138 339724 218010
rect 340524 217274 340552 218690
rect 340708 218074 340736 219406
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 339650 217110 339724 217138
rect 340478 217246 340552 217274
rect 341306 217246 341380 217274
rect 342088 217274 342116 224198
rect 342732 223582 342760 231676
rect 342720 223576 342772 223582
rect 342720 223518 342772 223524
rect 343376 222902 343404 231676
rect 343744 231662 344034 231690
rect 343548 223304 343600 223310
rect 343548 223246 343600 223252
rect 343364 222896 343416 222902
rect 343364 222838 343416 222844
rect 343560 218074 343588 223246
rect 343744 220114 343772 231662
rect 344664 228818 344692 231676
rect 345308 229906 345336 231676
rect 345664 230104 345716 230110
rect 345664 230046 345716 230052
rect 345296 229900 345348 229906
rect 345296 229842 345348 229848
rect 344652 228812 344704 228818
rect 344652 228754 344704 228760
rect 344652 224664 344704 224670
rect 344652 224606 344704 224612
rect 343732 220108 343784 220114
rect 343732 220050 343784 220056
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342996 218068 343048 218074
rect 342996 218010 343048 218016
rect 343548 218068 343600 218074
rect 343548 218010 343600 218016
rect 342088 217246 342162 217274
rect 339650 216988 339678 217110
rect 340478 216988 340506 217246
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 343008 217138 343036 218010
rect 343836 217138 343864 219370
rect 344664 217274 344692 224606
rect 345480 220108 345532 220114
rect 345480 220050 345532 220056
rect 345492 217274 345520 220050
rect 345676 219162 345704 230046
rect 345952 228954 345980 231676
rect 345940 228948 345992 228954
rect 345940 228890 345992 228896
rect 346216 228812 346268 228818
rect 346216 228754 346268 228760
rect 345664 219156 345716 219162
rect 345664 219098 345716 219104
rect 342962 217110 343036 217138
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 345446 217246 345520 217274
rect 346228 217274 346256 228754
rect 346596 227730 346624 231676
rect 346584 227724 346636 227730
rect 346584 227666 346636 227672
rect 347044 225888 347096 225894
rect 347044 225830 347096 225836
rect 347056 219434 347084 225830
rect 347240 224534 347268 231676
rect 347884 226030 347912 231676
rect 348160 231662 348542 231690
rect 347872 226024 347924 226030
rect 347872 225966 347924 225972
rect 347228 224528 347280 224534
rect 347228 224470 347280 224476
rect 347596 222896 347648 222902
rect 347596 222838 347648 222844
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347608 218074 347636 222838
rect 348160 220386 348188 231662
rect 349172 226166 349200 231676
rect 349160 226160 349212 226166
rect 349160 226102 349212 226108
rect 349068 226024 349120 226030
rect 349068 225966 349120 225972
rect 348148 220380 348200 220386
rect 348148 220322 348200 220328
rect 348792 218204 348844 218210
rect 348792 218146 348844 218152
rect 347136 218068 347188 218074
rect 347136 218010 347188 218016
rect 347596 218068 347648 218074
rect 347596 218010 347648 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 342962 216988 342990 217110
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345446 216988 345474 217246
rect 346274 216988 346302 217246
rect 347148 217138 347176 218010
rect 347976 217138 348004 218010
rect 348804 217138 348832 218146
rect 349080 218074 349108 225966
rect 349816 225622 349844 231676
rect 350460 229770 350488 231676
rect 350448 229764 350500 229770
rect 350448 229706 350500 229712
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 350172 228948 350224 228954
rect 350172 228890 350224 228896
rect 349804 225616 349856 225622
rect 349804 225558 349856 225564
rect 350184 218074 350212 228890
rect 350552 225026 350580 229570
rect 351104 228410 351132 231676
rect 351288 231662 351762 231690
rect 351288 229094 351316 231662
rect 351288 229066 351408 229094
rect 351092 228404 351144 228410
rect 351092 228346 351144 228352
rect 351184 225616 351236 225622
rect 351184 225558 351236 225564
rect 350368 224998 350580 225026
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 349632 217138 349660 218010
rect 350368 217274 350396 224998
rect 351196 218210 351224 225558
rect 351380 220658 351408 229066
rect 352392 227322 352420 231676
rect 353036 230110 353064 231676
rect 353024 230104 353076 230110
rect 353024 230046 353076 230052
rect 352564 229900 352616 229906
rect 352564 229842 352616 229848
rect 352380 227316 352432 227322
rect 352380 227258 352432 227264
rect 351368 220652 351420 220658
rect 351368 220594 351420 220600
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 351368 219020 351420 219026
rect 351368 218962 351420 218968
rect 351184 218204 351236 218210
rect 351184 218146 351236 218152
rect 351380 217274 351408 218962
rect 350368 217246 350442 217274
rect 347102 217110 347176 217138
rect 347930 217110 348004 217138
rect 348758 217110 348832 217138
rect 349586 217110 349660 217138
rect 347102 216988 347130 217110
rect 347930 216988 347958 217110
rect 348758 216988 348786 217110
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351408 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352576 219162 352604 229842
rect 353680 227186 353708 231676
rect 353956 231662 354338 231690
rect 353668 227180 353720 227186
rect 353668 227122 353720 227128
rect 353956 221746 353984 231662
rect 354588 227180 354640 227186
rect 354588 227122 354640 227128
rect 353944 221740 353996 221746
rect 353944 221682 353996 221688
rect 352932 220380 352984 220386
rect 352932 220322 352984 220328
rect 352564 219156 352616 219162
rect 352564 219098 352616 219104
rect 352944 217274 352972 220322
rect 354404 219156 354456 219162
rect 354404 219098 354456 219104
rect 353760 218068 353812 218074
rect 353760 218010 353812 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218010
rect 354416 217274 354444 219098
rect 354600 218074 354628 227122
rect 354968 223174 354996 231676
rect 355612 228682 355640 231676
rect 355600 228676 355652 228682
rect 355600 228618 355652 228624
rect 355232 228404 355284 228410
rect 355232 228346 355284 228352
rect 354956 223168 355008 223174
rect 354956 223110 355008 223116
rect 355244 219026 355272 228346
rect 355508 226908 355560 226914
rect 355508 226850 355560 226856
rect 355520 219162 355548 226850
rect 356256 224398 356284 231676
rect 356900 225758 356928 231676
rect 356888 225752 356940 225758
rect 356888 225694 356940 225700
rect 356244 224392 356296 224398
rect 356244 224334 356296 224340
rect 357348 224392 357400 224398
rect 357348 224334 357400 224340
rect 357072 223168 357124 223174
rect 357072 223110 357124 223116
rect 355508 219156 355560 219162
rect 355508 219098 355560 219104
rect 355232 219020 355284 219026
rect 355232 218962 355284 218968
rect 355416 219020 355468 219026
rect 355416 218962 355468 218968
rect 354588 218068 354640 218074
rect 354588 218010 354640 218016
rect 354416 217246 354582 217274
rect 353726 217110 353800 217138
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218962
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356256 217138 356284 218010
rect 357084 217274 357112 223110
rect 357360 218074 357388 224334
rect 357544 220250 357572 231676
rect 358188 229906 358216 231676
rect 358176 229900 358228 229906
rect 358176 229842 358228 229848
rect 358084 229288 358136 229294
rect 358084 229230 358136 229236
rect 357532 220244 357584 220250
rect 357532 220186 357584 220192
rect 358096 219434 358124 229230
rect 358832 228546 358860 231676
rect 359200 231662 359490 231690
rect 358820 228540 358872 228546
rect 358820 228482 358872 228488
rect 359200 223038 359228 231662
rect 359372 227588 359424 227594
rect 359372 227530 359424 227536
rect 359188 223032 359240 223038
rect 359188 222974 359240 222980
rect 357728 219406 358124 219434
rect 357728 218890 357756 219406
rect 358728 219156 358780 219162
rect 358728 219098 358780 219104
rect 357716 218884 357768 218890
rect 357716 218826 357768 218832
rect 357348 218068 357400 218074
rect 357348 218010 357400 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357112 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357912 217138 357940 218010
rect 358740 217138 358768 219098
rect 359384 218074 359412 227530
rect 360120 227050 360148 231676
rect 360764 229294 360792 231676
rect 360752 229288 360804 229294
rect 360752 229230 360804 229236
rect 360936 229288 360988 229294
rect 360936 229230 360988 229236
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359556 221740 359608 221746
rect 359556 221682 359608 221688
rect 359372 218068 359424 218074
rect 359372 218010 359424 218016
rect 359568 217274 359596 221682
rect 360384 220244 360436 220250
rect 360384 220186 360436 220192
rect 360396 217274 360424 220186
rect 360948 219434 360976 229230
rect 361408 227458 361436 231676
rect 361868 231662 362066 231690
rect 362328 231662 362710 231690
rect 361868 229094 361896 231662
rect 361868 229066 361988 229094
rect 361396 227452 361448 227458
rect 361396 227394 361448 227400
rect 361212 227316 361264 227322
rect 361212 227258 361264 227264
rect 361764 227316 361816 227322
rect 361764 227258 361816 227264
rect 360856 219406 360976 219434
rect 360856 218754 360884 219406
rect 360844 218748 360896 218754
rect 360844 218690 360896 218696
rect 361224 217274 361252 227258
rect 361776 226914 361804 227258
rect 361764 226908 361816 226914
rect 361764 226850 361816 226856
rect 361960 221610 361988 229066
rect 361948 221604 362000 221610
rect 361948 221546 362000 221552
rect 362040 221468 362092 221474
rect 362040 221410 362092 221416
rect 362052 217274 362080 221410
rect 362328 221338 362356 231662
rect 363340 229294 363368 231676
rect 363328 229288 363380 229294
rect 363328 229230 363380 229236
rect 362868 228404 362920 228410
rect 362868 228346 362920 228352
rect 362316 221332 362368 221338
rect 362316 221274 362368 221280
rect 362880 217274 362908 228346
rect 363984 223310 364012 231676
rect 364156 229900 364208 229906
rect 364156 229842 364208 229848
rect 363972 223304 364024 223310
rect 363972 223246 364024 223252
rect 364168 218074 364196 229842
rect 364628 224670 364656 231676
rect 364812 231662 365286 231690
rect 364616 224664 364668 224670
rect 364616 224606 364668 224612
rect 364812 224262 364840 231662
rect 365916 225894 365944 231676
rect 366560 228818 366588 231676
rect 366548 228812 366600 228818
rect 366548 228754 366600 228760
rect 366916 228540 366968 228546
rect 366916 228482 366968 228488
rect 366364 227792 366416 227798
rect 366364 227734 366416 227740
rect 365904 225888 365956 225894
rect 365904 225830 365956 225836
rect 364800 224256 364852 224262
rect 364800 224198 364852 224204
rect 364984 224256 365036 224262
rect 364984 224198 365036 224204
rect 364996 219162 365024 224198
rect 366376 219434 366404 227734
rect 366364 219428 366416 219434
rect 366364 219370 366416 219376
rect 364984 219156 365036 219162
rect 364984 219098 365036 219104
rect 366732 218884 366784 218890
rect 366732 218826 366784 218832
rect 365352 218340 365404 218346
rect 365352 218282 365404 218288
rect 364524 218204 364576 218210
rect 364524 218146 364576 218152
rect 363696 218068 363748 218074
rect 363696 218010 363748 218016
rect 364156 218068 364208 218074
rect 364156 218010 364208 218016
rect 357866 217110 357940 217138
rect 358694 217110 358768 217138
rect 359522 217246 359596 217274
rect 360350 217246 360424 217274
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362834 217246 362908 217274
rect 357866 216988 357894 217110
rect 358694 216988 358722 217110
rect 359522 216988 359550 217246
rect 360350 216988 360378 217246
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363708 217138 363736 218010
rect 364536 217138 364564 218146
rect 365364 217138 365392 218282
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366192 217138 366220 218010
rect 366744 217274 366772 218826
rect 366928 218074 366956 228482
rect 367204 226030 367232 231676
rect 367388 231662 367862 231690
rect 367192 226024 367244 226030
rect 367192 225966 367244 225972
rect 367388 220114 367416 231662
rect 367652 225888 367704 225894
rect 367652 225830 367704 225836
rect 367376 220108 367428 220114
rect 367376 220050 367428 220056
rect 367664 218210 367692 225830
rect 368492 222902 368520 231676
rect 369136 228954 369164 231676
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 369780 228682 369808 231676
rect 369768 228676 369820 228682
rect 369768 228618 369820 228624
rect 369124 227928 369176 227934
rect 369124 227870 369176 227876
rect 368480 222896 368532 222902
rect 368480 222838 368532 222844
rect 367836 220108 367888 220114
rect 367836 220050 367888 220056
rect 367652 218204 367704 218210
rect 367652 218146 367704 218152
rect 366916 218068 366968 218074
rect 366916 218010 366968 218016
rect 367848 217274 367876 220050
rect 369136 219026 369164 227870
rect 369768 227044 369820 227050
rect 369768 226986 369820 226992
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 369492 218204 369544 218210
rect 369492 218146 369544 218152
rect 368664 218068 368716 218074
rect 368664 218010 368716 218016
rect 366744 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367802 217246 367876 217274
rect 367802 216988 367830 217246
rect 368676 217138 368704 218010
rect 369504 217138 369532 218146
rect 369780 218074 369808 226986
rect 370424 225622 370452 231676
rect 371068 229770 371096 231676
rect 371436 231662 371726 231690
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 370964 229628 371016 229634
rect 370964 229570 371016 229576
rect 370412 225616 370464 225622
rect 370412 225558 370464 225564
rect 370504 223032 370556 223038
rect 370504 222974 370556 222980
rect 370516 218210 370544 222974
rect 370504 218204 370556 218210
rect 370504 218146 370556 218152
rect 370976 218074 371004 229570
rect 371148 220516 371200 220522
rect 371148 220458 371200 220464
rect 369768 218068 369820 218074
rect 369768 218010 369820 218016
rect 370320 218068 370372 218074
rect 370320 218010 370372 218016
rect 370964 218068 371016 218074
rect 370964 218010 371016 218016
rect 370332 217138 370360 218010
rect 371160 217274 371188 220458
rect 371436 220386 371464 231662
rect 372356 227322 372384 231676
rect 373000 227798 373028 231676
rect 372988 227792 373040 227798
rect 372988 227734 373040 227740
rect 372344 227316 372396 227322
rect 372344 227258 372396 227264
rect 373264 227316 373316 227322
rect 373264 227258 373316 227264
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371424 220380 371476 220386
rect 371424 220322 371476 220328
rect 372540 218074 372568 225558
rect 373276 218346 373304 227258
rect 373644 227186 373672 231676
rect 373816 228676 373868 228682
rect 373816 228618 373868 228624
rect 373632 227180 373684 227186
rect 373632 227122 373684 227128
rect 373632 219020 373684 219026
rect 373632 218962 373684 218968
rect 373264 218340 373316 218346
rect 373264 218282 373316 218288
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 368630 217110 368704 217138
rect 369458 217110 369532 217138
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 368630 216988 368658 217110
rect 369458 216988 369486 217110
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217138 373672 218962
rect 373828 218074 373856 228618
rect 374288 224398 374316 231676
rect 374932 227594 374960 231676
rect 375576 227934 375604 231676
rect 375564 227928 375616 227934
rect 375564 227870 375616 227876
rect 374920 227588 374972 227594
rect 374920 227530 374972 227536
rect 374276 224392 374328 224398
rect 374276 224334 374328 224340
rect 375288 224392 375340 224398
rect 375288 224334 375340 224340
rect 375104 222896 375156 222902
rect 375104 222838 375156 222844
rect 375116 219434 375144 222838
rect 375300 219434 375328 224334
rect 376220 223174 376248 231676
rect 376576 228812 376628 228818
rect 376576 228754 376628 228760
rect 376208 223168 376260 223174
rect 376208 223110 376260 223116
rect 374460 219428 374512 219434
rect 375116 219406 375236 219434
rect 375300 219428 375432 219434
rect 375300 219406 375380 219428
rect 374460 219370 374512 219376
rect 373816 218068 373868 218074
rect 373816 218010 373868 218016
rect 374472 217138 374500 219370
rect 375208 217274 375236 219406
rect 375380 219370 375432 219376
rect 376588 218074 376616 228754
rect 376864 221746 376892 231676
rect 377232 231662 377522 231690
rect 377232 227458 377260 231662
rect 377404 230444 377456 230450
rect 377404 230386 377456 230392
rect 377220 227452 377272 227458
rect 377220 227394 377272 227400
rect 376852 221740 376904 221746
rect 376852 221682 376904 221688
rect 377416 220250 377444 230386
rect 378152 224262 378180 231676
rect 378796 230450 378824 231676
rect 378784 230444 378836 230450
rect 378784 230386 378836 230392
rect 378968 229152 379020 229158
rect 378968 229094 379020 229100
rect 378140 224256 378192 224262
rect 378140 224198 378192 224204
rect 377772 221604 377824 221610
rect 377772 221546 377824 221552
rect 377404 220244 377456 220250
rect 377404 220186 377456 220192
rect 376944 218204 376996 218210
rect 376944 218146 376996 218152
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376576 218068 376628 218074
rect 376576 218010 376628 218016
rect 375208 217246 375282 217274
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217110 373672 217138
rect 374426 217110 374500 217138
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217110
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218146
rect 377784 217274 377812 221546
rect 378980 219434 379008 229094
rect 379440 228410 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 379624 225894 379652 231662
rect 380268 229094 380296 231662
rect 380440 230036 380492 230042
rect 380440 229978 380492 229984
rect 380452 229094 380480 229978
rect 381372 229906 381400 231676
rect 381360 229900 381412 229906
rect 381360 229842 381412 229848
rect 379900 229066 380296 229094
rect 380360 229066 380480 229094
rect 379612 225888 379664 225894
rect 379612 225830 379664 225836
rect 379336 225752 379388 225758
rect 379336 225694 379388 225700
rect 378796 219406 379008 219434
rect 378796 218890 378824 219406
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379152 218748 379204 218754
rect 379152 218690 379204 218696
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379164 217274 379192 218690
rect 379348 218074 379376 225694
rect 379900 221474 379928 229066
rect 380360 224210 380388 229066
rect 382016 228546 382044 231676
rect 382476 231662 382674 231690
rect 382004 228540 382056 228546
rect 382004 228482 382056 228488
rect 381728 228404 381780 228410
rect 381728 228346 381780 228352
rect 380084 224182 380388 224210
rect 379888 221468 379940 221474
rect 379888 221410 379940 221416
rect 380084 219026 380112 224182
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 379336 218068 379388 218074
rect 379336 218010 379388 218016
rect 379164 217246 379422 217274
rect 378566 217110 378640 217138
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381740 218074 381768 228346
rect 381912 227180 381964 227186
rect 381912 227122 381964 227128
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381728 218068 381780 218074
rect 381728 218010 381780 218016
rect 381096 217138 381124 218010
rect 381924 217274 381952 227122
rect 382476 220114 382504 231662
rect 383304 227458 383332 231676
rect 383948 229158 383976 231676
rect 384304 229900 384356 229906
rect 384304 229842 384356 229848
rect 383936 229152 383988 229158
rect 383936 229094 383988 229100
rect 383292 227452 383344 227458
rect 383292 227394 383344 227400
rect 382924 227316 382976 227322
rect 382924 227258 382976 227264
rect 382464 220108 382516 220114
rect 382464 220050 382516 220056
rect 382740 220108 382792 220114
rect 382740 220050 382792 220056
rect 382752 217274 382780 220050
rect 382936 218210 382964 227258
rect 384316 219434 384344 229842
rect 384592 223038 384620 231676
rect 384580 223032 384632 223038
rect 384580 222974 384632 222980
rect 385236 220522 385264 231676
rect 385880 227050 385908 231676
rect 386524 229770 386552 231676
rect 386512 229764 386564 229770
rect 386512 229706 386564 229712
rect 386972 229764 387024 229770
rect 386972 229706 387024 229712
rect 386984 229094 387012 229706
rect 387168 229094 387196 231676
rect 386984 229066 387104 229094
rect 387168 229066 387288 229094
rect 385868 227044 385920 227050
rect 385868 226986 385920 226992
rect 386328 227044 386380 227050
rect 386328 226986 386380 226992
rect 385224 220516 385276 220522
rect 385224 220458 385276 220464
rect 384304 219428 384356 219434
rect 384304 219370 384356 219376
rect 383568 219292 383620 219298
rect 383568 219234 383620 219240
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217246 381952 217274
rect 382706 217246 382780 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217246
rect 382706 216988 382734 217246
rect 383580 217138 383608 219234
rect 384396 219020 384448 219026
rect 384396 218962 384448 218968
rect 384408 217138 384436 218962
rect 386052 218884 386104 218890
rect 386052 218826 386104 218832
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 385236 217138 385264 218010
rect 386064 217138 386092 218826
rect 386340 218074 386368 226986
rect 387076 219298 387104 229066
rect 387260 228682 387288 229066
rect 387248 228676 387300 228682
rect 387248 228618 387300 228624
rect 387812 224398 387840 231676
rect 388088 231662 388470 231690
rect 388088 225622 388116 231662
rect 389100 230042 389128 231676
rect 389088 230036 389140 230042
rect 389088 229978 389140 229984
rect 389744 228818 389772 231676
rect 390020 231662 390402 231690
rect 389732 228812 389784 228818
rect 389732 228754 389784 228760
rect 388076 225616 388128 225622
rect 388076 225558 388128 225564
rect 388444 225616 388496 225622
rect 388444 225558 388496 225564
rect 387800 224392 387852 224398
rect 387800 224334 387852 224340
rect 387708 223032 387760 223038
rect 387708 222974 387760 222980
rect 387064 219292 387116 219298
rect 387064 219234 387116 219240
rect 386880 218204 386932 218210
rect 386880 218146 386932 218152
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 386892 217138 386920 218146
rect 387720 217274 387748 222974
rect 388456 218210 388484 225558
rect 389088 224256 389140 224262
rect 389088 224198 389140 224204
rect 388444 218204 388496 218210
rect 388444 218146 388496 218152
rect 389100 218074 389128 224198
rect 390020 221610 390048 231662
rect 390284 228676 390336 228682
rect 390284 228618 390336 228624
rect 390008 221604 390060 221610
rect 390008 221546 390060 221552
rect 390100 220244 390152 220250
rect 390100 220186 390152 220192
rect 388536 218068 388588 218074
rect 388536 218010 388588 218016
rect 389088 218068 389140 218074
rect 389088 218010 389140 218016
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 383534 217110 383608 217138
rect 384362 217110 384436 217138
rect 385190 217110 385264 217138
rect 386018 217110 386092 217138
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 383534 216988 383562 217110
rect 384362 216988 384390 217110
rect 385190 216988 385218 217110
rect 386018 216988 386046 217110
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388548 217138 388576 218010
rect 389376 217138 389404 218010
rect 390112 217274 390140 220186
rect 390296 218074 390324 228618
rect 391032 222902 391060 231676
rect 391676 227322 391704 231676
rect 392136 231662 392334 231690
rect 391848 228404 391900 228410
rect 391848 228346 391900 228352
rect 391664 227316 391716 227322
rect 391664 227258 391716 227264
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221468 391072 221474
rect 391020 221410 391072 221416
rect 390284 218068 390336 218074
rect 390284 218010 390336 218016
rect 391032 217274 391060 221410
rect 391860 217274 391888 228346
rect 392136 218754 392164 231662
rect 392964 228546 392992 231676
rect 392952 228540 393004 228546
rect 392952 228482 393004 228488
rect 393228 228540 393280 228546
rect 393228 228482 393280 228488
rect 392124 218748 392176 218754
rect 392124 218690 392176 218696
rect 393240 218074 393268 228482
rect 393608 225758 393636 231676
rect 394252 229906 394280 231676
rect 394804 231662 394910 231690
rect 394240 229900 394292 229906
rect 394240 229842 394292 229848
rect 393964 227792 394016 227798
rect 393964 227734 394016 227740
rect 393596 225752 393648 225758
rect 393596 225694 393648 225700
rect 393976 219026 394004 227734
rect 394608 225752 394660 225758
rect 394608 225694 394660 225700
rect 393964 219020 394016 219026
rect 393964 218962 394016 218968
rect 394332 218204 394384 218210
rect 394332 218146 394384 218152
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393228 218068 393280 218074
rect 393228 218010 393280 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 390112 217246 390186 217274
rect 388502 217110 388576 217138
rect 389330 217110 389404 217138
rect 388502 216988 388530 217110
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 217246 391060 217274
rect 391814 217246 391888 217274
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217138 394372 218146
rect 394620 218074 394648 225694
rect 394804 220114 394832 231662
rect 395540 227798 395568 231676
rect 395528 227792 395580 227798
rect 395528 227734 395580 227740
rect 395988 227316 396040 227322
rect 395988 227258 396040 227264
rect 394792 220108 394844 220114
rect 394792 220050 394844 220056
rect 395804 218748 395856 218754
rect 395804 218690 395856 218696
rect 394608 218068 394660 218074
rect 394608 218010 394660 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395172 217138 395200 218010
rect 395816 217274 395844 218690
rect 396000 218074 396028 227258
rect 396184 227186 396212 231676
rect 396828 229770 396856 231676
rect 396816 229764 396868 229770
rect 396816 229706 396868 229712
rect 397472 227798 397500 231676
rect 396632 227792 396684 227798
rect 396632 227734 396684 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396172 227180 396224 227186
rect 396172 227122 396224 227128
rect 396644 218890 396672 227734
rect 398116 223038 398144 231676
rect 398760 227050 398788 231676
rect 398748 227044 398800 227050
rect 398748 226986 398800 226992
rect 398472 226908 398524 226914
rect 398472 226850 398524 226856
rect 398104 223032 398156 223038
rect 398104 222974 398156 222980
rect 397368 222896 397420 222902
rect 397368 222838 397420 222844
rect 396632 218884 396684 218890
rect 396632 218826 396684 218832
rect 397380 218074 397408 222838
rect 397644 220108 397696 220114
rect 397644 220050 397696 220056
rect 395988 218068 396040 218074
rect 395988 218010 396040 218016
rect 396816 218068 396868 218074
rect 396816 218010 396868 218016
rect 397368 218068 397420 218074
rect 397368 218010 397420 218016
rect 395816 217246 395982 217274
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217110 394372 217138
rect 395126 217110 395200 217138
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217110
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396828 217138 396856 218010
rect 397656 217274 397684 220050
rect 398484 217274 398512 226850
rect 399404 225622 399432 231676
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399392 225616 399444 225622
rect 399392 225558 399444 225564
rect 399864 219434 399892 229706
rect 400048 228682 400076 231676
rect 400232 231662 400706 231690
rect 400968 231662 401350 231690
rect 401704 231662 401994 231690
rect 400232 229094 400260 231662
rect 400232 229066 400352 229094
rect 400036 228676 400088 228682
rect 400036 228618 400088 228624
rect 400128 228540 400180 228546
rect 400128 228482 400180 228488
rect 400140 219434 400168 228482
rect 400324 221474 400352 229066
rect 400968 224262 400996 231662
rect 401416 228812 401468 228818
rect 401416 228754 401468 228760
rect 400956 224256 401008 224262
rect 400956 224198 401008 224204
rect 400312 221468 400364 221474
rect 400312 221410 400364 221416
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 396782 217110 396856 217138
rect 397610 217246 397684 217274
rect 398438 217246 398512 217274
rect 396782 216988 396810 217110
rect 397610 216988 397638 217246
rect 398438 216988 398466 217246
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 401428 218074 401456 228754
rect 401704 220250 401732 231662
rect 402624 228410 402652 231676
rect 402612 228404 402664 228410
rect 402612 228346 402664 228352
rect 403268 227798 403296 231676
rect 403912 228274 403940 231676
rect 404268 230376 404320 230382
rect 404268 230318 404320 230324
rect 403900 228268 403952 228274
rect 403900 228210 403952 228216
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 404084 227792 404136 227798
rect 404084 227734 404136 227740
rect 401692 220244 401744 220250
rect 401692 220186 401744 220192
rect 401784 219020 401836 219026
rect 401784 218962 401836 218968
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 401416 218068 401468 218074
rect 401416 218010 401468 218016
rect 400048 217246 400122 217274
rect 399266 217110 399340 217138
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218962
rect 402256 218210 402284 227734
rect 404096 219434 404124 227734
rect 404280 219434 404308 230318
rect 404556 225758 404584 231676
rect 404740 231662 405214 231690
rect 404544 225752 404596 225758
rect 404544 225694 404596 225700
rect 404740 219434 404768 231662
rect 405096 221468 405148 221474
rect 405096 221410 405148 221416
rect 403440 219428 403492 219434
rect 404096 219406 404216 219434
rect 404280 219428 404412 219434
rect 404280 219406 404360 219428
rect 403440 219370 403492 219376
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402624 217138 402652 218826
rect 403452 217138 403480 219370
rect 404188 217274 404216 219406
rect 404360 219370 404412 219376
rect 404556 219406 404768 219434
rect 404556 218754 404584 219406
rect 404544 218748 404596 218754
rect 404544 218690 404596 218696
rect 405108 217274 405136 221410
rect 405844 220114 405872 231676
rect 406488 227322 406516 231676
rect 406476 227316 406528 227322
rect 406476 227258 406528 227264
rect 406752 224936 406804 224942
rect 406752 224878 406804 224884
rect 405832 220108 405884 220114
rect 405832 220050 405884 220056
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405936 217274 405964 219438
rect 406764 217274 406792 224878
rect 407132 222902 407160 231676
rect 407776 228546 407804 231676
rect 408420 228818 408448 231676
rect 408696 231662 409078 231690
rect 408408 228812 408460 228818
rect 408408 228754 408460 228760
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 407764 227928 407816 227934
rect 407764 227870 407816 227876
rect 407120 222896 407172 222902
rect 407120 222838 407172 222844
rect 407776 219026 407804 227870
rect 408696 226914 408724 231662
rect 408868 230240 408920 230246
rect 408868 230182 408920 230188
rect 408880 227798 408908 230182
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228404 409840 228410
rect 409788 228346 409840 228352
rect 408868 227792 408920 227798
rect 408868 227734 408920 227740
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 408684 226908 408736 226914
rect 408684 226850 408736 226856
rect 408408 222896 408460 222902
rect 408408 222838 408460 222844
rect 407764 219020 407816 219026
rect 407764 218962 407816 218968
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405062 217246 405136 217274
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217246
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 222838
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228346
rect 410352 227798 410380 231676
rect 410996 230246 411024 231676
rect 410984 230240 411036 230246
rect 410984 230182 411036 230188
rect 410892 230036 410944 230042
rect 410892 229978 410944 229984
rect 410904 229094 410932 229978
rect 410720 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410720 218074 410748 229066
rect 410892 228676 410944 228682
rect 410892 228618 410944 228624
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 228618
rect 411640 227934 411668 231676
rect 412284 230382 412312 231676
rect 412744 231662 412942 231690
rect 412272 230376 412324 230382
rect 412272 230318 412324 230324
rect 412456 229764 412508 229770
rect 412456 229706 412508 229712
rect 411628 227928 411680 227934
rect 411628 227870 411680 227876
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412468 218890 412496 229706
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229084 413888 229090
rect 413836 229026 413888 229032
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412456 218884 412508 218890
rect 412456 218826 412508 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229026
rect 414216 221474 414244 231676
rect 414860 224942 414888 231676
rect 415504 228410 415532 231676
rect 416148 228682 416176 231676
rect 416792 229094 416820 231676
rect 417436 230042 417464 231676
rect 417712 231662 418094 231690
rect 418264 231662 418738 231690
rect 417424 230036 417476 230042
rect 417424 229978 417476 229984
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416136 228676 416188 228682
rect 416136 228618 416188 228624
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416688 227792 416740 227798
rect 416688 227734 416740 227740
rect 414848 224936 414900 224942
rect 414848 224878 414900 224884
rect 416504 224256 416556 224262
rect 416504 224198 416556 224204
rect 414204 221468 414256 221474
rect 414204 221410 414256 221416
rect 415032 221060 415084 221066
rect 415032 221002 415084 221008
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 221002
rect 416516 219434 416544 224198
rect 416700 219434 416728 227734
rect 416884 222902 416912 229066
rect 417160 229066 417740 229094
rect 416872 222896 416924 222902
rect 416872 222838 416924 222844
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418264 220794 418292 231662
rect 419368 229770 419396 231676
rect 419356 229764 419408 229770
rect 419356 229706 419408 229712
rect 419448 229288 419500 229294
rect 419448 229230 419500 229236
rect 418252 220788 418304 220794
rect 418252 220730 418304 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 419172 219156 419224 219162
rect 419172 219098 419224 219104
rect 418344 218068 418396 218074
rect 418344 218010 418396 218016
rect 418356 217138 418384 218010
rect 419184 217138 419212 219098
rect 419460 218074 419488 229230
rect 420012 229158 420040 231676
rect 420000 229152 420052 229158
rect 420000 229094 420052 229100
rect 420184 229152 420236 229158
rect 420184 229094 420236 229100
rect 420196 221066 420224 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420184 221060 420236 221066
rect 420184 221002 420236 221008
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 420656 219434 420684 220798
rect 420656 219406 420776 219434
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 423784 231662 423890 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 224262 422248 229066
rect 422208 224256 422260 224262
rect 422208 224198 422260 224204
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423312 224256 423364 224262
rect 423312 224198 423364 224204
rect 422680 219406 422892 219434
rect 422680 219162 422708 219406
rect 422668 219156 422720 219162
rect 422668 219098 422720 219104
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 417482 217110 417556 217138
rect 418310 217110 418384 217138
rect 419138 217110 419212 217138
rect 419966 217110 420040 217138
rect 417482 216988 417510 217110
rect 418310 216988 418338 217110
rect 419138 216988 419166 217110
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 224198
rect 423784 220862 423812 231662
rect 424520 229294 424548 231676
rect 424508 229288 424560 229294
rect 424508 229230 424560 229236
rect 424324 229152 424376 229158
rect 424324 229094 424376 229100
rect 424336 224262 424364 229094
rect 424324 224256 424376 224262
rect 424324 224198 424376 224204
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 423772 220856 423824 220862
rect 423772 220798 423824 220804
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 223650 426480 231676
rect 426820 231662 427110 231690
rect 426440 223644 426492 223650
rect 426440 223586 426492 223592
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427924 231662 428398 231690
rect 428660 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 426992 223644 427044 223650
rect 426992 223586 427044 223592
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 223586
rect 427924 218210 427952 231662
rect 428660 219434 428688 231662
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 429948 219434 429976 231662
rect 430120 220244 430172 220250
rect 430120 220186 430172 220192
rect 428292 219406 428688 219434
rect 429580 219406 429976 219434
rect 427912 218204 427964 218210
rect 427912 218146 427964 218152
rect 428292 218074 428320 219406
rect 429580 218346 429608 219406
rect 429936 218612 429988 218618
rect 429936 218554 429988 218560
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 428280 218068 428332 218074
rect 428280 218010 428332 218016
rect 427464 217138 427492 218010
rect 428476 217274 428504 218146
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217274 429148 218010
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217246 428504 217274
rect 429074 217246 429148 217274
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217246
rect 429074 216988 429102 217246
rect 429948 217138 429976 218554
rect 430132 218210 430160 220186
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 220250 432092 231662
rect 432052 220244 432104 220250
rect 432052 220186 432104 220192
rect 431960 220108 432012 220114
rect 431960 220050 432012 220056
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 430120 218204 430172 218210
rect 430120 218146 430172 218152
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 220050
rect 432708 218618 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218612 432748 218618
rect 432696 218554 432748 218560
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220114 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436692 231690
rect 434812 220108 434864 220114
rect 434812 220050 434864 220056
rect 435284 218210 435312 231662
rect 436100 230308 436152 230314
rect 436100 230250 436152 230256
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218204 435784 218210
rect 435732 218146 435784 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434904 218068 434956 218074
rect 434904 218010 434956 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218010
rect 435744 217138 435772 218146
rect 436112 217258 436140 230250
rect 436284 220380 436336 220386
rect 436284 220322 436336 220328
rect 436296 218074 436324 220322
rect 436664 218210 436692 231662
rect 436756 230330 436784 231676
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436756 230314 436876 230330
rect 436756 230308 436888 230314
rect 436756 230302 436836 230308
rect 436836 230250 436888 230256
rect 437032 220386 437060 231662
rect 437020 220380 437072 220386
rect 437020 220322 437072 220328
rect 436652 218204 436704 218210
rect 436652 218146 436704 218152
rect 437768 218074 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 224954 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 224954 439360 230318
rect 438872 224926 438992 224954
rect 439056 224926 439360 224954
rect 438872 219434 438900 224926
rect 438216 219428 438268 219434
rect 438216 219370 438268 219376
rect 438860 219428 438912 219434
rect 438860 219370 438912 219376
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437756 218068 437808 218074
rect 437756 218010 437808 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 219370
rect 439056 217274 439084 224926
rect 440344 219434 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 219428 439924 219434
rect 439872 219370 439924 219376
rect 440332 219428 440384 219434
rect 440332 219370 440384 219376
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 219370
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 224954 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 224926 441752 224954
rect 441632 218090 441660 224926
rect 441540 218062 441660 218090
rect 441540 217274 441568 218062
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441494 217246 441568 217274
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230246 443868 231676
rect 444484 230450 444512 231676
rect 444668 231662 445142 231690
rect 444472 230444 444524 230450
rect 444472 230386 444524 230392
rect 444668 230330 444696 231662
rect 444484 230302 444696 230330
rect 443828 230240 443880 230246
rect 443828 230182 443880 230188
rect 443472 229066 443960 229094
rect 443932 217274 443960 229066
rect 444484 224954 444512 230302
rect 444656 230240 444708 230246
rect 444656 230182 444708 230188
rect 444668 224954 444696 230182
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 447060 230042 447088 231676
rect 447244 231662 447718 231690
rect 447048 230036 447100 230042
rect 447048 229978 447100 229984
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 445772 229066 446444 229094
rect 444484 224926 444604 224954
rect 444668 224926 445616 224954
rect 444576 217274 444604 224926
rect 445588 217274 445616 224926
rect 446416 217274 446444 229066
rect 447244 219434 447272 231662
rect 447600 230444 447652 230450
rect 447600 230386 447652 230392
rect 447612 219434 447640 230386
rect 448348 230382 448376 231676
rect 448336 230376 448388 230382
rect 448336 230318 448388 230324
rect 448992 229566 449020 231676
rect 449636 230382 449664 231676
rect 449164 230376 449216 230382
rect 449164 230318 449216 230324
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448612 229424 448664 229430
rect 448612 229366 448664 229372
rect 448624 229094 448652 229366
rect 449176 229094 449204 230318
rect 449900 230036 449952 230042
rect 449900 229978 449952 229984
rect 448624 229066 448928 229094
rect 449176 229066 449756 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444576 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441494 216988 441522 217246
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448900 217274 448928 229066
rect 449728 217274 449756 229066
rect 449912 219434 449940 229978
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 230318
rect 450924 229430 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451372 229560 451424 229566
rect 451372 229502 451424 229508
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 450556 229066 450768 229094
rect 449912 219406 450584 219434
rect 450556 217274 450584 219406
rect 450740 219298 450768 229066
rect 451384 224262 451412 229502
rect 451832 229288 451884 229294
rect 451832 229230 451884 229236
rect 451372 224256 451424 224262
rect 451372 224198 451424 224204
rect 451844 219434 451872 229230
rect 452200 224256 452252 224262
rect 452200 224198 452252 224204
rect 451476 219406 451872 219434
rect 450728 219292 450780 219298
rect 450728 219234 450780 219240
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448900 217246 448974 217274
rect 449728 217246 449802 217274
rect 450556 217246 450630 217274
rect 448106 217194 448158 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449774 216988 449802 217246
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 224198
rect 452580 221474 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 453028 229424 453080 229430
rect 453028 229366 453080 229372
rect 452568 221468 452620 221474
rect 452568 221410 452620 221416
rect 453040 217274 453068 229366
rect 453316 218074 453344 230182
rect 453500 230110 453528 231676
rect 454144 230246 454172 231676
rect 454802 231662 455092 231690
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230240 454184 230246
rect 454132 230182 454184 230188
rect 453488 230104 453540 230110
rect 453488 230046 453540 230052
rect 454328 229094 454356 230318
rect 454328 229066 454724 229094
rect 453856 219292 453908 219298
rect 453856 219234 453908 219240
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 219234
rect 454696 217274 454724 229066
rect 455064 218210 455092 231662
rect 455236 230240 455288 230246
rect 455236 230182 455288 230188
rect 455248 220794 455276 230182
rect 455432 229634 455460 231676
rect 455788 230104 455840 230110
rect 455788 230046 455840 230052
rect 455420 229628 455472 229634
rect 455420 229570 455472 229576
rect 455236 220788 455288 220794
rect 455236 220730 455288 220736
rect 455800 219434 455828 230046
rect 456076 224602 456104 231676
rect 456064 224596 456116 224602
rect 456064 224538 456116 224544
rect 456720 221610 456748 231676
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 457168 229628 457220 229634
rect 457168 229570 457220 229576
rect 456708 221604 456760 221610
rect 456708 221546 456760 221552
rect 456708 221468 456760 221474
rect 456708 221410 456760 221416
rect 455800 219406 456380 219434
rect 455052 218204 455104 218210
rect 455052 218146 455104 218152
rect 455512 218068 455564 218074
rect 455512 218010 455564 218016
rect 454696 217246 454770 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455524 217138 455552 218010
rect 456352 217274 456380 219406
rect 456720 218074 456748 221410
rect 457180 219434 457208 229570
rect 458008 223582 458036 231676
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 457996 223576 458048 223582
rect 457996 223518 458048 223524
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 457180 219406 458036 219434
rect 456708 218068 456760 218074
rect 456708 218010 456760 218016
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 456352 217246 456426 217274
rect 455524 217110 455598 217138
rect 455570 216988 455598 217110
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459652 224596 459704 224602
rect 459652 224538 459704 224544
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459664 217274 459692 224538
rect 459940 222902 459968 231676
rect 460584 224738 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224732 460624 224738
rect 460572 224674 460624 224680
rect 460204 223576 460256 223582
rect 460204 223518 460256 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 460216 218754 460244 223518
rect 460204 218748 460256 218754
rect 460204 218690 460256 218696
rect 461308 218748 461360 218754
rect 461308 218690 461360 218696
rect 460480 218204 460532 218210
rect 460480 218146 460532 218152
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 459664 217246 459738 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 216988 459738 217246
rect 460492 217138 460520 218146
rect 461320 217138 461348 218690
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224398 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224392 462556 224398
rect 462504 224334 462556 224340
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 221604 462188 221610
rect 462136 221546 462188 221552
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 221546
rect 462976 217274 463004 225762
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224732 463200 224738
rect 463148 224674 463200 224680
rect 463160 218074 463188 224674
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 230042 467052 231676
rect 467012 230036 467064 230042
rect 467012 229978 467064 229984
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 460492 217110 460566 217138
rect 461320 217110 461394 217138
rect 460538 216988 460566 217110
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 229770 468340 231676
rect 468956 229906 468984 231676
rect 469600 229906 469628 231676
rect 468944 229900 468996 229906
rect 468944 229842 468996 229848
rect 469588 229900 469640 229906
rect 469588 229842 469640 229848
rect 468300 229764 468352 229770
rect 468300 229706 468352 229712
rect 469128 229764 469180 229770
rect 469128 229706 469180 229712
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 469140 220386 469168 229706
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224392 469364 224398
rect 469312 224334 469364 224340
rect 469128 220380 469180 220386
rect 469128 220322 469180 220328
rect 468772 217246 468846 217274
rect 469324 217258 469352 224334
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224398 470272 231676
rect 470888 230246 470916 231676
rect 470876 230240 470928 230246
rect 470876 230182 470928 230188
rect 471532 227934 471560 231676
rect 471888 230240 471940 230246
rect 471888 230182 471940 230188
rect 471520 227928 471572 227934
rect 471520 227870 471572 227876
rect 470232 224392 470284 224398
rect 470232 224334 470284 224340
rect 471900 222154 471928 230182
rect 472176 227050 472204 231676
rect 472834 231662 473032 231690
rect 472164 227044 472216 227050
rect 472164 226986 472216 226992
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471704 220856 471756 220862
rect 471704 220798 471756 220804
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 471716 218074 471744 220798
rect 473004 220250 473032 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474766 231662 475056 231690
rect 474004 230036 474056 230042
rect 474004 229978 474056 229984
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 472992 220244 473044 220250
rect 472992 220186 473044 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471704 218068 471756 218074
rect 471704 218010 471756 218016
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220658 474044 229978
rect 474476 229094 474504 231662
rect 474476 229066 474780 229094
rect 474752 224262 474780 229066
rect 475028 227798 475056 231662
rect 475396 230382 475424 231676
rect 475384 230376 475436 230382
rect 475384 230318 475436 230324
rect 476040 230110 476068 231676
rect 476684 230246 476712 231676
rect 476672 230240 476724 230246
rect 476672 230182 476724 230188
rect 476028 230104 476080 230110
rect 476028 230046 476080 230052
rect 476764 229900 476816 229906
rect 476764 229842 476816 229848
rect 475384 229764 475436 229770
rect 475384 229706 475436 229712
rect 475016 227792 475068 227798
rect 475016 227734 475068 227740
rect 474740 224256 474792 224262
rect 474740 224198 474792 224204
rect 475396 220794 475424 229706
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474004 220652 474056 220658
rect 474004 220594 474056 220600
rect 475384 220652 475436 220658
rect 475384 220594 475436 220600
rect 474556 220380 474608 220386
rect 474556 220322 474608 220328
rect 474568 217274 474596 220322
rect 475396 217274 475424 220594
rect 475580 218346 475608 223518
rect 476212 220788 476264 220794
rect 476212 220730 476264 220736
rect 475568 218340 475620 218346
rect 475568 218282 475620 218288
rect 476224 217274 476252 220730
rect 476592 217274 476620 225558
rect 476776 220794 476804 229842
rect 477328 225622 477356 231676
rect 477986 231662 478552 231690
rect 478630 231662 478828 231690
rect 478328 230376 478380 230382
rect 478328 230318 478380 230324
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 478340 222902 478368 230318
rect 478328 222896 478380 222902
rect 478328 222838 478380 222844
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478524 220114 478552 231662
rect 478800 228682 478828 231662
rect 479260 229906 479288 231676
rect 479708 230240 479760 230246
rect 479708 230182 479760 230188
rect 479524 230104 479576 230110
rect 479524 230046 479576 230052
rect 479248 229900 479300 229906
rect 479248 229842 479300 229848
rect 478788 228676 478840 228682
rect 478788 228618 478840 228624
rect 479340 227928 479392 227934
rect 479340 227870 479392 227876
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478512 220108 478564 220114
rect 478512 220050 478564 220056
rect 478708 217274 478736 220730
rect 479352 219434 479380 227870
rect 479536 224534 479564 230046
rect 479720 228274 479748 230182
rect 479904 229294 479932 231676
rect 480548 230382 480576 231676
rect 480536 230376 480588 230382
rect 480536 230318 480588 230324
rect 479892 229288 479944 229294
rect 479892 229230 479944 229236
rect 479708 228268 479760 228274
rect 479708 228210 479760 228216
rect 481192 227186 481220 231676
rect 481548 230376 481600 230382
rect 481548 230318 481600 230324
rect 481180 227180 481232 227186
rect 481180 227122 481232 227128
rect 481180 227044 481232 227050
rect 481180 226986 481232 226992
rect 479524 224528 479576 224534
rect 479524 224470 479576 224476
rect 479708 224392 479760 224398
rect 479708 224334 479760 224340
rect 479352 219406 479564 219434
rect 479536 217274 479564 219406
rect 479720 219298 479748 224334
rect 479708 219292 479760 219298
rect 479708 219234 479760 219240
rect 480352 219292 480404 219298
rect 480352 219234 480404 219240
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480364 217138 480392 219234
rect 481192 217274 481220 226986
rect 481560 220386 481588 230318
rect 481836 229770 481864 231676
rect 481824 229764 481876 229770
rect 481824 229706 481876 229712
rect 482284 229288 482336 229294
rect 482284 229230 482336 229236
rect 482296 220522 482324 229230
rect 482480 228546 482508 231676
rect 483124 230042 483152 231676
rect 483112 230036 483164 230042
rect 483112 229978 483164 229984
rect 483768 229294 483796 231676
rect 484426 231662 484808 231690
rect 484780 230042 484808 231662
rect 484308 230036 484360 230042
rect 484308 229978 484360 229984
rect 484768 230036 484820 230042
rect 484768 229978 484820 229984
rect 484032 229900 484084 229906
rect 484032 229842 484084 229848
rect 483756 229288 483808 229294
rect 483756 229230 483808 229236
rect 483572 228676 483624 228682
rect 483572 228618 483624 228624
rect 482468 228540 482520 228546
rect 482468 228482 482520 228488
rect 482928 227792 482980 227798
rect 482928 227734 482980 227740
rect 482940 222222 482968 227734
rect 482928 222216 482980 222222
rect 482928 222158 482980 222164
rect 482284 220516 482336 220522
rect 482284 220458 482336 220464
rect 481548 220380 481600 220386
rect 481548 220322 481600 220328
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482940 218482 482968 222158
rect 483584 219162 483612 228618
rect 484044 228138 484072 229842
rect 484032 228132 484084 228138
rect 484032 228074 484084 228080
rect 484320 221746 484348 229978
rect 485056 227322 485084 231676
rect 485044 227316 485096 227322
rect 485044 227258 485096 227264
rect 485700 224262 485728 231676
rect 486344 229906 486372 231676
rect 486332 229900 486384 229906
rect 486332 229842 486384 229848
rect 486792 229288 486844 229294
rect 486792 229230 486844 229236
rect 486608 224528 486660 224534
rect 486608 224470 486660 224476
rect 484584 224256 484636 224262
rect 484584 224198 484636 224204
rect 485688 224256 485740 224262
rect 485688 224198 485740 224204
rect 484308 221740 484360 221746
rect 484308 221682 484360 221688
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 483572 219156 483624 219162
rect 483572 219098 483624 219104
rect 482928 218476 482980 218482
rect 482928 218418 482980 218424
rect 482836 218340 482888 218346
rect 482836 218282 482888 218288
rect 482848 217274 482876 218282
rect 483768 217274 483796 221410
rect 484596 219473 484624 224198
rect 486148 222896 486200 222902
rect 486148 222838 486200 222844
rect 484582 219464 484638 219473
rect 484582 219399 484638 219408
rect 484596 217274 484624 219399
rect 485320 218476 485372 218482
rect 485320 218418 485372 218424
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 482848 217246 482922 217274
rect 480364 217110 480438 217138
rect 480410 216988 480438 217110
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482894 216988 482922 217246
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485332 217138 485360 218418
rect 486160 217138 486188 222838
rect 486620 220969 486648 224470
rect 486804 224398 486832 229230
rect 486792 224392 486844 224398
rect 486792 224334 486844 224340
rect 486988 222902 487016 231676
rect 487632 228410 487660 231676
rect 488290 231662 488488 231690
rect 487620 228404 487672 228410
rect 487620 228346 487672 228352
rect 487804 228268 487856 228274
rect 487804 228210 487856 228216
rect 486976 222896 487028 222902
rect 486976 222838 487028 222844
rect 486606 220960 486662 220969
rect 486606 220895 486662 220904
rect 486620 217274 486648 220895
rect 487816 218113 487844 228210
rect 488460 220250 488488 231662
rect 488920 225894 488948 231676
rect 488908 225888 488960 225894
rect 488908 225830 488960 225836
rect 489184 225616 489236 225622
rect 489184 225558 489236 225564
rect 488448 220244 488500 220250
rect 488448 220186 488500 220192
rect 489196 219434 489224 225558
rect 489564 223310 489592 231676
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 489932 225010 489960 229706
rect 489920 225004 489972 225010
rect 489920 224946 489972 224952
rect 489552 223304 489604 223310
rect 489552 223246 489604 223252
rect 490208 223174 490236 231676
rect 490852 230110 490880 231676
rect 490840 230104 490892 230110
rect 490840 230046 490892 230052
rect 490656 230036 490708 230042
rect 490656 229978 490708 229984
rect 490668 229634 490696 229978
rect 490656 229628 490708 229634
rect 490656 229570 490708 229576
rect 490564 228132 490616 228138
rect 490564 228074 490616 228080
rect 490196 223168 490248 223174
rect 490196 223110 490248 223116
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 488724 219428 488776 219434
rect 488724 219370 488776 219376
rect 489184 219428 489236 219434
rect 489184 219370 489236 219376
rect 487802 218104 487858 218113
rect 488736 218074 488764 219370
rect 487802 218039 487858 218048
rect 488724 218068 488776 218074
rect 487816 217274 487844 218039
rect 488724 218010 488776 218016
rect 486620 217246 487062 217274
rect 487816 217246 487890 217274
rect 485332 217110 485406 217138
rect 486160 217110 486234 217138
rect 485378 216988 485406 217110
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488736 217138 488764 218010
rect 489472 217274 489500 220050
rect 490576 219201 490604 228074
rect 491496 225758 491524 231676
rect 492154 231662 492352 231690
rect 491484 225752 491536 225758
rect 491484 225694 491536 225700
rect 491944 220516 491996 220522
rect 491944 220458 491996 220464
rect 490562 219192 490618 219201
rect 490288 219156 490340 219162
rect 490562 219127 490618 219136
rect 491114 219192 491170 219201
rect 491114 219127 491170 219136
rect 490288 219098 490340 219104
rect 490300 218929 490328 219098
rect 490286 218920 490342 218929
rect 490286 218855 490342 218864
rect 489472 217246 489546 217274
rect 488690 217110 488764 217138
rect 488690 216988 488718 217110
rect 489518 216988 489546 217246
rect 490300 217138 490328 218855
rect 491128 218657 491156 219127
rect 491114 218648 491170 218657
rect 491114 218583 491170 218592
rect 491128 217138 491156 218583
rect 491956 217274 491984 220458
rect 492324 220114 492352 231662
rect 492784 230382 492812 231676
rect 492772 230376 492824 230382
rect 492772 230318 492824 230324
rect 493428 230246 493456 231676
rect 494086 231662 494376 231690
rect 493968 230376 494020 230382
rect 493968 230318 494020 230324
rect 493416 230240 493468 230246
rect 493416 230182 493468 230188
rect 493784 230104 493836 230110
rect 493784 230046 493836 230052
rect 493796 228818 493824 230046
rect 493784 228812 493836 228818
rect 493784 228754 493836 228760
rect 492956 227180 493008 227186
rect 492956 227122 493008 227128
rect 492772 220380 492824 220386
rect 492772 220322 492824 220328
rect 492312 220108 492364 220114
rect 492312 220050 492364 220056
rect 491956 217246 492168 217274
rect 490300 217110 490374 217138
rect 491128 217110 491202 217138
rect 490346 216988 490374 217110
rect 491174 216988 491202 217110
rect 492002 216988 492030 217246
rect 492140 217161 492168 217246
rect 492126 217152 492182 217161
rect 492784 217138 492812 220322
rect 492968 219201 492996 227122
rect 493980 220658 494008 230318
rect 494348 230110 494376 231662
rect 494336 230104 494388 230110
rect 494336 230046 494388 230052
rect 494716 229362 494744 231676
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494704 229356 494756 229362
rect 494704 229298 494756 229304
rect 494612 228540 494664 228546
rect 494612 228482 494664 228488
rect 493968 220652 494020 220658
rect 493968 220594 494020 220600
rect 492954 219192 493010 219201
rect 492954 219127 493010 219136
rect 493598 219192 493654 219201
rect 493598 219127 493654 219136
rect 493612 217297 493640 219127
rect 494624 218210 494652 228482
rect 495176 225622 495204 230182
rect 495360 228682 495388 231676
rect 496004 229770 496032 231676
rect 496188 231662 496662 231690
rect 495992 229764 496044 229770
rect 495992 229706 496044 229712
rect 496188 229094 496216 231662
rect 496360 229356 496412 229362
rect 496360 229298 496412 229304
rect 496372 229094 496400 229298
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 495348 228676 495400 228682
rect 495348 228618 495400 228624
rect 495164 225616 495216 225622
rect 495164 225558 495216 225564
rect 494796 225004 494848 225010
rect 494796 224946 494848 224952
rect 494808 219745 494836 224946
rect 496084 221740 496136 221746
rect 496084 221682 496136 221688
rect 494794 219736 494850 219745
rect 494794 219671 494850 219680
rect 494612 218204 494664 218210
rect 494612 218146 494664 218152
rect 493598 217288 493654 217297
rect 494808 217274 494836 219671
rect 495256 218204 495308 218210
rect 495256 218146 495308 218152
rect 493598 217223 493654 217232
rect 494486 217246 494836 217274
rect 493612 217138 493640 217223
rect 492784 217110 492858 217138
rect 493612 217110 493686 217138
rect 492126 217087 492182 217096
rect 492830 216988 492858 217110
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495268 217138 495296 218146
rect 496096 217138 496124 221682
rect 496280 221610 496308 229066
rect 496268 221604 496320 221610
rect 496268 221546 496320 221552
rect 496464 220386 496492 229066
rect 497292 227050 497320 231676
rect 497936 230314 497964 231676
rect 497924 230308 497976 230314
rect 497924 230250 497976 230256
rect 497464 229628 497516 229634
rect 497464 229570 497516 229576
rect 497280 227044 497332 227050
rect 497280 226986 497332 226992
rect 497476 224954 497504 229570
rect 498580 227186 498608 231676
rect 498752 227316 498804 227322
rect 498752 227258 498804 227264
rect 498568 227180 498620 227186
rect 498568 227122 498620 227128
rect 498764 224954 498792 227258
rect 497476 224926 497780 224954
rect 496912 224392 496964 224398
rect 496912 224334 496964 224340
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 496924 218385 496952 224334
rect 497752 219201 497780 224926
rect 498672 224926 498792 224954
rect 497738 219192 497794 219201
rect 497738 219127 497794 219136
rect 496910 218376 496966 218385
rect 496910 218311 496966 218320
rect 496924 217138 496952 218311
rect 497556 218068 497608 218074
rect 497556 218010 497608 218016
rect 497568 217297 497596 218010
rect 497554 217288 497610 217297
rect 497752 217274 497780 219127
rect 498672 217841 498700 224926
rect 499224 224398 499252 231676
rect 499868 229498 499896 231676
rect 500052 231662 500526 231690
rect 499856 229492 499908 229498
rect 499856 229434 499908 229440
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 499396 224256 499448 224262
rect 499396 224198 499448 224204
rect 498658 217832 498714 217841
rect 498658 217767 498714 217776
rect 498672 217274 498700 217767
rect 497752 217246 497826 217274
rect 497554 217223 497610 217232
rect 495268 217110 495342 217138
rect 496096 217110 496170 217138
rect 496924 217110 496998 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217110
rect 496970 216988 496998 217110
rect 497798 216988 497826 217246
rect 498626 217246 498700 217274
rect 498626 216988 498654 217246
rect 499408 217138 499436 224198
rect 500052 222018 500080 231662
rect 500224 229900 500276 229906
rect 500224 229842 500276 229848
rect 500040 222012 500092 222018
rect 500040 221954 500092 221960
rect 500236 218385 500264 229842
rect 501156 223038 501184 231676
rect 501328 229492 501380 229498
rect 501328 229434 501380 229440
rect 501340 227322 501368 229434
rect 501800 229430 501828 231676
rect 501788 229424 501840 229430
rect 501788 229366 501840 229372
rect 502444 228546 502472 231676
rect 503102 231662 503484 231690
rect 503260 230172 503312 230178
rect 503260 230114 503312 230120
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 501512 228404 501564 228410
rect 501512 228346 501564 228352
rect 501328 227316 501380 227322
rect 501328 227258 501380 227264
rect 501524 224954 501552 228346
rect 503272 226302 503300 230114
rect 503260 226296 503312 226302
rect 503260 226238 503312 226244
rect 503076 225888 503128 225894
rect 503076 225830 503128 225836
rect 501524 224926 501920 224954
rect 501144 223032 501196 223038
rect 501144 222974 501196 222980
rect 501052 222896 501104 222902
rect 501052 222838 501104 222844
rect 501064 218482 501092 222838
rect 501052 218476 501104 218482
rect 501052 218418 501104 218424
rect 500038 218376 500094 218385
rect 500038 218311 500040 218320
rect 500092 218311 500094 218320
rect 500222 218376 500278 218385
rect 500222 218311 500278 218320
rect 500040 218282 500092 218288
rect 500236 217274 500264 218311
rect 500236 217246 500310 217274
rect 499408 217110 499482 217138
rect 499454 216988 499482 217110
rect 500282 216988 500310 217246
rect 501064 217138 501092 218418
rect 501892 217274 501920 224926
rect 502708 220244 502760 220250
rect 502708 220186 502760 220192
rect 502720 219201 502748 220186
rect 502522 219192 502578 219201
rect 502522 219127 502578 219136
rect 502706 219192 502762 219201
rect 503088 219162 503116 225830
rect 503456 221746 503484 231662
rect 503732 230042 503760 231676
rect 504390 231662 504680 231690
rect 504364 230308 504416 230314
rect 504364 230250 504416 230256
rect 503720 230036 503772 230042
rect 503720 229978 503772 229984
rect 504376 229094 504404 230250
rect 504192 229066 504404 229094
rect 503444 221740 503496 221746
rect 503444 221682 503496 221688
rect 504192 220250 504220 229066
rect 504364 223304 504416 223310
rect 504364 223246 504416 223252
rect 504180 220244 504232 220250
rect 504180 220186 504232 220192
rect 502706 219127 502762 219136
rect 503076 219156 503128 219162
rect 502536 218686 502564 219127
rect 502524 218680 502576 218686
rect 502524 218622 502576 218628
rect 501892 217246 501966 217274
rect 501064 217110 501138 217138
rect 501110 216988 501138 217110
rect 501938 216988 501966 217246
rect 502720 217138 502748 219127
rect 503076 219098 503128 219104
rect 503536 219156 503588 219162
rect 503536 219098 503588 219104
rect 503548 217569 503576 219098
rect 503534 217560 503590 217569
rect 503534 217495 503590 217504
rect 503548 217138 503576 217495
rect 504376 217138 504404 223246
rect 504652 222902 504680 231662
rect 505020 229094 505048 231676
rect 505664 229906 505692 231676
rect 505652 229900 505704 229906
rect 505652 229842 505704 229848
rect 505020 229066 505140 229094
rect 505112 223310 505140 229066
rect 506020 228812 506072 228818
rect 506020 228754 506072 228760
rect 505100 223304 505152 223310
rect 505100 223246 505152 223252
rect 505652 223168 505704 223174
rect 505652 223110 505704 223116
rect 504640 222896 504692 222902
rect 504640 222838 504692 222844
rect 504640 219360 504692 219366
rect 504640 219302 504692 219308
rect 505284 219360 505336 219366
rect 505284 219302 505336 219308
rect 504652 218385 504680 219302
rect 505296 219201 505324 219302
rect 505098 219192 505154 219201
rect 505098 219127 505154 219136
rect 505282 219192 505338 219201
rect 505282 219127 505338 219136
rect 505112 218770 505140 219127
rect 505112 218742 505324 218770
rect 505008 218680 505060 218686
rect 504822 218648 504878 218657
rect 504822 218583 504878 218592
rect 505006 218648 505008 218657
rect 505060 218648 505062 218657
rect 505006 218583 505062 218592
rect 504638 218376 504694 218385
rect 504638 218311 504694 218320
rect 504836 217841 504864 218583
rect 505296 218385 505324 218742
rect 505282 218376 505338 218385
rect 505282 218311 505338 218320
rect 505664 218074 505692 223110
rect 505836 218884 505888 218890
rect 505836 218826 505888 218832
rect 505284 218068 505336 218074
rect 505284 218010 505336 218016
rect 505652 218068 505704 218074
rect 505652 218010 505704 218016
rect 504822 217832 504878 217841
rect 504822 217767 504878 217776
rect 505296 217138 505324 218010
rect 505848 217841 505876 218826
rect 506032 217841 506060 228754
rect 506308 228410 506336 231676
rect 506966 231662 507348 231690
rect 506940 230036 506992 230042
rect 506940 229978 506992 229984
rect 506952 228834 506980 229978
rect 507124 229424 507176 229430
rect 507124 229366 507176 229372
rect 507136 228954 507164 229366
rect 507124 228948 507176 228954
rect 507124 228890 507176 228896
rect 506952 228806 507072 228834
rect 506296 228404 506348 228410
rect 506296 228346 506348 228352
rect 506848 225752 506900 225758
rect 506848 225694 506900 225700
rect 505834 217832 505890 217841
rect 505834 217767 505890 217776
rect 506018 217832 506074 217841
rect 506018 217767 506074 217776
rect 506032 217274 506060 217767
rect 506860 217274 506888 225694
rect 507044 220522 507072 228806
rect 507320 225758 507348 231662
rect 507596 229158 507624 231676
rect 507584 229152 507636 229158
rect 507584 229094 507636 229100
rect 507308 225752 507360 225758
rect 507308 225694 507360 225700
rect 508240 224534 508268 231676
rect 508228 224528 508280 224534
rect 508228 224470 508280 224476
rect 508884 224262 508912 231676
rect 509528 230042 509556 231676
rect 509516 230036 509568 230042
rect 509516 229978 509568 229984
rect 509240 229764 509292 229770
rect 509240 229706 509292 229712
rect 509252 225010 509280 229706
rect 510172 229094 510200 231676
rect 510172 229066 510384 229094
rect 510160 226296 510212 226302
rect 510160 226238 510212 226244
rect 509700 225616 509752 225622
rect 509700 225558 509752 225564
rect 509240 225004 509292 225010
rect 509712 224954 509740 225558
rect 509240 224946 509292 224952
rect 509436 224926 509740 224954
rect 510172 224954 510200 226238
rect 510356 225622 510384 229066
rect 510816 226166 510844 231676
rect 511460 230246 511488 231676
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 511264 229152 511316 229158
rect 511264 229094 511316 229100
rect 510804 226160 510856 226166
rect 510804 226102 510856 226108
rect 510344 225616 510396 225622
rect 510344 225558 510396 225564
rect 510172 224926 510384 224954
rect 508872 224256 508924 224262
rect 508872 224198 508924 224204
rect 508504 220652 508556 220658
rect 508504 220594 508556 220600
rect 507032 220516 507084 220522
rect 507032 220458 507084 220464
rect 507676 220108 507728 220114
rect 507676 220050 507728 220056
rect 507124 219156 507176 219162
rect 507124 219098 507176 219104
rect 507136 218346 507164 219098
rect 507688 218346 507716 220050
rect 507124 218340 507176 218346
rect 507124 218282 507176 218288
rect 507676 218340 507728 218346
rect 507676 218282 507728 218288
rect 506032 217246 506106 217274
rect 506860 217246 506934 217274
rect 502720 217110 502794 217138
rect 503548 217110 503622 217138
rect 504376 217110 504450 217138
rect 502766 216988 502794 217110
rect 503594 216988 503622 217110
rect 504422 216988 504450 217110
rect 505250 217110 505324 217138
rect 505250 216988 505278 217110
rect 506078 216988 506106 217246
rect 506906 216988 506934 217246
rect 507688 217138 507716 218282
rect 508516 217841 508544 220594
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 508516 217138 508544 217767
rect 509436 217274 509464 224926
rect 510158 218648 510214 218657
rect 509712 218606 510158 218634
rect 509712 218385 509740 218606
rect 510158 218583 510214 218592
rect 510356 218482 510384 224926
rect 511276 220658 511304 229094
rect 512104 228682 512132 231676
rect 512762 231662 513144 231690
rect 511816 228676 511868 228682
rect 511816 228618 511868 228624
rect 512092 228676 512144 228682
rect 512092 228618 512144 228624
rect 511264 220652 511316 220658
rect 511264 220594 511316 220600
rect 510988 220380 511040 220386
rect 510988 220322 511040 220328
rect 511000 220017 511028 220322
rect 510986 220008 511042 220017
rect 510986 219943 511042 219952
rect 510344 218476 510396 218482
rect 510344 218418 510396 218424
rect 509698 218376 509754 218385
rect 509698 218311 509754 218320
rect 510356 217274 510384 218418
rect 509390 217246 509464 217274
rect 510218 217246 510384 217274
rect 507688 217110 507762 217138
rect 508516 217110 508590 217138
rect 507734 216988 507762 217110
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 219943
rect 511828 217274 511856 228618
rect 512644 225004 512696 225010
rect 512644 224946 512696 224952
rect 512656 220017 512684 224946
rect 513116 223174 513144 231662
rect 513392 230382 513420 231676
rect 513380 230376 513432 230382
rect 513380 230318 513432 230324
rect 514036 227050 514064 231676
rect 514024 227044 514076 227050
rect 514024 226986 514076 226992
rect 514300 226908 514352 226914
rect 514300 226850 514352 226856
rect 513104 223168 513156 223174
rect 513104 223110 513156 223116
rect 513378 221640 513434 221649
rect 513378 221575 513380 221584
rect 513432 221575 513434 221584
rect 513380 221546 513432 221552
rect 512642 220008 512698 220017
rect 512642 219943 512698 219952
rect 512656 217274 512684 219943
rect 513392 217274 513420 221546
rect 514312 217274 514340 226850
rect 514680 224670 514708 231676
rect 515338 231662 515720 231690
rect 515404 230376 515456 230382
rect 515404 230318 515456 230324
rect 514668 224664 514720 224670
rect 514668 224606 514720 224612
rect 515416 221882 515444 230318
rect 515692 229770 515720 231662
rect 515876 231662 515982 231690
rect 516626 231662 517192 231690
rect 517270 231662 517468 231690
rect 515680 229764 515732 229770
rect 515680 229706 515732 229712
rect 515876 227594 515904 231662
rect 516508 230240 516560 230246
rect 516508 230182 516560 230188
rect 516048 229900 516100 229906
rect 516048 229842 516100 229848
rect 515864 227588 515916 227594
rect 515864 227530 515916 227536
rect 516060 227186 516088 229842
rect 515864 227180 515916 227186
rect 515864 227122 515916 227128
rect 516048 227180 516100 227186
rect 516048 227122 516100 227128
rect 515876 224954 515904 227122
rect 515784 224926 515904 224954
rect 516520 224942 516548 230182
rect 516508 224936 516560 224942
rect 515404 221876 515456 221882
rect 515404 221818 515456 221824
rect 515784 221241 515812 224926
rect 516508 224878 516560 224884
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 515220 220244 515272 220250
rect 515220 220186 515272 220192
rect 514758 219192 514814 219201
rect 514758 219127 514814 219136
rect 514942 219192 514998 219201
rect 514942 219127 514944 219136
rect 514772 219026 514800 219127
rect 514996 219127 514998 219136
rect 514944 219098 514996 219104
rect 514760 219020 514812 219026
rect 514760 218962 514812 218968
rect 511828 217246 511902 217274
rect 512656 217246 512730 217274
rect 513392 217246 513558 217274
rect 514312 217246 514386 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515232 217138 515260 220186
rect 515784 217274 515812 221167
rect 515956 220244 516008 220250
rect 515956 220186 516008 220192
rect 515968 219570 515996 220186
rect 515956 219564 516008 219570
rect 515956 219506 516008 219512
rect 515784 217246 516042 217274
rect 515186 217110 515260 217138
rect 515186 216988 515214 217110
rect 516014 216988 516042 217246
rect 516796 217138 516824 224334
rect 517164 220386 517192 231662
rect 517440 229906 517468 231662
rect 517428 229900 517480 229906
rect 517428 229842 517480 229848
rect 517900 229090 517928 231676
rect 517888 229084 517940 229090
rect 517888 229026 517940 229032
rect 517704 227316 517756 227322
rect 517704 227258 517756 227264
rect 517716 221785 517744 227258
rect 518544 226030 518572 231676
rect 519188 230042 519216 231676
rect 518900 230036 518952 230042
rect 518900 229978 518952 229984
rect 519176 230036 519228 230042
rect 519176 229978 519228 229984
rect 518532 226024 518584 226030
rect 518532 225966 518584 225972
rect 518912 223446 518940 229978
rect 519832 228818 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 521120 230178 521148 231676
rect 521568 230376 521620 230382
rect 521568 230318 521620 230324
rect 521108 230172 521160 230178
rect 521108 230114 521160 230120
rect 520188 228948 520240 228954
rect 520188 228890 520240 228896
rect 519820 228812 519872 228818
rect 519820 228754 519872 228760
rect 518900 223440 518952 223446
rect 518900 223382 518952 223388
rect 519268 223032 519320 223038
rect 519268 222974 519320 222980
rect 518440 222012 518492 222018
rect 518440 221954 518492 221960
rect 517702 221776 517758 221785
rect 517702 221711 517758 221720
rect 517152 220380 517204 220386
rect 517152 220322 517204 220328
rect 517716 217274 517744 221711
rect 518452 220862 518480 221954
rect 518440 220856 518492 220862
rect 518440 220798 518492 220804
rect 517670 217246 517744 217274
rect 516796 217110 516870 217138
rect 516842 216988 516870 217110
rect 517670 216988 517698 217246
rect 518452 217138 518480 220798
rect 518808 219428 518860 219434
rect 518808 219370 518860 219376
rect 518820 218754 518848 219370
rect 518808 218748 518860 218754
rect 518808 218690 518860 218696
rect 519280 217138 519308 222974
rect 519542 220280 519598 220289
rect 519542 220215 519598 220224
rect 519556 219745 519584 220215
rect 519542 219736 519598 219745
rect 519542 219671 519598 219680
rect 519818 219736 519874 219745
rect 519818 219671 519874 219680
rect 519832 219434 519860 219671
rect 520200 219638 520228 228890
rect 520924 228540 520976 228546
rect 520924 228482 520976 228488
rect 520188 219632 520240 219638
rect 520188 219574 520240 219580
rect 519820 219428 519872 219434
rect 519820 219370 519872 219376
rect 519820 219020 519872 219026
rect 519820 218962 519872 218968
rect 519544 218884 519596 218890
rect 519544 218826 519596 218832
rect 519556 218210 519584 218826
rect 519832 218210 519860 218962
rect 519544 218204 519596 218210
rect 519544 218146 519596 218152
rect 519820 218204 519872 218210
rect 519820 218146 519872 218152
rect 520200 217274 520228 219574
rect 520154 217246 520228 217274
rect 520936 217274 520964 228482
rect 521580 220250 521608 230318
rect 521764 227322 521792 231676
rect 522422 231662 522896 231690
rect 522304 229900 522356 229906
rect 522304 229842 522356 229848
rect 521752 227316 521804 227322
rect 521752 227258 521804 227264
rect 521752 221740 521804 221746
rect 521752 221682 521804 221688
rect 521568 220244 521620 220250
rect 521568 220186 521620 220192
rect 520936 217246 521010 217274
rect 518452 217110 518526 217138
rect 519280 217110 519354 217138
rect 518498 216988 518526 217110
rect 519326 216988 519354 217110
rect 520154 216988 520182 217246
rect 520982 217122 521010 217246
rect 521764 217138 521792 221682
rect 522316 220522 522344 229842
rect 522868 221746 522896 231662
rect 523052 229906 523080 231676
rect 523040 229900 523092 229906
rect 523040 229842 523092 229848
rect 523696 223038 523724 231676
rect 524340 227458 524368 231676
rect 524984 229634 525012 231676
rect 525628 229922 525656 231676
rect 525628 229894 525748 229922
rect 525524 229764 525576 229770
rect 525524 229706 525576 229712
rect 524972 229628 525024 229634
rect 524972 229570 525024 229576
rect 525536 227730 525564 229706
rect 525524 227724 525576 227730
rect 525524 227666 525576 227672
rect 524328 227452 524380 227458
rect 524328 227394 524380 227400
rect 525064 227180 525116 227186
rect 525064 227122 525116 227128
rect 524236 223304 524288 223310
rect 524236 223246 524288 223252
rect 523684 223032 523736 223038
rect 523684 222974 523736 222980
rect 523408 222896 523460 222902
rect 523408 222838 523460 222844
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 522028 220516 522080 220522
rect 522028 220458 522080 220464
rect 522304 220516 522356 220522
rect 522304 220458 522356 220464
rect 522040 219774 522068 220458
rect 522028 219768 522080 219774
rect 522580 219768 522632 219774
rect 522028 219710 522080 219716
rect 522578 219736 522580 219745
rect 522632 219736 522634 219745
rect 522578 219671 522634 219680
rect 522592 217138 522620 219671
rect 523420 217530 523448 222838
rect 523408 217524 523460 217530
rect 523408 217466 523460 217472
rect 523420 217138 523448 217466
rect 524248 217138 524276 223246
rect 524420 219020 524472 219026
rect 524420 218962 524472 218968
rect 524432 218210 524460 218962
rect 525076 218754 525104 227122
rect 525720 224398 525748 229894
rect 526272 228954 526300 231676
rect 526916 230382 526944 231676
rect 526904 230376 526956 230382
rect 526904 230318 526956 230324
rect 526260 228948 526312 228954
rect 526260 228890 526312 228896
rect 525892 228404 525944 228410
rect 525892 228346 525944 228352
rect 525708 224392 525760 224398
rect 525708 224334 525760 224340
rect 525904 222018 525932 228346
rect 527560 225758 527588 231676
rect 528008 230444 528060 230450
rect 528008 230386 528060 230392
rect 527824 230376 527876 230382
rect 527824 230318 527876 230324
rect 526352 225752 526404 225758
rect 526352 225694 526404 225700
rect 527548 225752 527600 225758
rect 527548 225694 527600 225700
rect 526364 224954 526392 225694
rect 526364 224926 526760 224954
rect 525892 222012 525944 222018
rect 525892 221954 525944 221960
rect 524604 218748 524656 218754
rect 524604 218690 524656 218696
rect 525064 218748 525116 218754
rect 525064 218690 525116 218696
rect 524420 218204 524472 218210
rect 524420 218146 524472 218152
rect 524616 217734 524644 218690
rect 524604 217728 524656 217734
rect 524604 217670 524656 217676
rect 525076 217274 525104 218690
rect 525904 217274 525932 221954
rect 526442 220008 526498 220017
rect 526442 219943 526498 219952
rect 526456 218890 526484 219943
rect 526444 218884 526496 218890
rect 526444 218826 526496 218832
rect 526732 217274 526760 224926
rect 527548 220652 527600 220658
rect 527548 220594 527600 220600
rect 527560 218482 527588 220594
rect 527836 220114 527864 230318
rect 528020 230042 528048 230386
rect 528008 230036 528060 230042
rect 528008 229978 528060 229984
rect 528204 225894 528232 231676
rect 528848 230314 528876 231676
rect 529506 231662 529796 231690
rect 529020 230444 529072 230450
rect 529020 230386 529072 230392
rect 528836 230308 528888 230314
rect 528836 230250 528888 230256
rect 528192 225888 528244 225894
rect 528192 225830 528244 225836
rect 528376 224528 528428 224534
rect 528376 224470 528428 224476
rect 527824 220108 527876 220114
rect 527824 220050 527876 220056
rect 527548 218476 527600 218482
rect 527548 218418 527600 218424
rect 525076 217246 525150 217274
rect 525904 217246 525978 217274
rect 526732 217246 526806 217274
rect 520970 217116 521022 217122
rect 521764 217110 521838 217138
rect 522592 217110 522666 217138
rect 523420 217110 523494 217138
rect 524248 217110 524322 217138
rect 520970 217058 521022 217064
rect 520982 216988 521010 217058
rect 521810 216988 521838 217110
rect 522638 216988 522666 217110
rect 523466 216988 523494 217110
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527560 217138 527588 218418
rect 528388 217870 528416 224470
rect 529032 223310 529060 230386
rect 529204 224256 529256 224262
rect 529204 224198 529256 224204
rect 529020 223304 529072 223310
rect 529020 223246 529072 223252
rect 528376 217864 528428 217870
rect 528376 217806 528428 217812
rect 528388 217138 528416 217806
rect 529216 217138 529244 224198
rect 529768 221610 529796 231662
rect 529940 230172 529992 230178
rect 529940 230114 529992 230120
rect 529952 226302 529980 230114
rect 529940 226296 529992 226302
rect 529940 226238 529992 226244
rect 530136 224534 530164 231676
rect 530780 230042 530808 231676
rect 530768 230036 530820 230042
rect 530768 229978 530820 229984
rect 531424 228546 531452 231676
rect 531412 228540 531464 228546
rect 531412 228482 531464 228488
rect 531688 226160 531740 226166
rect 531688 226102 531740 226108
rect 530952 225616 531004 225622
rect 530952 225558 531004 225564
rect 530124 224528 530176 224534
rect 530124 224470 530176 224476
rect 530032 223440 530084 223446
rect 530032 223382 530084 223388
rect 529756 221604 529808 221610
rect 529756 221546 529808 221552
rect 530044 220017 530072 223382
rect 530030 220008 530086 220017
rect 530030 219943 530086 219952
rect 529388 218748 529440 218754
rect 529388 218690 529440 218696
rect 529400 218346 529428 218690
rect 529388 218340 529440 218346
rect 529388 218282 529440 218288
rect 530044 217138 530072 219943
rect 530964 217274 530992 225558
rect 531320 224936 531372 224942
rect 531320 224878 531372 224884
rect 531332 219774 531360 224878
rect 531320 219768 531372 219774
rect 531320 219710 531372 219716
rect 530918 217246 530992 217274
rect 531700 217274 531728 226102
rect 532068 225622 532096 231676
rect 532712 229770 532740 231676
rect 533370 231662 533752 231690
rect 532700 229764 532752 229770
rect 532700 229706 532752 229712
rect 532424 229628 532476 229634
rect 532424 229570 532476 229576
rect 532056 225616 532108 225622
rect 532056 225558 532108 225564
rect 532436 224806 532464 229570
rect 532424 224800 532476 224806
rect 532424 224742 532476 224748
rect 533724 222902 533752 231662
rect 534000 228682 534028 231676
rect 534644 230450 534672 231676
rect 534632 230444 534684 230450
rect 534632 230386 534684 230392
rect 534724 229900 534776 229906
rect 534724 229842 534776 229848
rect 533988 228676 534040 228682
rect 533988 228618 534040 228624
rect 533896 228404 533948 228410
rect 533896 228346 533948 228352
rect 533712 222896 533764 222902
rect 533712 222838 533764 222844
rect 533710 220552 533766 220561
rect 533710 220487 533766 220496
rect 533724 220017 533752 220487
rect 533710 220008 533766 220017
rect 533710 219943 533766 219952
rect 532516 219768 532568 219774
rect 532516 219710 532568 219716
rect 531700 217246 531774 217274
rect 530918 217190 530946 217246
rect 530906 217184 530958 217190
rect 527560 217110 527634 217138
rect 528388 217110 528462 217138
rect 529216 217110 529290 217138
rect 530044 217110 530118 217138
rect 530906 217126 530958 217132
rect 527606 216988 527634 217110
rect 528434 216988 528462 217110
rect 529262 216988 529290 217110
rect 530090 216988 530118 217110
rect 530918 216988 530946 217126
rect 531746 216988 531774 217246
rect 532528 217138 532556 219710
rect 533908 218890 533936 228346
rect 534736 223174 534764 229842
rect 535288 224262 535316 231676
rect 535932 227186 535960 231676
rect 536576 230178 536604 231676
rect 536564 230172 536616 230178
rect 536564 230114 536616 230120
rect 535920 227180 535972 227186
rect 535920 227122 535972 227128
rect 537220 227050 537248 231676
rect 537864 228410 537892 231676
rect 538508 229906 538536 231676
rect 538692 231662 539166 231690
rect 538496 229900 538548 229906
rect 538496 229842 538548 229848
rect 537852 228404 537904 228410
rect 537852 228346 537904 228352
rect 537576 227724 537628 227730
rect 537576 227666 537628 227672
rect 536012 227044 536064 227050
rect 536012 226986 536064 226992
rect 537208 227044 537260 227050
rect 537208 226986 537260 226992
rect 536024 224954 536052 226986
rect 535932 224926 536052 224954
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 534172 223168 534224 223174
rect 534172 223110 534224 223116
rect 534724 223168 534776 223174
rect 534724 223110 534776 223116
rect 534184 219298 534212 223110
rect 535000 221876 535052 221882
rect 535000 221818 535052 221824
rect 534172 219292 534224 219298
rect 534172 219234 534224 219240
rect 534632 219292 534684 219298
rect 534632 219234 534684 219240
rect 533436 218884 533488 218890
rect 533436 218826 533488 218832
rect 533896 218884 533948 218890
rect 533896 218826 533948 218832
rect 533448 217326 533476 218826
rect 533620 218748 533672 218754
rect 533620 218690 533672 218696
rect 534356 218748 534408 218754
rect 534356 218690 534408 218696
rect 533632 217841 533660 218690
rect 533618 217832 533674 217841
rect 533618 217767 533674 217776
rect 534368 217734 534396 218690
rect 534356 217728 534408 217734
rect 533632 217654 534258 217682
rect 534356 217670 534408 217676
rect 533632 217598 533660 217654
rect 533620 217592 533672 217598
rect 534230 217580 534258 217654
rect 534230 217569 534488 217580
rect 534230 217560 534502 217569
rect 534230 217552 534446 217560
rect 533620 217534 533672 217540
rect 534446 217495 534502 217504
rect 533436 217320 533488 217326
rect 533436 217262 533488 217268
rect 533448 217138 533476 217262
rect 534644 217138 534672 219234
rect 535012 218754 535040 221818
rect 535184 219156 535236 219162
rect 535184 219098 535236 219104
rect 535000 218748 535052 218754
rect 535000 218690 535052 218696
rect 532528 217110 532602 217138
rect 532574 216988 532602 217110
rect 533402 217110 533476 217138
rect 534230 217110 534672 217138
rect 535012 217138 535040 218690
rect 535196 217598 535224 219098
rect 535932 217598 535960 224926
rect 536656 224664 536708 224670
rect 536656 224606 536708 224612
rect 535184 217592 535236 217598
rect 535184 217534 535236 217540
rect 535920 217592 535972 217598
rect 535920 217534 535972 217540
rect 535932 217274 535960 217534
rect 535886 217246 535960 217274
rect 535012 217110 535086 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217110
rect 535058 216988 535086 217110
rect 535886 216988 535914 217246
rect 536668 217138 536696 224606
rect 537588 218890 537616 227666
rect 538692 221474 538720 231662
rect 544200 230444 544252 230450
rect 544200 230386 544252 230392
rect 541624 230308 541676 230314
rect 541624 230250 541676 230256
rect 540244 229084 540296 229090
rect 540244 229026 540296 229032
rect 538864 227588 538916 227594
rect 538864 227530 538916 227536
rect 538680 221468 538732 221474
rect 538680 221410 538732 221416
rect 537576 218884 537628 218890
rect 537576 218826 537628 218832
rect 537588 217274 537616 218826
rect 538876 217598 538904 227530
rect 539968 220516 540020 220522
rect 539968 220458 540020 220464
rect 539140 220380 539192 220386
rect 539140 220322 539192 220328
rect 538864 217592 538916 217598
rect 538864 217534 538916 217540
rect 538876 217274 538904 217534
rect 537542 217246 537616 217274
rect 538370 217246 538904 217274
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 216988 538398 217246
rect 539152 217138 539180 220322
rect 539980 217138 540008 220458
rect 540256 219366 540284 229026
rect 541440 226024 541492 226030
rect 541440 225966 541492 225972
rect 541452 224954 541480 225966
rect 541636 224954 541664 230250
rect 543188 228812 543240 228818
rect 543188 228754 543240 228760
rect 541452 224926 541572 224954
rect 541636 224926 541756 224954
rect 540244 219360 540296 219366
rect 540244 219302 540296 219308
rect 540796 219360 540848 219366
rect 540796 219302 540848 219308
rect 540808 217138 540836 219302
rect 541544 217274 541572 224926
rect 541728 220658 541756 224926
rect 542452 223304 542504 223310
rect 542452 223246 542504 223252
rect 542084 221128 542136 221134
rect 542084 221070 542136 221076
rect 541716 220652 541768 220658
rect 541716 220594 541768 220600
rect 541898 220552 541954 220561
rect 541898 220487 541954 220496
rect 541544 217246 541710 217274
rect 539152 217110 539226 217138
rect 539980 217110 540054 217138
rect 540808 217110 540882 217138
rect 539198 216988 539226 217110
rect 540026 216988 540054 217110
rect 540854 216988 540882 217110
rect 541682 216988 541710 217246
rect 541912 217190 541940 220487
rect 542096 217734 542124 221070
rect 542268 219904 542320 219910
rect 542268 219846 542320 219852
rect 542280 219366 542308 219846
rect 542464 219366 542492 223246
rect 543200 221882 543228 228754
rect 544212 226030 544240 230386
rect 549260 230172 549312 230178
rect 549260 230114 549312 230120
rect 547144 230036 547196 230042
rect 547144 229978 547196 229984
rect 545764 227316 545816 227322
rect 545764 227258 545816 227264
rect 544936 226296 544988 226302
rect 544936 226238 544988 226244
rect 544200 226024 544252 226030
rect 544200 225966 544252 225972
rect 542728 221876 542780 221882
rect 542728 221818 542780 221824
rect 543188 221876 543240 221882
rect 543188 221818 543240 221824
rect 542740 220814 542768 221818
rect 542740 220786 542860 220814
rect 542268 219360 542320 219366
rect 542268 219302 542320 219308
rect 542452 219360 542504 219366
rect 542452 219302 542504 219308
rect 542084 217728 542136 217734
rect 542084 217670 542136 217676
rect 542268 217728 542320 217734
rect 542268 217670 542320 217676
rect 542280 217462 542308 217670
rect 542268 217456 542320 217462
rect 542268 217398 542320 217404
rect 542464 217274 542492 219302
rect 542464 217246 542538 217274
rect 541900 217184 541952 217190
rect 541900 217126 541952 217132
rect 542510 216988 542538 217246
rect 542832 217172 542860 220786
rect 544658 220552 544714 220561
rect 543832 220516 543884 220522
rect 544658 220487 544714 220496
rect 543832 220458 543884 220464
rect 543844 220402 543872 220458
rect 543706 220374 543872 220402
rect 543706 220114 543734 220374
rect 544198 220280 544254 220289
rect 543832 220244 543884 220250
rect 543832 220186 543884 220192
rect 544016 220244 544068 220250
rect 544198 220215 544254 220224
rect 544016 220186 544068 220192
rect 543694 220108 543746 220114
rect 543694 220050 543746 220056
rect 543844 217818 543872 220186
rect 544028 219162 544056 220186
rect 544016 219156 544068 219162
rect 544016 219098 544068 219104
rect 544212 219026 544240 220215
rect 544476 219088 544528 219094
rect 544476 219030 544528 219036
rect 544200 219020 544252 219026
rect 544200 218962 544252 218968
rect 544488 218618 544516 219030
rect 544476 218612 544528 218618
rect 544476 218554 544528 218560
rect 543844 217790 544424 217818
rect 543004 217592 543056 217598
rect 543004 217534 543056 217540
rect 543016 217444 543044 217534
rect 543280 217456 543332 217462
rect 543016 217416 543280 217444
rect 544396 217410 544424 217790
rect 543280 217398 543332 217404
rect 544016 217388 544068 217394
rect 543384 217348 544016 217376
rect 543188 217320 543240 217326
rect 543384 217308 543412 217348
rect 544016 217330 544068 217336
rect 544304 217382 544424 217410
rect 544304 217308 544332 217382
rect 543240 217280 543412 217308
rect 544166 217280 544332 217308
rect 543188 217262 543240 217268
rect 543832 217252 543884 217258
rect 543832 217194 543884 217200
rect 543464 217184 543516 217190
rect 542832 217144 543366 217172
rect 543338 216988 543366 217144
rect 543844 217138 543872 217194
rect 543516 217132 543872 217138
rect 543464 217126 543872 217132
rect 543476 217110 543872 217126
rect 544166 216988 544194 217280
rect 544672 217190 544700 220487
rect 544948 219230 544976 226238
rect 545776 220998 545804 227258
rect 547156 221746 547184 229978
rect 547880 227452 547932 227458
rect 547880 227394 547932 227400
rect 547892 224954 547920 227394
rect 547892 224926 548932 224954
rect 547420 223168 547472 223174
rect 547420 223110 547472 223116
rect 546592 221740 546644 221746
rect 546592 221682 546644 221688
rect 547144 221740 547196 221746
rect 547144 221682 547196 221688
rect 545764 220992 545816 220998
rect 545764 220934 545816 220940
rect 544936 219224 544988 219230
rect 544936 219166 544988 219172
rect 544948 217274 544976 219166
rect 545776 217274 545804 220934
rect 545948 220652 546000 220658
rect 545948 220594 546000 220600
rect 545960 220504 545988 220594
rect 546316 220516 546368 220522
rect 545960 220476 546316 220504
rect 546316 220458 546368 220464
rect 544948 217246 545022 217274
rect 545776 217246 545850 217274
rect 544660 217184 544712 217190
rect 544660 217126 544712 217132
rect 544994 216988 545022 217246
rect 545822 216988 545850 217246
rect 546604 217138 546632 221682
rect 547432 220561 547460 223110
rect 548064 223032 548116 223038
rect 548064 222974 548116 222980
rect 548076 221270 548104 222974
rect 548064 221264 548116 221270
rect 548064 221206 548116 221212
rect 547418 220552 547474 220561
rect 547418 220487 547474 220496
rect 547432 217308 547460 220487
rect 548076 219994 548104 221206
rect 547892 219966 548104 219994
rect 547604 219904 547656 219910
rect 547604 219846 547656 219852
rect 547616 219201 547644 219846
rect 547892 219314 547920 219966
rect 547800 219286 547920 219314
rect 547602 219192 547658 219201
rect 547602 219127 547658 219136
rect 547800 218634 547828 219286
rect 548154 219192 548210 219201
rect 548154 219127 548210 219136
rect 547972 218748 548024 218754
rect 547972 218690 548024 218696
rect 547800 218606 547920 218634
rect 547432 217280 547506 217308
rect 546604 217110 546678 217138
rect 546650 216988 546678 217110
rect 547478 216988 547506 217280
rect 547892 217274 547920 218606
rect 547984 218090 548012 218690
rect 548168 218657 548196 219127
rect 548708 218748 548760 218754
rect 548708 218690 548760 218696
rect 548154 218648 548210 218657
rect 548154 218583 548210 218592
rect 548720 218210 548748 218690
rect 548904 218362 548932 224926
rect 549272 223038 549300 230114
rect 555436 230042 555464 251194
rect 558196 236094 558224 265610
rect 645872 261526 645900 277766
rect 647252 265674 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 265668 647292 265674
rect 647240 265610 647292 265616
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 567844 259480 567896 259486
rect 567844 259422 567896 259428
rect 562324 256760 562376 256766
rect 562324 256702 562376 256708
rect 559564 253428 559616 253434
rect 559564 253370 559616 253376
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 555424 230036 555476 230042
rect 555424 229978 555476 229984
rect 556804 229900 556856 229906
rect 556804 229842 556856 229848
rect 555608 229764 555660 229770
rect 555608 229706 555660 229712
rect 551652 228948 551704 228954
rect 551652 228890 551704 228896
rect 550456 224800 550508 224806
rect 550456 224742 550508 224748
rect 549260 223032 549312 223038
rect 549260 222974 549312 222980
rect 550468 221134 550496 224742
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 550652 221474 550680 224334
rect 550640 221468 550692 221474
rect 550640 221410 550692 221416
rect 549260 221128 549312 221134
rect 549260 221070 549312 221076
rect 550456 221128 550508 221134
rect 550456 221070 550508 221076
rect 549074 220552 549130 220561
rect 549074 220487 549130 220496
rect 549088 218890 549116 220487
rect 549076 218884 549128 218890
rect 549076 218826 549128 218832
rect 549272 218385 549300 221070
rect 550468 220114 550496 221070
rect 549996 220108 550048 220114
rect 549996 220050 550048 220056
rect 550456 220108 550508 220114
rect 550456 220050 550508 220056
rect 549444 220040 549496 220046
rect 549444 219982 549496 219988
rect 549258 218376 549314 218385
rect 548904 218334 549116 218362
rect 548708 218204 548760 218210
rect 548708 218146 548760 218152
rect 548892 218204 548944 218210
rect 548892 218146 548944 218152
rect 548904 218090 548932 218146
rect 547984 218062 548932 218090
rect 548432 217728 548484 217734
rect 548484 217676 548564 217682
rect 548432 217670 548564 217676
rect 548444 217654 548564 217670
rect 548536 217444 548564 217654
rect 548800 217456 548852 217462
rect 548536 217416 548800 217444
rect 548800 217398 548852 217404
rect 549088 217274 549116 218334
rect 549258 218311 549314 218320
rect 549456 217598 549484 219982
rect 549444 217592 549496 217598
rect 549444 217534 549496 217540
rect 547892 217246 548334 217274
rect 549088 217246 549162 217274
rect 548306 216988 548334 217246
rect 549134 216988 549162 217246
rect 550008 217138 550036 220050
rect 550652 217274 550680 221410
rect 551664 217274 551692 228890
rect 554044 225888 554096 225894
rect 554044 225830 554096 225836
rect 553308 225752 553360 225758
rect 553308 225694 553360 225700
rect 553320 224954 553348 225694
rect 553228 224926 553348 224954
rect 553228 222154 553256 224926
rect 554056 222194 554084 225830
rect 554056 222166 554452 222194
rect 553216 222148 553268 222154
rect 553216 222090 553268 222096
rect 552388 220652 552440 220658
rect 552388 220594 552440 220600
rect 550652 217246 550818 217274
rect 549962 217110 550036 217138
rect 549962 216988 549990 217110
rect 550790 216988 550818 217246
rect 551618 217246 551692 217274
rect 551618 216988 551646 217246
rect 552400 217138 552428 220594
rect 553228 217274 553256 222090
rect 554228 221128 554280 221134
rect 554228 221070 554280 221076
rect 553490 220552 553546 220561
rect 554240 220522 554268 221070
rect 553490 220487 553492 220496
rect 553544 220487 553546 220496
rect 554228 220516 554280 220522
rect 553492 220458 553544 220464
rect 554228 220458 554280 220464
rect 553492 220108 553544 220114
rect 553492 220050 553544 220056
rect 553504 219230 553532 220050
rect 553676 219904 553728 219910
rect 553676 219846 553728 219852
rect 553688 219586 553716 219846
rect 553688 219558 554084 219586
rect 553492 219224 553544 219230
rect 553492 219166 553544 219172
rect 553860 219020 553912 219026
rect 553504 218980 553860 219008
rect 553504 218210 553532 218980
rect 553860 218962 553912 218968
rect 554056 218385 554084 219558
rect 553674 218376 553730 218385
rect 553674 218311 553730 218320
rect 554042 218376 554098 218385
rect 554042 218311 554098 218320
rect 553688 218210 553716 218311
rect 553492 218204 553544 218210
rect 553492 218146 553544 218152
rect 553676 218204 553728 218210
rect 553676 218146 553728 218152
rect 554424 217274 554452 222166
rect 555422 222048 555478 222057
rect 555422 221983 555478 221992
rect 555436 221610 555464 221983
rect 555424 221604 555476 221610
rect 555424 221546 555476 221552
rect 554962 220552 555018 220561
rect 554962 220487 555018 220496
rect 554976 220114 555004 220487
rect 555238 220280 555294 220289
rect 555238 220215 555294 220224
rect 554964 220108 555016 220114
rect 554964 220050 555016 220056
rect 553228 217246 553302 217274
rect 552400 217110 552474 217138
rect 552446 216988 552474 217110
rect 553274 216988 553302 217246
rect 554102 217246 554452 217274
rect 554102 216988 554130 217246
rect 554976 217138 555004 220050
rect 555252 219026 555280 220215
rect 555240 219020 555292 219026
rect 555240 218962 555292 218968
rect 555436 217274 555464 221546
rect 555620 220697 555648 229706
rect 556528 224528 556580 224534
rect 556528 224470 556580 224476
rect 556068 221740 556120 221746
rect 556068 221682 556120 221688
rect 555606 220688 555662 220697
rect 555606 220623 555662 220632
rect 556080 220114 556108 221682
rect 556344 221604 556396 221610
rect 556344 221546 556396 221552
rect 556356 220114 556384 221546
rect 556068 220108 556120 220114
rect 556068 220050 556120 220056
rect 556344 220108 556396 220114
rect 556344 220050 556396 220056
rect 555608 219360 555660 219366
rect 555608 219302 555660 219308
rect 555792 219360 555844 219366
rect 555792 219302 555844 219308
rect 555620 219026 555648 219302
rect 555608 219020 555660 219026
rect 555608 218962 555660 218968
rect 555804 218754 555832 219302
rect 556160 218884 556212 218890
rect 556160 218826 556212 218832
rect 555792 218748 555844 218754
rect 555792 218690 555844 218696
rect 556172 218618 556200 218826
rect 556160 218612 556212 218618
rect 556160 218554 556212 218560
rect 555436 217246 555786 217274
rect 554930 217110 555004 217138
rect 554930 216988 554958 217110
rect 555758 216988 555786 217246
rect 556540 217138 556568 224470
rect 556816 221610 556844 229842
rect 558184 228540 558236 228546
rect 558184 228482 558236 228488
rect 558196 224954 558224 228482
rect 558920 225616 558972 225622
rect 558920 225558 558972 225564
rect 558012 224926 558224 224954
rect 558932 224954 558960 225558
rect 558932 224926 559052 224954
rect 557356 222420 557408 222426
rect 557356 222362 557408 222368
rect 556804 221604 556856 221610
rect 556804 221546 556856 221552
rect 557368 220114 557396 222362
rect 558012 222306 558040 224926
rect 558012 222278 558408 222306
rect 558012 220814 558040 222278
rect 558380 222154 558408 222278
rect 559024 222194 559052 224926
rect 558932 222166 559052 222194
rect 558184 222148 558236 222154
rect 558184 222090 558236 222096
rect 558368 222148 558420 222154
rect 558368 222090 558420 222096
rect 558196 221134 558224 222090
rect 558184 221128 558236 221134
rect 558184 221070 558236 221076
rect 557736 220786 558040 220814
rect 557540 220652 557592 220658
rect 557540 220594 557592 220600
rect 557552 220114 557580 220594
rect 557356 220108 557408 220114
rect 557356 220050 557408 220056
rect 557540 220108 557592 220114
rect 557540 220050 557592 220056
rect 557368 217138 557396 220050
rect 557736 219586 557764 220786
rect 558550 220688 558606 220697
rect 558550 220623 558552 220632
rect 558604 220623 558606 220632
rect 558552 220594 558604 220600
rect 558550 219736 558606 219745
rect 558550 219671 558606 219680
rect 558564 219586 558592 219671
rect 557552 219558 557764 219586
rect 558380 219558 558592 219586
rect 557552 217274 557580 219558
rect 557724 219496 557776 219502
rect 557724 219438 557776 219444
rect 557736 219008 557764 219438
rect 558380 219314 558408 219558
rect 558736 219496 558788 219502
rect 558736 219438 558788 219444
rect 558748 219314 558776 219438
rect 558288 219286 558408 219314
rect 558656 219286 558776 219314
rect 558288 219162 558316 219286
rect 558656 219212 558684 219286
rect 558472 219184 558684 219212
rect 558276 219156 558328 219162
rect 558276 219098 558328 219104
rect 558472 219008 558500 219184
rect 558736 219156 558788 219162
rect 558736 219098 558788 219104
rect 557736 218980 558500 219008
rect 558748 218634 558776 219098
rect 558564 218618 558776 218634
rect 558552 218612 558776 218618
rect 558604 218606 558776 218612
rect 558932 218634 558960 222166
rect 559576 220250 559604 253370
rect 561588 228676 561640 228682
rect 561588 228618 561640 228624
rect 560760 222896 560812 222902
rect 560760 222838 560812 222844
rect 559932 220652 559984 220658
rect 559932 220594 559984 220600
rect 559746 220552 559802 220561
rect 559746 220487 559802 220496
rect 559380 220244 559432 220250
rect 559380 220186 559432 220192
rect 559564 220244 559616 220250
rect 559564 220186 559616 220192
rect 559392 219745 559420 220186
rect 559102 219736 559158 219745
rect 559102 219671 559158 219680
rect 559378 219736 559434 219745
rect 559378 219671 559434 219680
rect 559116 218754 559144 219671
rect 559760 218890 559788 220487
rect 559748 218884 559800 218890
rect 559748 218826 559800 218832
rect 559104 218748 559156 218754
rect 559104 218690 559156 218696
rect 558932 218606 559144 218634
rect 558552 218554 558604 218560
rect 559116 217274 559144 218606
rect 557552 217246 558270 217274
rect 556540 217110 556614 217138
rect 557368 217110 557442 217138
rect 556586 216988 556614 217110
rect 557414 216988 557442 217110
rect 558242 216988 558270 217246
rect 559070 217246 559144 217274
rect 559070 216988 559098 217246
rect 559944 217138 559972 220594
rect 560772 217138 560800 222838
rect 561600 217274 561628 228618
rect 562336 226302 562364 256702
rect 566372 228404 566424 228410
rect 566372 228346 566424 228352
rect 564072 227180 564124 227186
rect 564072 227122 564124 227128
rect 562324 226296 562376 226302
rect 562324 226238 562376 226244
rect 561956 226024 562008 226030
rect 561956 225966 562008 225972
rect 561968 224954 561996 225966
rect 561968 224926 562272 224954
rect 562244 222329 562272 224926
rect 563704 224256 563756 224262
rect 563704 224198 563756 224204
rect 562968 222896 563020 222902
rect 562968 222838 563020 222844
rect 562416 222556 562468 222562
rect 562416 222498 562468 222504
rect 562230 222320 562286 222329
rect 562230 222255 562286 222264
rect 562046 220552 562102 220561
rect 562046 220487 562102 220496
rect 562060 217598 562088 220487
rect 562048 217592 562100 217598
rect 562048 217534 562100 217540
rect 559898 217110 559972 217138
rect 560726 217110 560800 217138
rect 561554 217246 561628 217274
rect 562244 217274 562272 222255
rect 562428 222154 562456 222498
rect 562784 222420 562836 222426
rect 562784 222362 562836 222368
rect 562416 222148 562468 222154
rect 562416 222090 562468 222096
rect 562598 222048 562654 222057
rect 562598 221983 562654 221992
rect 562612 221898 562640 221983
rect 562520 221870 562640 221898
rect 562520 217598 562548 221870
rect 562796 220130 562824 222362
rect 562980 222154 563008 222838
rect 563428 222420 563480 222426
rect 563428 222362 563480 222368
rect 562968 222148 563020 222154
rect 562968 222090 563020 222096
rect 563150 222048 563206 222057
rect 563150 221983 563206 221992
rect 562968 221740 563020 221746
rect 562968 221682 563020 221688
rect 562796 220102 562916 220130
rect 562692 219972 562744 219978
rect 562692 219914 562744 219920
rect 562704 218226 562732 219914
rect 562888 219910 562916 220102
rect 562980 219994 563008 221682
rect 563164 220402 563192 221983
rect 563440 221898 563468 222362
rect 563716 222194 563744 224198
rect 564084 222194 564112 227122
rect 565728 227044 565780 227050
rect 565728 226986 565780 226992
rect 564808 223032 564860 223038
rect 564808 222974 564860 222980
rect 564624 222828 564676 222834
rect 564624 222770 564676 222776
rect 563716 222166 563836 222194
rect 563072 220374 563192 220402
rect 563256 221870 563468 221898
rect 563072 220130 563100 220374
rect 563256 220250 563284 221870
rect 563808 221746 563836 222166
rect 563992 222166 564112 222194
rect 563796 221740 563848 221746
rect 563796 221682 563848 221688
rect 563426 220552 563482 220561
rect 563426 220487 563482 220496
rect 563244 220244 563296 220250
rect 563244 220186 563296 220192
rect 563440 220182 563468 220487
rect 563428 220176 563480 220182
rect 563072 220102 563192 220130
rect 563428 220118 563480 220124
rect 562980 219966 563100 219994
rect 562876 219904 562928 219910
rect 562876 219846 562928 219852
rect 562874 219736 562930 219745
rect 562874 219671 562930 219680
rect 562888 218754 562916 219671
rect 563072 219586 563100 219966
rect 562980 219558 563100 219586
rect 562980 219042 563008 219558
rect 563164 219042 563192 220102
rect 562980 219014 563192 219042
rect 562876 218748 562928 218754
rect 562876 218690 562928 218696
rect 563060 218748 563112 218754
rect 563060 218690 563112 218696
rect 562876 218612 562928 218618
rect 563072 218600 563100 218690
rect 562928 218572 563100 218600
rect 562876 218554 562928 218560
rect 563520 218476 563572 218482
rect 563520 218418 563572 218424
rect 563072 218334 563376 218362
rect 563072 218226 563100 218334
rect 562704 218198 563100 218226
rect 563348 218210 563376 218334
rect 563336 218204 563388 218210
rect 563336 218146 563388 218152
rect 563014 218136 563066 218142
rect 562874 218104 562930 218113
rect 563066 218084 563100 218090
rect 563014 218078 563100 218084
rect 563026 218062 563100 218078
rect 562874 218039 562930 218048
rect 562508 217592 562560 217598
rect 562508 217534 562560 217540
rect 562888 217546 562916 218039
rect 563072 217682 563100 218062
rect 563242 217696 563298 217705
rect 563072 217654 563242 217682
rect 563242 217631 563298 217640
rect 563532 217546 563560 218418
rect 562888 217518 563560 217546
rect 563808 217274 563836 221682
rect 562244 217246 562410 217274
rect 559898 216988 559926 217110
rect 560726 216988 560754 217110
rect 561554 216988 561582 217246
rect 562382 216988 562410 217246
rect 563210 217246 563836 217274
rect 563992 217274 564020 222166
rect 563992 217246 564066 217274
rect 563210 216988 563238 217246
rect 564038 216988 564066 217246
rect 564636 217190 564664 222770
rect 564820 222698 564848 222974
rect 564808 222692 564860 222698
rect 564808 222634 564860 222640
rect 564820 222194 564848 222634
rect 565740 222601 565768 226986
rect 565726 222592 565782 222601
rect 565726 222527 565782 222536
rect 564820 222166 564940 222194
rect 564912 217274 564940 222166
rect 566384 218226 566412 228346
rect 567856 224954 567884 259422
rect 568592 229094 568620 260850
rect 570616 234598 570644 261462
rect 571340 249076 571392 249082
rect 571340 249018 571392 249024
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 569960 230036 570012 230042
rect 569960 229978 570012 229984
rect 569972 229094 570000 229978
rect 571352 229094 571380 249018
rect 632704 246356 632756 246362
rect 632704 246298 632756 246304
rect 591304 245676 591356 245682
rect 591304 245618 591356 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 568592 229066 568988 229094
rect 569972 229066 570736 229094
rect 571352 229066 572300 229094
rect 568396 226296 568448 226302
rect 568396 226238 568448 226244
rect 568408 224954 568436 226238
rect 567856 224926 567976 224954
rect 567382 222592 567438 222601
rect 567382 222527 567438 222536
rect 567396 221746 567424 222527
rect 567568 222148 567620 222154
rect 567568 222090 567620 222096
rect 567752 222148 567804 222154
rect 567752 222090 567804 222096
rect 567580 221746 567608 222090
rect 567384 221740 567436 221746
rect 567384 221682 567436 221688
rect 567568 221740 567620 221746
rect 567568 221682 567620 221688
rect 567764 221610 567792 222090
rect 567476 221604 567528 221610
rect 567476 221546 567528 221552
rect 567752 221604 567804 221610
rect 567752 221546 567804 221552
rect 566568 220374 566964 220402
rect 566568 219230 566596 220374
rect 566936 220250 566964 220374
rect 566924 220244 566976 220250
rect 566924 220186 566976 220192
rect 566740 220176 566792 220182
rect 566740 220118 566792 220124
rect 566556 219224 566608 219230
rect 566556 219166 566608 219172
rect 566752 218498 566780 220118
rect 567016 219156 567068 219162
rect 567016 219098 567068 219104
rect 567028 218618 567056 219098
rect 567200 219020 567252 219026
rect 567200 218962 567252 218968
rect 567212 218618 567240 218962
rect 567016 218612 567068 218618
rect 567016 218554 567068 218560
rect 567200 218612 567252 218618
rect 567200 218554 567252 218560
rect 566752 218470 567240 218498
rect 566384 218198 566596 218226
rect 565280 217654 565860 217682
rect 565280 217326 565308 217654
rect 565680 217424 565736 217433
rect 565680 217359 565736 217368
rect 564866 217246 564940 217274
rect 565268 217320 565320 217326
rect 565268 217262 565320 217268
rect 564624 217184 564676 217190
rect 564624 217126 564676 217132
rect 564866 216988 564894 217246
rect 565694 216988 565722 217359
rect 565832 217326 565860 217654
rect 566002 217458 566058 217467
rect 566002 217393 566058 217402
rect 566188 217456 566240 217462
rect 566188 217398 566240 217404
rect 565820 217320 565872 217326
rect 565820 217262 565872 217268
rect 566016 217190 566044 217393
rect 566004 217184 566056 217190
rect 566004 217126 566056 217132
rect 566200 217122 566228 217398
rect 566568 217274 566596 218198
rect 567016 217456 567068 217462
rect 567016 217398 567068 217404
rect 566522 217246 566596 217274
rect 566188 217116 566240 217122
rect 566188 217058 566240 217064
rect 566522 216988 566550 217246
rect 567028 217122 567056 217398
rect 567212 217190 567240 218470
rect 567200 217184 567252 217190
rect 567488 217172 567516 221546
rect 567948 221270 567976 224926
rect 568316 224926 568436 224954
rect 568960 224954 568988 229066
rect 568960 224926 569816 224954
rect 568120 221604 568172 221610
rect 568120 221546 568172 221552
rect 567752 221264 567804 221270
rect 567752 221206 567804 221212
rect 567936 221264 567988 221270
rect 567936 221206 567988 221212
rect 567764 221082 567792 221206
rect 568132 221082 568160 221546
rect 567764 221054 568160 221082
rect 568026 219736 568082 219745
rect 568026 219671 568082 219680
rect 567844 219224 567896 219230
rect 567844 219166 567896 219172
rect 567856 218890 567884 219166
rect 568040 218890 568068 219671
rect 567844 218884 567896 218890
rect 567844 218826 567896 218832
rect 568028 218884 568080 218890
rect 568028 218826 568080 218832
rect 567200 217126 567252 217132
rect 567350 217144 567516 217172
rect 567016 217116 567068 217122
rect 567016 217058 567068 217064
rect 567350 216988 567378 217144
rect 568316 217104 568344 224926
rect 569316 222828 569368 222834
rect 569316 222770 569368 222776
rect 569132 222556 569184 222562
rect 569132 222498 569184 222504
rect 569144 221270 569172 222498
rect 568948 221264 569000 221270
rect 568948 221206 569000 221212
rect 569132 221264 569184 221270
rect 569132 221206 569184 221212
rect 568960 218464 568988 221206
rect 568960 218436 569264 218464
rect 569236 217274 569264 218436
rect 568178 217076 568344 217104
rect 569006 217246 569264 217274
rect 568178 216988 568206 217076
rect 569006 216988 569034 217246
rect 569328 217190 569356 222770
rect 569788 217274 569816 224926
rect 570708 217274 570736 229066
rect 572272 224954 572300 229066
rect 577516 224954 577544 240110
rect 591316 235278 591344 245618
rect 624424 244316 624476 244322
rect 624424 244258 624476 244264
rect 591304 235272 591356 235278
rect 591304 235214 591356 235220
rect 571628 224926 572300 224954
rect 577424 224926 577544 224954
rect 571432 222420 571484 222426
rect 571432 222362 571484 222368
rect 571248 220244 571300 220250
rect 571248 220186 571300 220192
rect 571260 218215 571288 220186
rect 571246 218206 571302 218215
rect 571246 218141 571302 218150
rect 569788 217246 569862 217274
rect 569316 217184 569368 217190
rect 569316 217126 569368 217132
rect 569834 216988 569862 217246
rect 570662 217246 570736 217274
rect 570662 216988 570690 217246
rect 571444 217138 571472 222362
rect 571628 222194 571656 224926
rect 572168 222692 572220 222698
rect 572168 222634 572220 222640
rect 571890 222320 571946 222329
rect 571890 222255 571946 222264
rect 571536 222166 571656 222194
rect 571536 218328 571564 222166
rect 571904 220250 571932 222255
rect 572180 222217 572208 222634
rect 572626 222592 572682 222601
rect 572626 222527 572682 222536
rect 572352 222420 572404 222426
rect 572352 222362 572404 222368
rect 572166 222208 572222 222217
rect 572364 222154 572392 222362
rect 572640 222154 572668 222527
rect 573180 222420 573232 222426
rect 573180 222362 573232 222368
rect 572166 222143 572222 222152
rect 572352 222148 572404 222154
rect 572352 222090 572404 222096
rect 572628 222148 572680 222154
rect 572628 222090 572680 222096
rect 572088 220646 572576 220674
rect 571892 220244 571944 220250
rect 571892 220186 571944 220192
rect 572088 219910 572116 220646
rect 572350 220552 572406 220561
rect 572350 220487 572406 220496
rect 572076 219904 572128 219910
rect 572076 219846 572128 219852
rect 572166 219736 572222 219745
rect 572166 219671 572222 219680
rect 571984 219360 572036 219366
rect 572180 219348 572208 219671
rect 572364 219450 572392 220487
rect 572548 220130 572576 220646
rect 572994 220144 573050 220153
rect 572548 220102 572994 220130
rect 572994 220079 573050 220088
rect 573192 219910 573220 222362
rect 575938 222184 575994 222193
rect 575938 222119 575994 222128
rect 573180 219904 573232 219910
rect 573180 219846 573232 219852
rect 572364 219422 573864 219450
rect 573836 219366 573864 219422
rect 573824 219360 573876 219366
rect 572180 219320 572668 219348
rect 571984 219302 572036 219308
rect 571996 219212 572024 219302
rect 571996 219184 572300 219212
rect 572272 219094 572300 219184
rect 572260 219088 572312 219094
rect 572260 219030 572312 219036
rect 571800 219020 571852 219026
rect 571800 218962 571852 218968
rect 571812 218498 571840 218962
rect 572640 218872 572668 219320
rect 572916 219286 573680 219314
rect 573824 219302 573876 219308
rect 575296 219360 575348 219366
rect 575296 219302 575348 219308
rect 572916 218958 572944 219286
rect 573272 219224 573324 219230
rect 573272 219166 573324 219172
rect 573456 219224 573508 219230
rect 573456 219166 573508 219172
rect 572904 218952 572956 218958
rect 572904 218894 572956 218900
rect 573088 218884 573140 218890
rect 572640 218844 572852 218872
rect 572076 218748 572128 218754
rect 572076 218690 572128 218696
rect 572444 218748 572496 218754
rect 572444 218690 572496 218696
rect 572088 218634 572116 218690
rect 572456 218634 572484 218690
rect 572088 218606 572484 218634
rect 572626 218648 572682 218657
rect 572626 218583 572682 218592
rect 571812 218470 572484 218498
rect 571892 218340 571944 218346
rect 571536 218300 571748 218328
rect 571720 217682 571748 218300
rect 571944 218300 572392 218328
rect 571892 218282 571944 218288
rect 571984 218204 572036 218210
rect 571984 218146 572036 218152
rect 572168 218204 572220 218210
rect 572168 218146 572220 218152
rect 571720 217654 571932 217682
rect 571904 217274 571932 217654
rect 571996 217546 572024 218146
rect 572180 217977 572208 218146
rect 572364 218090 572392 218300
rect 572456 218226 572484 218470
rect 572640 218362 572668 218583
rect 572824 218521 572852 218844
rect 573088 218826 573140 218832
rect 572810 218512 572866 218521
rect 572810 218447 572866 218456
rect 573100 218362 573128 218826
rect 572640 218334 573128 218362
rect 573284 218346 573312 219166
rect 573468 218482 573496 219166
rect 573652 218482 573680 219286
rect 574560 219088 574612 219094
rect 574560 219030 574612 219036
rect 573456 218476 573508 218482
rect 573456 218418 573508 218424
rect 573640 218476 573692 218482
rect 573640 218418 573692 218424
rect 574572 218346 574600 219030
rect 574744 219020 574796 219026
rect 574744 218962 574796 218968
rect 574756 218351 574784 218962
rect 575112 218748 575164 218754
rect 575112 218690 575164 218696
rect 573272 218340 573324 218346
rect 573272 218282 573324 218288
rect 574376 218340 574428 218346
rect 574376 218282 574428 218288
rect 574560 218340 574612 218346
rect 574560 218282 574612 218288
rect 574742 218342 574798 218351
rect 574388 218226 574416 218282
rect 574742 218277 574798 218286
rect 572456 218198 573128 218226
rect 574388 218198 574600 218226
rect 572364 218062 572760 218090
rect 572166 217968 572222 217977
rect 572166 217903 572222 217912
rect 572442 217560 572498 217569
rect 571996 217518 572442 217546
rect 572442 217495 572498 217504
rect 571904 217246 572346 217274
rect 571444 217110 571518 217138
rect 571490 216988 571518 217110
rect 572318 216988 572346 217246
rect 572732 217138 572760 218062
rect 573100 217410 573128 218198
rect 574572 218192 574600 218198
rect 574928 218204 574980 218210
rect 574572 218164 574784 218192
rect 574466 218104 574522 218113
rect 574466 218039 574522 218048
rect 574282 217560 574338 217569
rect 574282 217495 574338 217504
rect 573100 217382 574140 217410
rect 572732 217110 574048 217138
rect 574020 216492 574048 217110
rect 574112 216730 574140 217382
rect 574296 216918 574324 217495
rect 574480 217274 574508 218039
rect 574480 217246 574600 217274
rect 574284 216912 574336 216918
rect 574284 216854 574336 216860
rect 574572 216782 574600 217246
rect 574560 216776 574612 216782
rect 574112 216702 574232 216730
rect 574560 216718 574612 216724
rect 574204 216646 574232 216702
rect 574192 216640 574244 216646
rect 574192 216582 574244 216588
rect 574020 216464 574324 216492
rect 574296 215150 574324 216464
rect 574756 215286 574784 218164
rect 574928 218146 574980 218152
rect 574940 217569 574968 218146
rect 574926 217560 574982 217569
rect 574926 217495 574982 217504
rect 574928 216912 574980 216918
rect 574928 216854 574980 216860
rect 574744 215280 574796 215286
rect 574744 215222 574796 215228
rect 574284 215144 574336 215150
rect 574284 215086 574336 215092
rect 574940 213246 574968 216854
rect 575124 214878 575152 218690
rect 575112 214872 575164 214878
rect 575112 214814 575164 214820
rect 575308 213654 575336 219302
rect 575664 216776 575716 216782
rect 575664 216718 575716 216724
rect 575478 215112 575534 215121
rect 575478 215047 575534 215056
rect 575296 213648 575348 213654
rect 575296 213590 575348 213596
rect 575492 213518 575520 215047
rect 575676 214742 575704 216718
rect 575664 214736 575716 214742
rect 575664 214678 575716 214684
rect 575952 214606 575980 222119
rect 577424 217410 577452 224926
rect 593972 222284 594024 222290
rect 593972 222226 594024 222232
rect 577594 220688 577650 220697
rect 577594 220623 577650 220632
rect 577424 217382 577544 217410
rect 576124 216640 576176 216646
rect 576124 216582 576176 216588
rect 575940 214600 575992 214606
rect 575940 214542 575992 214548
rect 576136 214470 576164 216582
rect 576860 216504 576912 216510
rect 576860 216446 576912 216452
rect 576872 215121 576900 216446
rect 576858 215112 576914 215121
rect 576858 215047 576914 215056
rect 576306 214976 576362 214985
rect 576306 214911 576362 214920
rect 576124 214464 576176 214470
rect 576124 214406 576176 214412
rect 575480 213512 575532 213518
rect 575480 213454 575532 213460
rect 576320 213382 576348 214911
rect 576308 213376 576360 213382
rect 576308 213318 576360 213324
rect 574928 213240 574980 213246
rect 574928 213182 574980 213188
rect 577516 99346 577544 217382
rect 577608 215098 577636 220623
rect 582102 220144 582158 220153
rect 582102 220079 582158 220088
rect 582116 219994 582144 220079
rect 582116 219978 582420 219994
rect 582116 219972 582432 219978
rect 582116 219966 582380 219972
rect 582380 219914 582432 219920
rect 582196 219904 582248 219910
rect 582196 219846 582248 219852
rect 582208 219366 582236 219846
rect 582196 219360 582248 219366
rect 582196 219302 582248 219308
rect 582288 219224 582340 219230
rect 582102 219192 582158 219201
rect 582102 219127 582158 219136
rect 582286 219192 582288 219201
rect 582340 219192 582342 219201
rect 582286 219127 582342 219136
rect 586150 219192 586206 219201
rect 586150 219127 586206 219136
rect 586334 219192 586390 219201
rect 586334 219127 586390 219136
rect 582116 218906 582144 219127
rect 582116 218878 582374 218906
rect 582196 218748 582248 218754
rect 582196 218690 582248 218696
rect 582208 218521 582236 218690
rect 582346 218657 582374 218878
rect 582332 218648 582388 218657
rect 582332 218583 582388 218592
rect 582194 218512 582250 218521
rect 582194 218447 582250 218456
rect 586164 218090 586192 219127
rect 586348 218754 586376 219127
rect 586520 219020 586572 219026
rect 586520 218962 586572 218968
rect 586336 218748 586388 218754
rect 586336 218690 586388 218696
rect 586532 218385 586560 218962
rect 591672 218884 591724 218890
rect 591672 218826 591724 218832
rect 586518 218376 586574 218385
rect 586518 218311 586574 218320
rect 586334 218240 586390 218249
rect 586334 218175 586336 218184
rect 586388 218175 586390 218184
rect 586336 218146 586388 218152
rect 586518 218104 586574 218113
rect 586164 218062 586518 218090
rect 586518 218039 586574 218048
rect 591684 217841 591712 218826
rect 591486 217832 591542 217841
rect 591486 217767 591542 217776
rect 591670 217832 591726 217841
rect 591670 217767 591726 217776
rect 591026 217560 591082 217569
rect 591026 217495 591082 217504
rect 590842 217288 590898 217297
rect 590842 217223 590898 217232
rect 590856 216918 590884 217223
rect 590844 216912 590896 216918
rect 590844 216854 590896 216860
rect 590844 216776 590896 216782
rect 590842 216744 590844 216753
rect 591040 216753 591068 217495
rect 591500 217297 591528 217767
rect 591486 217288 591542 217297
rect 591486 217223 591542 217232
rect 592038 217016 592094 217025
rect 592038 216951 592094 216960
rect 592052 216782 592080 216951
rect 592040 216776 592092 216782
rect 590896 216744 590898 216753
rect 590842 216679 590898 216688
rect 591026 216744 591082 216753
rect 592040 216718 592092 216724
rect 591026 216679 591082 216688
rect 586704 216504 586756 216510
rect 586704 216446 586756 216452
rect 582102 215928 582158 215937
rect 582102 215863 582104 215872
rect 582156 215863 582158 215872
rect 582104 215834 582156 215840
rect 586716 215393 586744 216446
rect 586702 215384 586758 215393
rect 586702 215319 586758 215328
rect 577608 215070 577728 215098
rect 577700 215014 577728 215070
rect 577688 215008 577740 215014
rect 577688 214950 577740 214956
rect 578606 214024 578662 214033
rect 578606 213959 578662 213968
rect 578620 208350 578648 213959
rect 579434 211712 579490 211721
rect 579490 211670 579660 211698
rect 579434 211647 579490 211656
rect 578790 209944 578846 209953
rect 578790 209879 578792 209888
rect 578844 209879 578846 209888
rect 578792 209850 578844 209856
rect 578608 208344 578660 208350
rect 578608 208286 578660 208292
rect 579632 207670 579660 211670
rect 593984 210202 594012 222226
rect 600964 222148 601016 222154
rect 600964 222090 601016 222096
rect 607772 222148 607824 222154
rect 607772 222090 607824 222096
rect 597466 222048 597522 222057
rect 597466 221983 597468 221992
rect 597520 221983 597522 221992
rect 600596 222012 600648 222018
rect 597468 221954 597520 221960
rect 600596 221954 600648 221960
rect 597836 221876 597888 221882
rect 597836 221818 597888 221824
rect 597848 221610 597876 221818
rect 597836 221604 597888 221610
rect 597836 221546 597888 221552
rect 599490 221504 599546 221513
rect 599490 221439 599546 221448
rect 599030 220280 599086 220289
rect 599030 220215 599086 220224
rect 599044 219366 599072 220215
rect 599032 219360 599084 219366
rect 599032 219302 599084 219308
rect 597468 218612 597520 218618
rect 597468 218554 597520 218560
rect 594984 218204 595036 218210
rect 594984 218146 595036 218152
rect 596916 218204 596968 218210
rect 596916 218146 596968 218152
rect 594996 216918 595024 218146
rect 596928 217734 596956 218146
rect 596916 217728 596968 217734
rect 596916 217670 596968 217676
rect 597100 217728 597152 217734
rect 597100 217670 597152 217676
rect 597112 217462 597140 217670
rect 597100 217456 597152 217462
rect 597100 217398 597152 217404
rect 597480 217326 597508 218554
rect 597926 217560 597982 217569
rect 597926 217495 597982 217504
rect 597100 217320 597152 217326
rect 597100 217262 597152 217268
rect 597468 217320 597520 217326
rect 597468 217262 597520 217268
rect 595166 217016 595222 217025
rect 595166 216951 595222 216960
rect 594800 216912 594852 216918
rect 594800 216854 594852 216860
rect 594984 216912 595036 216918
rect 594984 216854 595036 216860
rect 594812 210202 594840 216854
rect 595180 210202 595208 216951
rect 597112 216782 597140 217262
rect 595628 216776 595680 216782
rect 595626 216744 595628 216753
rect 596272 216776 596324 216782
rect 595680 216744 595682 216753
rect 595626 216679 595682 216688
rect 595810 216744 595866 216753
rect 596272 216718 596324 216724
rect 597100 216776 597152 216782
rect 597100 216718 597152 216724
rect 595810 216679 595866 216688
rect 595824 215393 595852 216679
rect 595994 216472 596050 216481
rect 595994 216407 595996 216416
rect 596048 216407 596050 216416
rect 595996 216378 596048 216384
rect 595996 215892 596048 215898
rect 595996 215834 596048 215840
rect 596008 215393 596036 215834
rect 595810 215384 595866 215393
rect 595810 215319 595866 215328
rect 595994 215384 596050 215393
rect 595994 215319 596050 215328
rect 595718 215112 595774 215121
rect 595718 215047 595774 215056
rect 595732 210202 595760 215047
rect 596284 210202 596312 216718
rect 597558 216608 597614 216617
rect 597558 216543 597614 216552
rect 596824 216436 596876 216442
rect 596824 216378 596876 216384
rect 596836 210202 596864 216378
rect 597572 210202 597600 216543
rect 597940 210202 597968 217495
rect 598478 217288 598534 217297
rect 598478 217223 598534 217232
rect 598492 210202 598520 217223
rect 598848 217184 598900 217190
rect 598848 217126 598900 217132
rect 598860 216918 598888 217126
rect 598848 216912 598900 216918
rect 598848 216854 598900 216860
rect 599030 216200 599086 216209
rect 599030 216135 599086 216144
rect 599044 210202 599072 216135
rect 599504 210202 599532 221439
rect 600608 220862 600636 221954
rect 600976 221474 601004 222090
rect 602250 222048 602306 222057
rect 601148 222012 601200 222018
rect 602250 221983 602306 221992
rect 601148 221954 601200 221960
rect 601160 221474 601188 221954
rect 601332 221740 601384 221746
rect 601332 221682 601384 221688
rect 600964 221468 601016 221474
rect 600964 221410 601016 221416
rect 601148 221468 601200 221474
rect 601148 221410 601200 221416
rect 600778 221232 600834 221241
rect 600778 221167 600834 221176
rect 600412 220856 600464 220862
rect 600412 220798 600464 220804
rect 600596 220856 600648 220862
rect 600596 220798 600648 220804
rect 599766 219192 599822 219201
rect 599766 219127 599822 219136
rect 599780 215966 599808 219127
rect 599768 215960 599820 215966
rect 599768 215902 599820 215908
rect 600424 214334 600452 220798
rect 600792 219434 600820 221167
rect 601344 220998 601372 221682
rect 601332 220992 601384 220998
rect 601332 220934 601384 220940
rect 601976 220788 602028 220794
rect 601976 220730 602028 220736
rect 601790 220280 601846 220289
rect 601790 220215 601846 220224
rect 601804 219502 601832 220215
rect 601792 219496 601844 219502
rect 601792 219438 601844 219444
rect 600608 219406 600820 219434
rect 600412 214328 600464 214334
rect 600412 214270 600464 214276
rect 600608 210202 600636 219406
rect 601988 219366 602016 220730
rect 601976 219360 602028 219366
rect 601976 219302 602028 219308
rect 600962 218920 601018 218929
rect 600962 218855 601018 218864
rect 600976 218385 601004 218855
rect 600962 218376 601018 218385
rect 600962 218311 601018 218320
rect 601146 218376 601202 218385
rect 601146 218311 601202 218320
rect 601160 217841 601188 218311
rect 601332 218204 601384 218210
rect 601332 218146 601384 218152
rect 601146 217832 601202 217841
rect 601146 217767 601202 217776
rect 601344 217326 601372 218146
rect 601148 217320 601200 217326
rect 601148 217262 601200 217268
rect 601332 217320 601384 217326
rect 601332 217262 601384 217268
rect 601160 217054 601188 217262
rect 601148 217048 601200 217054
rect 601148 216990 601200 216996
rect 600962 216200 601018 216209
rect 600962 216135 601018 216144
rect 600976 215393 601004 216135
rect 600962 215384 601018 215393
rect 600962 215319 601018 215328
rect 600780 214328 600832 214334
rect 600780 214270 600832 214276
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596284 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600636 210202
rect 600792 210202 600820 214270
rect 601792 213648 601844 213654
rect 601792 213590 601844 213596
rect 601240 213512 601292 213518
rect 601240 213454 601292 213460
rect 601252 210202 601280 213454
rect 601804 210202 601832 213590
rect 602264 210202 602292 221983
rect 607312 221876 607364 221882
rect 607312 221818 607364 221824
rect 606576 221740 606628 221746
rect 606576 221682 606628 221688
rect 606024 220992 606076 220998
rect 606024 220934 606076 220940
rect 604090 219192 604146 219201
rect 604090 219127 604146 219136
rect 604104 217870 604132 219127
rect 605288 218340 605340 218346
rect 605288 218282 605340 218288
rect 602896 217864 602948 217870
rect 602896 217806 602948 217812
rect 604092 217864 604144 217870
rect 604092 217806 604144 217812
rect 602908 212534 602936 217806
rect 605300 217734 605328 218282
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 605288 217728 605340 217734
rect 605288 217670 605340 217676
rect 603448 217456 603500 217462
rect 603448 217398 603500 217404
rect 602908 212506 603120 212534
rect 603092 210202 603120 212506
rect 603460 210202 603488 217398
rect 604000 216776 604052 216782
rect 604000 216718 604052 216724
rect 604012 210202 604040 216718
rect 604472 210202 604500 217670
rect 605104 217320 605156 217326
rect 605104 217262 605156 217268
rect 605116 210202 605144 217262
rect 605840 216912 605892 216918
rect 605840 216854 605892 216860
rect 605852 210202 605880 216854
rect 606036 210338 606064 220934
rect 606588 219586 606616 221682
rect 606758 220280 606814 220289
rect 606758 220215 606814 220224
rect 606772 219745 606800 220215
rect 606758 219736 606814 219745
rect 606758 219671 606814 219680
rect 606588 219558 606708 219586
rect 606484 218476 606536 218482
rect 606484 218418 606536 218424
rect 606496 217326 606524 218418
rect 606484 217320 606536 217326
rect 606484 217262 606536 217268
rect 606036 210310 606156 210338
rect 606128 210202 606156 210310
rect 606680 210202 606708 219558
rect 607324 210202 607352 221818
rect 607784 210202 607812 222090
rect 616878 221776 616934 221785
rect 616878 221711 616934 221720
rect 610256 221604 610308 221610
rect 610256 221546 610308 221552
rect 610072 221468 610124 221474
rect 610072 221410 610124 221416
rect 608692 221264 608744 221270
rect 608692 221206 608744 221212
rect 608704 214334 608732 221206
rect 608876 221128 608928 221134
rect 608876 221070 608928 221076
rect 608692 214328 608744 214334
rect 608692 214270 608744 214276
rect 608888 210202 608916 221070
rect 609060 217592 609112 217598
rect 609060 217534 609112 217540
rect 600792 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602264 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604472 210174 604900 210202
rect 605116 210174 605452 210202
rect 605852 210174 606004 210202
rect 606128 210174 606556 210202
rect 606680 210174 607108 210202
rect 607324 210174 607660 210202
rect 607784 210174 608212 210202
rect 608764 210174 608916 210202
rect 609072 210202 609100 217534
rect 609520 214328 609572 214334
rect 609520 214270 609572 214276
rect 609532 210202 609560 214270
rect 610084 210322 610112 221410
rect 610072 210316 610124 210322
rect 610072 210258 610124 210264
rect 610268 210202 610296 221546
rect 611634 220960 611690 220969
rect 611634 220895 611690 220904
rect 611358 215928 611414 215937
rect 611358 215863 611414 215872
rect 610624 210316 610676 210322
rect 610624 210258 610676 210264
rect 610636 210202 610664 210258
rect 611372 210202 611400 215863
rect 611648 210202 611676 220895
rect 614486 218648 614542 218657
rect 614486 218583 614542 218592
rect 613844 218068 613896 218074
rect 613844 218010 613896 218016
rect 612280 217864 612332 217870
rect 612280 217806 612332 217812
rect 612292 210202 612320 217806
rect 613384 215960 613436 215966
rect 613384 215902 613436 215908
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 215902
rect 613856 215422 613884 218010
rect 614120 217184 614172 217190
rect 614120 217126 614172 217132
rect 613844 215416 613896 215422
rect 613844 215358 613896 215364
rect 614132 210202 614160 217126
rect 614500 210202 614528 218583
rect 615684 217728 615736 217734
rect 615684 217670 615736 217676
rect 615040 215416 615092 215422
rect 615040 215358 615092 215364
rect 615052 210202 615080 215358
rect 615696 210202 615724 217670
rect 616144 217320 616196 217326
rect 616144 217262 616196 217268
rect 616156 210202 616184 217262
rect 616892 214742 616920 221711
rect 617248 220788 617300 220794
rect 617248 220730 617300 220736
rect 617062 220008 617118 220017
rect 617062 219943 617118 219952
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616880 214736 616932 214742
rect 616880 214678 616932 214684
rect 616708 214334 616736 214678
rect 616696 214328 616748 214334
rect 616696 214270 616748 214276
rect 617076 210202 617104 219943
rect 609072 210174 609316 210202
rect 609532 210174 609868 210202
rect 610268 210174 610420 210202
rect 610636 210174 610972 210202
rect 611372 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 617044 210174 617104 210202
rect 617260 210202 617288 220730
rect 622676 220380 622728 220386
rect 622676 220322 622728 220328
rect 621020 219768 621072 219774
rect 621020 219710 621072 219716
rect 618260 219632 618312 219638
rect 618260 219574 618312 219580
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 219574
rect 620558 215928 620614 215937
rect 620558 215863 620614 215872
rect 618902 215656 618958 215665
rect 618902 215591 618958 215600
rect 618916 210202 618944 215591
rect 619640 215144 619692 215150
rect 619640 215086 619692 215092
rect 619652 210202 619680 215086
rect 620008 214464 620060 214470
rect 620008 214406 620060 214412
rect 620020 210202 620048 214406
rect 620572 210202 620600 215863
rect 621032 210202 621060 219710
rect 621664 215280 621716 215286
rect 621664 215222 621716 215228
rect 621676 210202 621704 215222
rect 622400 214872 622452 214878
rect 622400 214814 622452 214820
rect 622412 210202 622440 214814
rect 622688 210202 622716 220322
rect 623320 217048 623372 217054
rect 623320 216990 623372 216996
rect 623332 210202 623360 216990
rect 624436 214742 624464 244258
rect 628564 241528 628616 241534
rect 628564 241470 628616 241476
rect 628576 229094 628604 241470
rect 628576 229066 628696 229094
rect 626632 220652 626684 220658
rect 626632 220594 626684 220600
rect 625252 220516 625304 220522
rect 625252 220458 625304 220464
rect 625264 219434 625292 220458
rect 625436 220108 625488 220114
rect 625436 220050 625488 220056
rect 625264 219406 625384 219434
rect 624424 214736 624476 214742
rect 624424 214678 624476 214684
rect 624424 214328 624476 214334
rect 624424 214270 624476 214276
rect 623872 213240 623924 213246
rect 623872 213182 623924 213188
rect 623884 210202 623912 213182
rect 624436 210202 624464 214270
rect 625356 210202 625384 219406
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621032 210174 621460 210202
rect 621676 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625384 210202
rect 625448 210202 625476 220050
rect 626446 218104 626502 218113
rect 626446 218039 626502 218048
rect 626080 215008 626132 215014
rect 626080 214950 626132 214956
rect 626092 210202 626120 214950
rect 626460 213926 626488 218039
rect 626644 214606 626672 220594
rect 628012 220244 628064 220250
rect 628012 220186 628064 220192
rect 626816 219904 626868 219910
rect 626816 219846 626868 219852
rect 626632 214600 626684 214606
rect 626632 214542 626684 214548
rect 626448 213920 626500 213926
rect 626448 213862 626500 213868
rect 626828 210202 626856 219846
rect 627184 214600 627236 214606
rect 627184 214542 627236 214548
rect 627196 210202 627224 214542
rect 628024 210202 628052 220186
rect 628196 219496 628248 219502
rect 628196 219438 628248 219444
rect 628208 214554 628236 219438
rect 628208 214526 628512 214554
rect 628288 214464 628340 214470
rect 628288 214406 628340 214412
rect 628300 210202 628328 214406
rect 628484 210338 628512 214526
rect 628668 212770 628696 229066
rect 630954 219736 631010 219745
rect 630954 219671 631010 219680
rect 630770 219464 630826 219473
rect 630770 219399 630826 219408
rect 629942 218376 629998 218385
rect 629942 218311 629998 218320
rect 629392 213920 629444 213926
rect 629392 213862 629444 213868
rect 628656 212764 628708 212770
rect 628656 212706 628708 212712
rect 628484 210310 628788 210338
rect 628760 210202 628788 210310
rect 629404 210202 629432 213862
rect 629956 210202 629984 218311
rect 630784 214606 630812 219399
rect 630772 214600 630824 214606
rect 630772 214542 630824 214548
rect 630968 210202 630996 219671
rect 631138 218648 631194 218657
rect 631138 218583 631194 218592
rect 625448 210174 625876 210202
rect 626092 210174 626428 210202
rect 626828 210174 626980 210202
rect 627196 210174 627532 210202
rect 628024 210174 628084 210202
rect 628300 210174 628636 210202
rect 628760 210174 629188 210202
rect 629404 210174 629740 210202
rect 629956 210174 630292 210202
rect 630844 210174 630996 210202
rect 631152 210202 631180 218583
rect 631600 214600 631652 214606
rect 631600 214542 631652 214548
rect 631612 210202 631640 214542
rect 632716 212906 632744 246298
rect 648632 242214 648660 277366
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 633624 235272 633676 235278
rect 633624 235214 633676 235220
rect 632704 212900 632756 212906
rect 632704 212842 632756 212848
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 632716 210202 632744 212706
rect 633636 210202 633664 235214
rect 652036 232558 652064 378111
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652024 232552 652076 232558
rect 652024 232494 652076 232500
rect 640246 231432 640302 231441
rect 640246 231367 640302 231376
rect 639602 230072 639658 230081
rect 639602 230007 639658 230016
rect 638866 219192 638922 219201
rect 638866 219127 638922 219136
rect 636660 215348 636712 215354
rect 636660 215290 636712 215296
rect 633808 214736 633860 214742
rect 633808 214678 633860 214684
rect 631152 210174 631396 210202
rect 631612 210174 631948 210202
rect 632716 210174 633052 210202
rect 633604 210174 633664 210202
rect 633820 210202 633848 214678
rect 635556 213240 635608 213246
rect 635556 213182 635608 213188
rect 634360 212900 634412 212906
rect 634360 212842 634412 212848
rect 634372 210202 634400 212842
rect 635568 210202 635596 213182
rect 636672 210202 636700 215290
rect 638316 213920 638368 213926
rect 638316 213862 638368 213868
rect 637212 212764 637264 212770
rect 637212 212706 637264 212712
rect 637224 210202 637252 212706
rect 638328 210202 638356 213862
rect 638880 210202 638908 219127
rect 639616 215354 639644 230007
rect 640062 218920 640118 218929
rect 640062 218855 640118 218864
rect 639604 215348 639656 215354
rect 639604 215290 639656 215296
rect 640076 213926 640104 218855
rect 640064 213920 640116 213926
rect 640064 213862 640116 213868
rect 639972 213512 640024 213518
rect 639972 213454 640024 213460
rect 639984 210202 640012 213454
rect 640260 210202 640288 231367
rect 650642 223136 650698 223145
rect 650642 223071 650698 223080
rect 643190 220416 643246 220425
rect 643190 220351 643246 220360
rect 641442 220144 641498 220153
rect 641442 220079 641498 220088
rect 641456 212770 641484 220079
rect 642086 217288 642142 217297
rect 642086 217223 642142 217232
rect 642100 213518 642128 217223
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 642088 213512 642140 213518
rect 642088 213454 642140 213460
rect 641628 213376 641680 213382
rect 641628 213318 641680 213324
rect 641444 212764 641496 212770
rect 641444 212706 641496 212712
rect 641640 210202 641668 213318
rect 642178 213208 642234 213217
rect 642178 213143 642234 213152
rect 642192 210202 642220 213143
rect 643020 210202 643048 215863
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637252 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643204 210202 643232 220351
rect 647240 220108 647292 220114
rect 647240 220050 647292 220056
rect 644938 217560 644994 217569
rect 644938 217495 644994 217504
rect 644952 210202 644980 217495
rect 646594 215656 646650 215665
rect 646594 215591 646650 215600
rect 645492 213784 645544 213790
rect 645492 213726 645544 213732
rect 645504 210202 645532 213726
rect 646608 210202 646636 215591
rect 647252 214690 647280 220050
rect 649906 218648 649962 218657
rect 649906 218583 649962 218592
rect 647252 214662 647556 214690
rect 647146 214568 647202 214577
rect 647146 214503 647202 214512
rect 647160 210202 647188 214503
rect 643204 210174 643540 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647528 210202 647556 214662
rect 648528 213920 648580 213926
rect 648528 213862 648580 213868
rect 648540 210202 648568 213862
rect 649920 210202 649948 218583
rect 650656 213926 650684 223071
rect 651838 222864 651894 222873
rect 651838 222799 651894 222808
rect 651194 221504 651250 221513
rect 651194 221439 651250 221448
rect 651010 214840 651066 214849
rect 651010 214775 651066 214784
rect 650644 213920 650696 213926
rect 650644 213862 650696 213868
rect 650460 213512 650512 213518
rect 650460 213454 650512 213460
rect 650472 210202 650500 213454
rect 647528 210174 647956 210202
rect 648508 210174 648568 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651024 210202 651052 214775
rect 651208 213790 651236 221439
rect 651196 213784 651248 213790
rect 651196 213726 651248 213732
rect 651852 213246 651880 222799
rect 652024 213648 652076 213654
rect 652024 213590 652076 213596
rect 651840 213240 651892 213246
rect 651840 213182 651892 213188
rect 652036 210202 652064 213590
rect 651024 210174 651268 210202
rect 651820 210174 652064 210202
rect 581000 209908 581052 209914
rect 581000 209850 581052 209856
rect 579620 207664 579672 207670
rect 579620 207606 579672 207612
rect 579434 207360 579490 207369
rect 579490 207318 579660 207346
rect 579434 207295 579490 207304
rect 578238 205864 578294 205873
rect 578238 205799 578240 205808
rect 578292 205799 578294 205808
rect 578240 205770 578292 205776
rect 579632 205634 579660 207318
rect 581012 206310 581040 209850
rect 652220 209574 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 405657 660344 550598
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661684 416832 661736 416838
rect 661684 416774 661736 416780
rect 660302 405648 660358 405657
rect 660302 405583 660358 405592
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 661696 268161 661724 416774
rect 661880 406337 661908 522990
rect 662064 492017 662092 590650
rect 664456 579737 664484 709310
rect 665836 626113 665864 749362
rect 666296 705537 666324 776999
rect 666466 742792 666522 742801
rect 666466 742727 666522 742736
rect 666282 705528 666338 705537
rect 666282 705463 666338 705472
rect 666480 665417 666508 742727
rect 667216 671129 667244 803150
rect 667754 786720 667810 786729
rect 667754 786655 667810 786664
rect 667570 743200 667626 743209
rect 667570 743135 667626 743144
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 667584 665961 667612 743135
rect 667768 710841 667796 786655
rect 668228 752321 668256 868119
rect 668584 789404 668636 789410
rect 668584 789346 668636 789352
rect 668398 783864 668454 783873
rect 668398 783799 668454 783808
rect 668214 752312 668270 752321
rect 668214 752247 668270 752256
rect 668214 733680 668270 733689
rect 668214 733615 668270 733624
rect 667754 710832 667810 710841
rect 667754 710767 667810 710776
rect 667754 688936 667810 688945
rect 667754 688871 667810 688880
rect 667570 665952 667626 665961
rect 667570 665887 667626 665896
rect 666466 665408 666522 665417
rect 666466 665343 666522 665352
rect 667204 629332 667256 629338
rect 667204 629274 667256 629280
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 664628 603152 664680 603158
rect 664628 603094 664680 603100
rect 666466 603120 666522 603129
rect 664442 579728 664498 579737
rect 664442 579663 664498 579672
rect 664640 494057 664668 603094
rect 666466 603055 666522 603064
rect 666008 576904 666060 576910
rect 666008 576846 666060 576852
rect 665824 494760 665876 494766
rect 666020 494737 666048 576846
rect 666480 529961 666508 603055
rect 667216 534177 667244 629274
rect 667768 621217 667796 688871
rect 668228 662561 668256 733615
rect 668412 708801 668440 783799
rect 668398 708792 668454 708801
rect 668398 708727 668454 708736
rect 668398 692880 668454 692889
rect 668398 692815 668454 692824
rect 668214 662552 668270 662561
rect 668214 662487 668270 662496
rect 668214 654256 668270 654265
rect 668214 654191 668270 654200
rect 667754 621208 667810 621217
rect 667754 621143 667810 621152
rect 668228 574161 668256 654191
rect 668412 620265 668440 692815
rect 668596 670585 668624 789346
rect 668768 775600 668820 775606
rect 668768 775542 668820 775548
rect 668780 734369 668808 775542
rect 668950 773800 669006 773809
rect 668950 773735 669006 773744
rect 668766 734360 668822 734369
rect 668766 734295 668822 734304
rect 668766 731504 668822 731513
rect 668766 731439 668822 731448
rect 668582 670576 668638 670585
rect 668582 670511 668638 670520
rect 668780 664601 668808 731439
rect 668964 710025 668992 773735
rect 669240 755177 669268 879135
rect 671158 872264 671214 872273
rect 671158 872199 671214 872208
rect 670606 867912 670662 867921
rect 670606 867847 670662 867856
rect 669778 864240 669834 864249
rect 669778 864175 669834 864184
rect 669594 789440 669650 789449
rect 669594 789375 669650 789384
rect 669226 755168 669282 755177
rect 669226 755103 669282 755112
rect 669410 741160 669466 741169
rect 669410 741095 669466 741104
rect 668950 710016 669006 710025
rect 668950 709951 669006 709960
rect 669226 705120 669282 705129
rect 669226 705055 669282 705064
rect 668766 664592 668822 664601
rect 668766 664527 668822 664536
rect 669042 648680 669098 648689
rect 669042 648615 669098 648624
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668398 620256 668454 620265
rect 668398 620191 668454 620200
rect 668398 601760 668454 601769
rect 668398 601695 668454 601704
rect 668214 574152 668270 574161
rect 668214 574087 668270 574096
rect 668214 564496 668270 564505
rect 668214 564431 668270 564440
rect 667202 534168 667258 534177
rect 667202 534103 667258 534112
rect 666466 529952 666522 529961
rect 666466 529887 666522 529896
rect 665824 494702 665876 494708
rect 666006 494728 666062 494737
rect 664626 494048 664682 494057
rect 664626 493983 664682 493992
rect 662050 492008 662106 492017
rect 662050 491943 662106 491952
rect 663064 470620 663116 470626
rect 663064 470562 663116 470568
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 663076 315489 663104 470562
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663248 364404 663300 364410
rect 663248 364346 663300 364352
rect 663062 315480 663118 315489
rect 663062 315415 663118 315424
rect 661682 268152 661738 268161
rect 661682 268087 661738 268096
rect 663260 234161 663288 364346
rect 664456 271153 664484 404330
rect 665836 358737 665864 494702
rect 666006 494663 666062 494672
rect 668228 485217 668256 564431
rect 668412 526561 668440 601695
rect 668596 535945 668624 643078
rect 668858 593736 668914 593745
rect 668858 593671 668914 593680
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668872 528601 668900 593671
rect 669056 573209 669084 648615
rect 669042 573200 669098 573209
rect 669042 573135 669098 573144
rect 669042 559056 669098 559065
rect 669042 558991 669098 559000
rect 668858 528592 668914 528601
rect 668858 528527 668914 528536
rect 668398 526552 668454 526561
rect 668398 526487 668454 526496
rect 668214 485208 668270 485217
rect 668214 485143 668270 485152
rect 668768 484424 668820 484430
rect 668768 484366 668820 484372
rect 667204 456816 667256 456822
rect 667204 456758 667256 456764
rect 665822 358728 665878 358737
rect 665822 358663 665878 358672
rect 666192 338156 666244 338162
rect 666192 338098 666244 338104
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 663246 234152 663302 234161
rect 663246 234087 663302 234096
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 662328 232348 662380 232354
rect 662328 232290 662380 232296
rect 661682 229528 661738 229537
rect 661682 229463 661738 229472
rect 660946 229256 661002 229265
rect 660946 229191 661002 229200
rect 652758 226400 652814 226409
rect 652758 226335 652814 226344
rect 652772 220114 652800 226335
rect 654782 225584 654838 225593
rect 654782 225519 654838 225528
rect 654140 221468 654192 221474
rect 654140 221410 654192 221416
rect 653034 220688 653090 220697
rect 653034 220623 653090 220632
rect 652760 220108 652812 220114
rect 652760 220050 652812 220056
rect 652852 213240 652904 213246
rect 652852 213182 652904 213188
rect 652864 210202 652892 213182
rect 653048 210202 653076 220623
rect 654152 210202 654180 221410
rect 654796 213382 654824 225519
rect 655886 225312 655942 225321
rect 655886 225247 655942 225256
rect 655704 221604 655756 221610
rect 655704 221546 655756 221552
rect 655426 216472 655482 216481
rect 655426 216407 655482 216416
rect 654784 213376 654836 213382
rect 654784 213318 654836 213324
rect 655440 210202 655468 216407
rect 655716 213926 655744 221546
rect 655900 221474 655928 225247
rect 660210 225040 660266 225049
rect 660210 224975 660266 224984
rect 658186 224496 658242 224505
rect 658186 224431 658242 224440
rect 656622 223680 656678 223689
rect 656622 223615 656678 223624
rect 655888 221468 655940 221474
rect 655888 221410 655940 221416
rect 655704 213920 655756 213926
rect 655704 213862 655756 213868
rect 656636 210202 656664 223615
rect 658002 221776 658058 221785
rect 658002 221711 658058 221720
rect 656808 213920 656860 213926
rect 656808 213862 656860 213868
rect 656820 210202 656848 213862
rect 658016 213654 658044 221711
rect 658004 213648 658056 213654
rect 658004 213590 658056 213596
rect 658200 210202 658228 224431
rect 659566 223952 659622 223961
rect 659566 223887 659622 223896
rect 658922 223408 658978 223417
rect 658922 223343 658978 223352
rect 658740 214396 658792 214402
rect 658740 214338 658792 214344
rect 658752 210202 658780 214338
rect 658936 213518 658964 223343
rect 659580 221610 659608 223887
rect 659568 221604 659620 221610
rect 659568 221546 659620 221552
rect 659568 213648 659620 213654
rect 659568 213590 659620 213596
rect 658924 213512 658976 213518
rect 658924 213454 658976 213460
rect 659580 210202 659608 213590
rect 660224 213246 660252 224975
rect 660960 213926 660988 229191
rect 661696 214402 661724 229463
rect 662052 214600 662104 214606
rect 662052 214542 662104 214548
rect 661684 214396 661736 214402
rect 661684 214338 661736 214344
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 660212 213240 660264 213246
rect 660212 213182 660264 213188
rect 660408 210202 660436 213862
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660960 210202 660988 213726
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 214542
rect 662340 210202 662368 232290
rect 665088 232212 665140 232218
rect 665088 232154 665140 232160
rect 663062 231840 663118 231849
rect 663062 231775 663118 231784
rect 663076 219434 663104 231775
rect 663246 231160 663302 231169
rect 663246 231095 663302 231104
rect 662984 219406 663104 219434
rect 662984 213790 663012 219406
rect 663260 214606 663288 231095
rect 664442 230616 664498 230625
rect 664442 230551 664498 230560
rect 663708 227588 663760 227594
rect 663708 227530 663760 227536
rect 663524 214940 663576 214946
rect 663524 214882 663576 214888
rect 663248 214600 663300 214606
rect 663248 214542 663300 214548
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 662972 213784 663024 213790
rect 662972 213726 663024 213732
rect 663168 210202 663196 213862
rect 663536 210202 663564 214882
rect 663720 213926 663748 227530
rect 664456 214946 664484 230551
rect 664626 215112 664682 215121
rect 664626 215047 664682 215056
rect 664444 214940 664496 214946
rect 664444 214882 664496 214888
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664640 213654 664668 215047
rect 664810 213752 664866 213761
rect 664810 213687 664866 213696
rect 664628 213648 664680 213654
rect 664628 213590 664680 213596
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 213687
rect 665100 213042 665128 232154
rect 665546 230888 665602 230897
rect 665546 230823 665602 230832
rect 665560 227594 665588 230823
rect 665548 227588 665600 227594
rect 665548 227530 665600 227536
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654152 210174 654580 210202
rect 655132 210174 655468 210202
rect 656236 210174 656664 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652208 209568 652260 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652208 209510 652260 209516
rect 632164 209494 632500 209510
rect 591304 208684 591356 208690
rect 591304 208626 591356 208632
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 207664 589516 207670
rect 589464 207606 589516 207612
rect 589476 206417 589504 207606
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 581000 206304 581052 206310
rect 581000 206246 581052 206252
rect 589648 206304 589700 206310
rect 589648 206246 589700 206252
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579632 205606 579752 205634
rect 579724 204270 579752 205606
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 589660 204785 589688 206246
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 589648 186312 589700 186318
rect 579580 186280 579582 186289
rect 589648 186254 589700 186260
rect 579526 186215 579582 186224
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 578804 180169 578832 180746
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 578804 175137 578832 178026
rect 589660 177954 589688 180231
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 583024 175296 583076 175302
rect 583024 175238 583076 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 579526 171048 579582 171057
rect 579526 170983 579528 170992
rect 579580 170983 579582 170992
rect 579528 170954 579580 170960
rect 580920 169726 580948 172518
rect 581644 171148 581696 171154
rect 581644 171090 581696 171096
rect 578332 169720 578384 169726
rect 578332 169662 578384 169668
rect 580908 169720 580960 169726
rect 580908 169662 580960 169668
rect 578344 169289 578372 169662
rect 578330 169280 578386 169289
rect 578330 169215 578386 169224
rect 579620 168428 579672 168434
rect 579620 168370 579672 168376
rect 578976 167204 579028 167210
rect 578976 167146 579028 167152
rect 578988 166977 579016 167146
rect 578974 166968 579030 166977
rect 578974 166903 579030 166912
rect 578884 165572 578936 165578
rect 578884 165514 578936 165520
rect 578896 164529 578924 165514
rect 578882 164520 578938 164529
rect 578882 164455 578938 164464
rect 579434 162480 579490 162489
rect 579632 162466 579660 168370
rect 581656 167210 581684 171090
rect 583036 171018 583064 175238
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 583024 171012 583076 171018
rect 583024 170954 583076 170960
rect 589462 170504 589518 170513
rect 589462 170439 589518 170448
rect 589476 169794 589504 170439
rect 582380 169788 582432 169794
rect 582380 169730 582432 169736
rect 589464 169788 589516 169794
rect 589464 169730 589516 169736
rect 581644 167204 581696 167210
rect 581644 167146 581696 167152
rect 581644 167068 581696 167074
rect 581644 167010 581696 167016
rect 579490 162438 579660 162466
rect 579434 162415 579490 162424
rect 580264 161492 580316 161498
rect 580264 161434 580316 161440
rect 579252 160064 579304 160070
rect 579252 160006 579304 160012
rect 579264 159905 579292 160006
rect 579250 159896 579306 159905
rect 579250 159831 579306 159840
rect 579160 158704 579212 158710
rect 579160 158646 579212 158652
rect 579172 158273 579200 158646
rect 579158 158264 579214 158273
rect 579158 158199 579214 158208
rect 579526 155952 579582 155961
rect 579526 155887 579528 155896
rect 579580 155887 579582 155896
rect 579528 155858 579580 155864
rect 580276 154562 580304 161434
rect 581656 160070 581684 167010
rect 582392 165578 582420 169730
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589462 165608 589518 165617
rect 582380 165572 582432 165578
rect 589462 165543 589518 165552
rect 582380 165514 582432 165520
rect 589476 164286 589504 165543
rect 585968 164280 586020 164286
rect 585968 164222 586020 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 584404 162920 584456 162926
rect 584404 162862 584456 162868
rect 582380 160132 582432 160138
rect 582380 160074 582432 160080
rect 581644 160064 581696 160070
rect 581644 160006 581696 160012
rect 581828 158840 581880 158846
rect 581828 158782 581880 158788
rect 578240 154556 578292 154562
rect 578240 154498 578292 154504
rect 580264 154556 580316 154562
rect 580264 154498 580316 154504
rect 578252 154057 578280 154498
rect 578238 154048 578294 154057
rect 578238 153983 578294 153992
rect 580448 153264 580500 153270
rect 580448 153206 580500 153212
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 578252 151745 578280 152730
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 147416 579580 147422
rect 579528 147358 579580 147364
rect 579540 147257 579568 147358
rect 579526 147248 579582 147257
rect 579526 147183 579582 147192
rect 578884 145580 578936 145586
rect 578884 145522 578936 145528
rect 578608 143200 578660 143206
rect 578608 143142 578660 143148
rect 578620 143041 578648 143142
rect 578606 143032 578662 143041
rect 578606 142967 578662 142976
rect 578700 139392 578752 139398
rect 578700 139334 578752 139340
rect 578712 138825 578740 139334
rect 578698 138816 578754 138825
rect 578698 138751 578754 138760
rect 578896 136649 578924 145522
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 580460 143206 580488 153206
rect 581840 150618 581868 158782
rect 582392 152794 582420 160074
rect 584416 155922 584444 162862
rect 585980 158710 586008 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158846 589504 159015
rect 589464 158840 589516 158846
rect 589464 158782 589516 158788
rect 585968 158704 586020 158710
rect 585968 158646 586020 158652
rect 589462 157448 589518 157457
rect 585784 157412 585836 157418
rect 589462 157383 589464 157392
rect 585784 157354 585836 157360
rect 589516 157383 589518 157392
rect 589464 157354 589516 157360
rect 584404 155916 584456 155922
rect 584404 155858 584456 155864
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 582380 152788 582432 152794
rect 582380 152730 582432 152736
rect 583024 151836 583076 151842
rect 583024 151778 583076 151784
rect 581828 150612 581880 150618
rect 581828 150554 581880 150560
rect 581644 150476 581696 150482
rect 581644 150418 581696 150424
rect 580448 143200 580500 143206
rect 580448 143142 580500 143148
rect 580264 142180 580316 142186
rect 580264 142122 580316 142128
rect 579528 140616 579580 140622
rect 579526 140584 579528 140593
rect 579580 140584 579582 140593
rect 579526 140519 579582 140528
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 578332 135924 578384 135930
rect 578332 135866 578384 135872
rect 578344 134473 578372 135866
rect 578330 134464 578386 134473
rect 578330 134399 578386 134408
rect 578240 134292 578292 134298
rect 578240 134234 578292 134240
rect 578252 132297 578280 134234
rect 579252 133204 579304 133210
rect 579252 133146 579304 133152
rect 578238 132288 578294 132297
rect 578238 132223 578294 132232
rect 578332 128308 578384 128314
rect 578332 128250 578384 128256
rect 578344 127809 578372 128250
rect 578330 127800 578386 127809
rect 578330 127735 578386 127744
rect 579264 125361 579292 133146
rect 579528 129736 579580 129742
rect 579526 129704 579528 129713
rect 579580 129704 579582 129713
rect 579526 129639 579582 129648
rect 580276 128314 580304 142122
rect 581656 139398 581684 150418
rect 583036 140622 583064 151778
rect 584416 144702 584444 154566
rect 585796 147422 585824 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 589462 150920 589518 150929
rect 589462 150855 589518 150864
rect 589476 150482 589504 150855
rect 589464 150476 589516 150482
rect 589464 150418 589516 150424
rect 589186 149288 589242 149297
rect 589186 149223 589242 149232
rect 585784 147416 585836 147422
rect 585784 147358 585836 147364
rect 587348 146328 587400 146334
rect 587348 146270 587400 146276
rect 585784 144968 585836 144974
rect 585784 144910 585836 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 140616 583076 140622
rect 583024 140558 583076 140564
rect 584404 139460 584456 139466
rect 584404 139402 584456 139408
rect 581644 139392 581696 139398
rect 581644 139334 581696 139340
rect 581644 136672 581696 136678
rect 581644 136614 581696 136620
rect 580264 128308 580316 128314
rect 580264 128250 580316 128256
rect 580448 127016 580500 127022
rect 580448 126958 580500 126964
rect 579250 125352 579306 125361
rect 579250 125287 579306 125296
rect 579252 124160 579304 124166
rect 579252 124102 579304 124108
rect 579264 123593 579292 124102
rect 579250 123584 579306 123593
rect 579250 123519 579306 123528
rect 579252 122868 579304 122874
rect 579252 122810 579304 122816
rect 579068 121168 579120 121174
rect 579066 121136 579068 121145
rect 579120 121136 579122 121145
rect 579066 121071 579122 121080
rect 578516 118652 578568 118658
rect 578516 118594 578568 118600
rect 578528 118425 578556 118594
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 579068 115252 579120 115258
rect 579068 115194 579120 115200
rect 578332 108384 578384 108390
rect 578330 108352 578332 108361
rect 578384 108352 578386 108361
rect 578330 108287 578386 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578332 106548 578384 106554
rect 578332 106490 578384 106496
rect 578344 105913 578372 106490
rect 578330 105904 578386 105913
rect 578330 105839 578386 105848
rect 577504 99340 577556 99346
rect 577504 99282 577556 99288
rect 577504 95940 577556 95946
rect 577504 95882 577556 95888
rect 574928 56160 574980 56166
rect 574928 56102 574980 56108
rect 574560 56024 574612 56030
rect 574560 55966 574612 55972
rect 574572 53990 574600 55966
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 54126 574784 55830
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 56102
rect 577516 55214 577544 95882
rect 578516 93832 578568 93838
rect 578516 93774 578568 93780
rect 578528 93129 578556 93774
rect 578514 93120 578570 93129
rect 578514 93055 578570 93064
rect 578516 86760 578568 86766
rect 578516 86702 578568 86708
rect 578528 86465 578556 86702
rect 578514 86456 578570 86465
rect 578514 86391 578570 86400
rect 578896 80073 578924 107578
rect 579080 90953 579108 115194
rect 579264 101833 579292 122810
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579526 114472 579582 114481
rect 579526 114407 579528 114416
rect 579580 114407 579582 114416
rect 579528 114378 579580 114384
rect 579528 113144 579580 113150
rect 579528 113086 579580 113092
rect 579540 112713 579568 113086
rect 579526 112704 579582 112713
rect 579526 112639 579582 112648
rect 579436 110288 579488 110294
rect 579434 110256 579436 110265
rect 579488 110256 579490 110265
rect 579434 110191 579490 110200
rect 580264 106956 580316 106962
rect 580264 106898 580316 106904
rect 579528 103352 579580 103358
rect 579526 103320 579528 103329
rect 579580 103320 579582 103329
rect 579526 103255 579582 103264
rect 579250 101824 579306 101833
rect 579250 101759 579306 101768
rect 579526 99240 579582 99249
rect 579526 99175 579528 99184
rect 579580 99175 579582 99184
rect 579528 99146 579580 99152
rect 579528 97504 579580 97510
rect 579526 97472 579528 97481
rect 579580 97472 579582 97481
rect 579526 97407 579582 97416
rect 579528 95056 579580 95062
rect 579526 95024 579528 95033
rect 579580 95024 579582 95033
rect 579526 94959 579582 94968
rect 579066 90944 579122 90953
rect 579066 90879 579122 90888
rect 579068 89752 579120 89758
rect 579068 89694 579120 89700
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579080 77897 579108 89694
rect 579528 88324 579580 88330
rect 579528 88266 579580 88272
rect 579540 88097 579568 88266
rect 579526 88088 579582 88097
rect 579526 88023 579582 88032
rect 580276 86766 580304 106898
rect 580460 106554 580488 126958
rect 581656 121174 581684 136614
rect 582380 131776 582432 131782
rect 582380 131718 582432 131724
rect 582392 129742 582420 131718
rect 582380 129736 582432 129742
rect 582380 129678 582432 129684
rect 583024 128376 583076 128382
rect 583024 128318 583076 128324
rect 581644 121168 581696 121174
rect 581644 121110 581696 121116
rect 582012 120760 582064 120766
rect 582012 120702 582064 120708
rect 582024 110294 582052 120702
rect 582012 110288 582064 110294
rect 582012 110230 582064 110236
rect 581828 109744 581880 109750
rect 581828 109686 581880 109692
rect 580448 106548 580500 106554
rect 580448 106490 580500 106496
rect 580632 106344 580684 106350
rect 580632 106286 580684 106292
rect 580448 93152 580500 93158
rect 580448 93094 580500 93100
rect 580264 86760 580316 86766
rect 580264 86702 580316 86708
rect 579344 84040 579396 84046
rect 579342 84008 579344 84017
rect 579396 84008 579398 84017
rect 579342 83943 579398 83952
rect 579252 82816 579304 82822
rect 579252 82758 579304 82764
rect 579264 82249 579292 82758
rect 579250 82240 579306 82249
rect 579250 82175 579306 82184
rect 579252 80096 579304 80102
rect 579252 80038 579304 80044
rect 579066 77888 579122 77897
rect 579066 77823 579122 77832
rect 579264 77738 579292 80038
rect 579080 77710 579292 77738
rect 578884 77444 578936 77450
rect 578884 77386 578936 77392
rect 578608 73160 578660 73166
rect 578606 73128 578608 73137
rect 578660 73128 578662 73137
rect 578606 73063 578662 73072
rect 578516 62076 578568 62082
rect 578516 62018 578568 62024
rect 578528 61849 578556 62018
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 577504 55208 577556 55214
rect 577504 55150 577556 55156
rect 578896 54398 578924 77386
rect 579080 71369 579108 77710
rect 579252 75608 579304 75614
rect 579250 75576 579252 75585
rect 579304 75576 579306 75585
rect 579250 75511 579306 75520
rect 580460 73166 580488 93094
rect 580644 89758 580672 106286
rect 581644 104916 581696 104922
rect 581644 104858 581696 104864
rect 580632 89752 580684 89758
rect 580632 89694 580684 89700
rect 581656 75614 581684 104858
rect 581840 84046 581868 109686
rect 583036 103358 583064 128318
rect 584416 124166 584444 139402
rect 585796 134298 585824 144910
rect 587360 135930 587388 146270
rect 589200 145586 589228 149223
rect 589370 147656 589426 147665
rect 589370 147591 589426 147600
rect 589384 146334 589412 147591
rect 589372 146328 589424 146334
rect 589372 146270 589424 146276
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589188 145580 589240 145586
rect 589188 145522 589240 145528
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589922 144392 589978 144401
rect 589922 144327 589978 144336
rect 589462 142760 589518 142769
rect 589462 142695 589518 142704
rect 589476 142186 589504 142695
rect 589464 142180 589516 142186
rect 589464 142122 589516 142128
rect 589094 141128 589150 141137
rect 589094 141063 589150 141072
rect 587348 135924 587400 135930
rect 587348 135866 587400 135872
rect 587164 135312 587216 135318
rect 587164 135254 587216 135260
rect 585784 134292 585836 134298
rect 585784 134234 585836 134240
rect 585968 133952 586020 133958
rect 585968 133894 586020 133900
rect 585784 124228 585836 124234
rect 585784 124170 585836 124176
rect 584404 124160 584456 124166
rect 584404 124102 584456 124108
rect 584404 121508 584456 121514
rect 584404 121450 584456 121456
rect 583024 103352 583076 103358
rect 583024 103294 583076 103300
rect 582380 102808 582432 102814
rect 582380 102750 582432 102756
rect 582392 95062 582420 102750
rect 584416 97510 584444 121450
rect 585140 115388 585192 115394
rect 585140 115330 585192 115336
rect 585152 108390 585180 115330
rect 585140 108384 585192 108390
rect 585140 108326 585192 108332
rect 585796 99210 585824 124170
rect 585980 116958 586008 133894
rect 587176 118658 587204 135254
rect 589108 133210 589136 141063
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589278 136232 589334 136241
rect 589278 136167 589334 136176
rect 589292 135318 589320 136167
rect 589280 135312 589332 135318
rect 589280 135254 589332 135260
rect 589462 134600 589518 134609
rect 589462 134535 589518 134544
rect 589476 133958 589504 134535
rect 589464 133952 589516 133958
rect 589464 133894 589516 133900
rect 589096 133204 589148 133210
rect 589096 133146 589148 133152
rect 588542 132968 588598 132977
rect 588542 132903 588598 132912
rect 587164 118652 587216 118658
rect 587164 118594 587216 118600
rect 585968 116952 586020 116958
rect 585968 116894 586020 116900
rect 587808 116000 587860 116006
rect 587808 115942 587860 115948
rect 587820 115258 587848 115942
rect 587808 115252 587860 115258
rect 587808 115194 587860 115200
rect 587164 114572 587216 114578
rect 587164 114514 587216 114520
rect 585968 100768 586020 100774
rect 585968 100710 586020 100716
rect 585784 99204 585836 99210
rect 585784 99146 585836 99152
rect 584404 97504 584456 97510
rect 584404 97446 584456 97452
rect 583024 96076 583076 96082
rect 583024 96018 583076 96024
rect 582380 95056 582432 95062
rect 582380 94998 582432 95004
rect 581828 84040 581880 84046
rect 581828 83982 581880 83988
rect 581644 75608 581696 75614
rect 581644 75550 581696 75556
rect 580448 73160 580500 73166
rect 580448 73102 580500 73108
rect 579066 71360 579122 71369
rect 579066 71295 579122 71304
rect 579526 68096 579582 68105
rect 579526 68031 579582 68040
rect 579540 67658 579568 68031
rect 579528 67652 579580 67658
rect 579528 67594 579580 67600
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 581644 65544 581696 65550
rect 581644 65486 581696 65492
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 580264 62824 580316 62830
rect 580264 62766 580316 62772
rect 579528 60716 579580 60722
rect 579528 60658 579580 60664
rect 579540 60353 579568 60658
rect 579526 60344 579582 60353
rect 579526 60279 579582 60288
rect 579068 58676 579120 58682
rect 579068 58618 579120 58624
rect 578884 54392 578936 54398
rect 578884 54334 578936 54340
rect 579080 54262 579108 58618
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 579528 56568 579580 56574
rect 579528 56510 579580 56516
rect 579540 56137 579568 56510
rect 579526 56128 579582 56137
rect 579526 56063 579582 56072
rect 579068 54256 579120 54262
rect 580276 54233 580304 62766
rect 581656 55049 581684 65486
rect 581642 55040 581698 55049
rect 581642 54975 581698 54984
rect 583036 54942 583064 96018
rect 584404 94512 584456 94518
rect 584404 94454 584456 94460
rect 583024 54936 583076 54942
rect 583024 54878 583076 54884
rect 584416 54777 584444 94454
rect 585980 80102 586008 100710
rect 587176 88330 587204 114514
rect 588556 113150 588584 132903
rect 589936 131782 589964 144327
rect 589924 131776 589976 131782
rect 589924 131718 589976 131724
rect 590106 131336 590162 131345
rect 590106 131271 590162 131280
rect 589462 129704 589518 129713
rect 589462 129639 589518 129648
rect 589476 128382 589504 129639
rect 589464 128376 589516 128382
rect 589464 128318 589516 128324
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589462 124808 589518 124817
rect 589462 124743 589518 124752
rect 589476 124234 589504 124743
rect 589464 124228 589516 124234
rect 589464 124170 589516 124176
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589462 121544 589518 121553
rect 589462 121479 589464 121488
rect 589516 121479 589518 121488
rect 589464 121450 589516 121456
rect 590120 120766 590148 131271
rect 590290 126440 590346 126449
rect 590290 126375 590346 126384
rect 590108 120760 590160 120766
rect 590108 120702 590160 120708
rect 589922 119912 589978 119921
rect 589922 119847 589978 119856
rect 588726 118280 588782 118289
rect 588726 118215 588782 118224
rect 588544 113144 588596 113150
rect 588544 113086 588596 113092
rect 588544 110492 588596 110498
rect 588544 110434 588596 110440
rect 587164 88324 587216 88330
rect 587164 88266 587216 88272
rect 588556 82822 588584 110434
rect 588740 93838 588768 118215
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589646 115016 589702 115025
rect 589646 114951 589702 114960
rect 589660 114578 589688 114951
rect 589648 114572 589700 114578
rect 589648 114514 589700 114520
rect 589554 113384 589610 113393
rect 589554 113319 589610 113328
rect 589568 113174 589596 113319
rect 589568 113146 589688 113174
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589278 110120 589334 110129
rect 589278 110055 589334 110064
rect 589292 106962 589320 110055
rect 589476 109750 589504 111687
rect 589660 110498 589688 113146
rect 589648 110492 589700 110498
rect 589648 110434 589700 110440
rect 589464 109744 589516 109750
rect 589464 109686 589516 109692
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589280 106956 589332 106962
rect 589280 106898 589332 106904
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589936 102814 589964 119847
rect 590304 115394 590332 126375
rect 590292 115388 590344 115394
rect 590292 115330 590344 115336
rect 591316 114442 591344 208626
rect 666204 186969 666232 338098
rect 667216 313721 667244 456758
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667388 350600 667440 350606
rect 667388 350542 667440 350548
rect 667202 313712 667258 313721
rect 667202 313647 667258 313656
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 666836 226500 666888 226506
rect 666836 226442 666888 226448
rect 666848 223145 666876 226442
rect 667020 226092 667072 226098
rect 667020 226034 667072 226040
rect 667032 223417 667060 226034
rect 667018 223408 667074 223417
rect 667018 223343 667074 223352
rect 666834 223136 666890 223145
rect 666834 223071 666890 223080
rect 667018 222184 667074 222193
rect 667018 222119 667074 222128
rect 666834 219464 666890 219473
rect 666834 219399 666890 219408
rect 666466 215384 666522 215393
rect 666466 215319 666522 215328
rect 666480 200977 666508 215319
rect 666466 200968 666522 200977
rect 666466 200903 666522 200912
rect 666190 186960 666246 186969
rect 666190 186895 666246 186904
rect 666848 174865 666876 219399
rect 667032 214577 667060 222119
rect 667018 214568 667074 214577
rect 667018 214503 667074 214512
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 174856 666890 174865
rect 666834 174791 666890 174800
rect 667032 133113 667060 209034
rect 667216 134609 667244 310490
rect 667400 181393 667428 350542
rect 667756 324352 667808 324358
rect 667756 324294 667808 324300
rect 667572 284368 667624 284374
rect 667572 284310 667624 284316
rect 667386 181384 667442 181393
rect 667386 181319 667442 181328
rect 667584 135969 667612 284310
rect 667768 178809 667796 324294
rect 668596 312905 668624 444382
rect 668780 360913 668808 484366
rect 669056 483177 669084 558991
rect 669042 483168 669098 483177
rect 669042 483103 669098 483112
rect 669240 456249 669268 705055
rect 669424 663649 669452 741095
rect 669608 709617 669636 789375
rect 669792 750961 669820 864175
rect 669964 815652 670016 815658
rect 669964 815594 670016 815600
rect 669778 750952 669834 750961
rect 669778 750887 669834 750896
rect 669778 738576 669834 738585
rect 669778 738511 669834 738520
rect 669594 709608 669650 709617
rect 669594 709543 669650 709552
rect 669594 695192 669650 695201
rect 669594 695127 669650 695136
rect 669410 663640 669466 663649
rect 669410 663575 669466 663584
rect 669608 620673 669636 695127
rect 669792 666233 669820 738511
rect 669976 673169 670004 815594
rect 670330 783048 670386 783057
rect 670330 782983 670386 782992
rect 670146 780600 670202 780609
rect 670146 780535 670202 780544
rect 670160 710433 670188 780535
rect 670146 710424 670202 710433
rect 670146 710359 670202 710368
rect 670344 707577 670372 782983
rect 670620 751777 670648 867847
rect 670974 781144 671030 781153
rect 670974 781079 671030 781088
rect 670606 751768 670662 751777
rect 670606 751703 670662 751712
rect 670790 750136 670846 750145
rect 670790 750071 670846 750080
rect 670804 727977 670832 750071
rect 670988 736934 671016 781079
rect 671172 752593 671200 872199
rect 671356 763065 671384 895630
rect 671342 763056 671398 763065
rect 671342 762991 671398 763000
rect 671632 758554 671660 935711
rect 671816 758713 671844 936663
rect 672644 930134 672672 937479
rect 672828 930134 672856 937751
rect 673012 930617 673040 958695
rect 673196 934697 673224 962503
rect 673182 934688 673238 934697
rect 673182 934623 673238 934632
rect 673380 932657 673408 962775
rect 674194 957128 674250 957137
rect 674194 957063 674250 957072
rect 673366 932648 673422 932657
rect 673366 932583 673422 932592
rect 672998 930608 673054 930617
rect 672998 930543 673054 930552
rect 674208 930209 674236 957063
rect 674392 933065 674420 966039
rect 675036 963254 675064 966709
rect 675206 966104 675262 966113
rect 675262 966062 675418 966090
rect 675206 966039 675262 966048
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675206 963656 675262 963665
rect 675206 963591 675262 963600
rect 675220 963254 675248 963591
rect 675404 963393 675432 963595
rect 675390 963384 675446 963393
rect 675390 963319 675446 963328
rect 674944 963226 675064 963254
rect 675128 963226 675248 963254
rect 674944 962577 674972 963226
rect 674930 962568 674986 962577
rect 674930 962503 674986 962512
rect 674654 962160 674710 962169
rect 674654 962095 674710 962104
rect 674378 933056 674434 933065
rect 674378 932991 674434 933000
rect 674668 932249 674696 962095
rect 675128 961769 675156 963226
rect 675496 962849 675524 963016
rect 675482 962840 675538 962849
rect 675482 962775 675538 962784
rect 675404 962169 675432 962404
rect 675390 962160 675446 962169
rect 675390 962095 675446 962104
rect 675128 961741 675418 961769
rect 675206 959304 675262 959313
rect 675262 959262 675418 959290
rect 675206 959239 675262 959248
rect 675114 958760 675170 958769
rect 675170 958718 675418 958746
rect 675114 958695 675170 958704
rect 675772 957817 675800 958052
rect 675298 957808 675354 957817
rect 675298 957743 675354 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 675312 955482 675340 957743
rect 675496 957137 675524 957440
rect 675482 957128 675538 957137
rect 675482 957063 675538 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675022 954544 675078 954553
rect 675022 954479 675078 954488
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 932240 674710 932249
rect 674654 932175 674710 932184
rect 674194 930200 674250 930209
rect 674194 930135 674250 930144
rect 672184 930106 672672 930134
rect 672736 930106 672856 930134
rect 671986 928296 672042 928305
rect 671986 928231 672042 928240
rect 671802 758704 671858 758713
rect 671802 758639 671858 758648
rect 671632 758526 671752 758554
rect 671526 758296 671582 758305
rect 671526 758231 671582 758240
rect 671158 752584 671214 752593
rect 671158 752519 671214 752528
rect 671158 737080 671214 737089
rect 671158 737015 671214 737024
rect 670896 736906 671016 736934
rect 670896 728090 670924 736906
rect 671172 734210 671200 737015
rect 671344 735616 671396 735622
rect 671344 735558 671396 735564
rect 671172 734182 671292 734210
rect 671066 730552 671122 730561
rect 671066 730487 671122 730496
rect 670896 728062 671016 728090
rect 670790 727968 670846 727977
rect 670790 727903 670846 727912
rect 670988 727274 671016 728062
rect 670896 727246 671016 727274
rect 670896 721834 670924 727246
rect 670896 721806 671016 721834
rect 670790 712464 670846 712473
rect 670790 712399 670846 712408
rect 670330 707568 670386 707577
rect 670330 707503 670386 707512
rect 670606 699816 670662 699825
rect 670606 699751 670662 699760
rect 670330 687440 670386 687449
rect 670330 687375 670386 687384
rect 669962 673160 670018 673169
rect 669962 673095 670018 673104
rect 669778 666224 669834 666233
rect 669778 666159 669834 666168
rect 670148 656940 670200 656946
rect 670148 656882 670200 656888
rect 669778 645416 669834 645425
rect 669778 645351 669834 645360
rect 669594 620664 669650 620673
rect 669594 620599 669650 620608
rect 669792 574977 669820 645351
rect 669962 644872 670018 644881
rect 669962 644807 670018 644816
rect 669778 574968 669834 574977
rect 669778 574903 669834 574912
rect 669976 571577 670004 644807
rect 669962 571568 670018 571577
rect 669962 571503 670018 571512
rect 669410 570344 669466 570353
rect 669410 570279 669466 570288
rect 669424 500993 669452 570279
rect 669778 556200 669834 556209
rect 669778 556135 669834 556144
rect 669594 553480 669650 553489
rect 669594 553415 669650 553424
rect 669410 500984 669466 500993
rect 669410 500919 669466 500928
rect 669608 482361 669636 553415
rect 669792 483585 669820 556135
rect 670160 537849 670188 656882
rect 670344 621014 670372 687375
rect 670620 621014 670648 699751
rect 670804 667729 670832 712399
rect 670988 706761 671016 721806
rect 671080 721754 671108 730487
rect 671080 721726 671200 721754
rect 670974 706752 671030 706761
rect 670974 706687 671030 706696
rect 670974 685536 671030 685545
rect 670974 685471 671030 685480
rect 670790 667720 670846 667729
rect 670790 667655 670846 667664
rect 670988 666482 671016 685471
rect 670896 666454 671016 666482
rect 670896 661858 670924 666454
rect 671172 666346 671200 721726
rect 671080 666318 671200 666346
rect 671080 666262 671108 666318
rect 671068 666256 671120 666262
rect 671068 666198 671120 666204
rect 671264 666074 671292 734182
rect 671172 666046 671292 666074
rect 671172 662425 671200 666046
rect 671158 662416 671214 662425
rect 671158 662351 671214 662360
rect 670896 661830 671016 661858
rect 670790 623928 670846 623937
rect 670790 623863 670846 623872
rect 670252 620986 670372 621014
rect 670436 620986 670648 621014
rect 670252 619290 670280 620986
rect 670436 619449 670464 620986
rect 670422 619440 670478 619449
rect 670422 619375 670478 619384
rect 670252 619262 670464 619290
rect 670436 618225 670464 619262
rect 670422 618216 670478 618225
rect 670422 618151 670478 618160
rect 670606 607336 670662 607345
rect 670606 607271 670662 607280
rect 670330 598904 670386 598913
rect 670330 598839 670386 598848
rect 670146 537840 670202 537849
rect 670146 537775 670202 537784
rect 669964 536852 670016 536858
rect 669964 536794 670016 536800
rect 669778 483576 669834 483585
rect 669778 483511 669834 483520
rect 669594 482352 669650 482361
rect 669594 482287 669650 482296
rect 669226 456240 669282 456249
rect 669226 456175 669282 456184
rect 669976 403753 670004 536794
rect 670344 528193 670372 598839
rect 670620 529689 670648 607271
rect 670804 579057 670832 623863
rect 670988 619857 671016 661830
rect 671158 640520 671214 640529
rect 671158 640455 671214 640464
rect 670974 619848 671030 619857
rect 670974 619783 671030 619792
rect 671172 596174 671200 640455
rect 671356 627881 671384 735558
rect 671540 713697 671568 758231
rect 671724 757897 671752 758526
rect 671710 757888 671766 757897
rect 671710 757823 671766 757832
rect 671710 757480 671766 757489
rect 671710 757415 671766 757424
rect 671526 713688 671582 713697
rect 671526 713623 671582 713632
rect 671526 713280 671582 713289
rect 671526 713215 671582 713224
rect 671540 712094 671568 713215
rect 671724 712881 671752 757415
rect 672000 732873 672028 928231
rect 672184 770681 672212 930106
rect 672538 873624 672594 873633
rect 672538 873559 672594 873568
rect 672354 784408 672410 784417
rect 672354 784343 672410 784352
rect 672170 770672 672226 770681
rect 672170 770607 672226 770616
rect 672170 733952 672226 733961
rect 672170 733887 672226 733896
rect 671986 732864 672042 732873
rect 671986 732799 672042 732808
rect 671710 712872 671766 712881
rect 671710 712807 671766 712816
rect 671540 712066 671660 712094
rect 671632 668545 671660 712066
rect 671986 688664 672042 688673
rect 671986 688599 672042 688608
rect 671618 668536 671674 668545
rect 671618 668471 671674 668480
rect 671802 668128 671858 668137
rect 671802 668063 671858 668072
rect 671526 667312 671582 667321
rect 671526 667247 671582 667256
rect 671540 649994 671568 667247
rect 671540 649966 671660 649994
rect 671342 627872 671398 627881
rect 671342 627807 671398 627816
rect 671632 626634 671660 649966
rect 671448 626606 671660 626634
rect 671448 622713 671476 626606
rect 671618 624472 671674 624481
rect 671618 624407 671674 624416
rect 671632 623234 671660 624407
rect 671816 623529 671844 668063
rect 671802 623520 671858 623529
rect 671802 623455 671858 623464
rect 671632 623206 671936 623234
rect 671710 623112 671766 623121
rect 671710 623047 671766 623056
rect 671434 622704 671490 622713
rect 671434 622639 671490 622648
rect 671436 612196 671488 612202
rect 671436 612138 671488 612144
rect 671080 596146 671200 596174
rect 670790 579048 670846 579057
rect 670790 578983 670846 578992
rect 670790 578640 670846 578649
rect 670790 578575 670846 578584
rect 670804 571962 670832 578575
rect 671080 578066 671108 596146
rect 671250 594824 671306 594833
rect 671250 594759 671306 594768
rect 671068 578060 671120 578066
rect 671068 578002 671120 578008
rect 671066 577824 671122 577833
rect 671066 577759 671122 577768
rect 671080 572714 671108 577759
rect 671080 572686 671200 572714
rect 670804 571934 671016 571962
rect 670790 569528 670846 569537
rect 670790 569463 670846 569472
rect 670804 567194 670832 569463
rect 670804 567166 670924 567194
rect 670896 538214 670924 567166
rect 670804 538186 670924 538214
rect 670804 534074 670832 538186
rect 670988 535129 671016 571934
rect 671172 567194 671200 572686
rect 671080 567166 671200 567194
rect 671080 557534 671108 567166
rect 671080 557506 671200 557534
rect 670974 535120 671030 535129
rect 670974 535055 671030 535064
rect 671172 534970 671200 557506
rect 671080 534942 671200 534970
rect 670804 534046 670924 534074
rect 670606 529680 670662 529689
rect 670606 529615 670662 529624
rect 670330 528184 670386 528193
rect 670330 528119 670386 528128
rect 670896 455161 670924 534046
rect 671080 533497 671108 534942
rect 671066 533488 671122 533497
rect 671066 533423 671122 533432
rect 671066 532944 671122 532953
rect 671066 532879 671122 532888
rect 671080 489297 671108 532879
rect 671264 525745 671292 594759
rect 671448 579873 671476 612138
rect 671434 579864 671490 579873
rect 671434 579799 671490 579808
rect 671526 579456 671582 579465
rect 671526 579391 671582 579400
rect 671540 572714 671568 579391
rect 671724 578241 671752 623047
rect 671908 612338 671936 623206
rect 672000 618254 672028 688599
rect 672184 661609 672212 733887
rect 672368 709209 672396 784343
rect 672552 754225 672580 873559
rect 672736 760345 672764 930106
rect 673366 929520 673422 929529
rect 673366 929455 673422 929464
rect 672998 870088 673054 870097
rect 672998 870023 673054 870032
rect 672722 760336 672778 760345
rect 672722 760271 672778 760280
rect 672722 759928 672778 759937
rect 672722 759863 672778 759872
rect 672538 754216 672594 754225
rect 672538 754151 672594 754160
rect 672538 738304 672594 738313
rect 672538 738239 672594 738248
rect 672552 736934 672580 738239
rect 672736 736934 672764 759863
rect 673012 755449 673040 870023
rect 673182 759112 673238 759121
rect 673182 759047 673238 759056
rect 672998 755440 673054 755449
rect 672998 755375 673054 755384
rect 672906 751360 672962 751369
rect 672906 751295 672962 751304
rect 672920 736934 672948 751295
rect 672552 736906 672672 736934
rect 672736 736906 672856 736934
rect 672920 736906 673040 736934
rect 672354 709200 672410 709209
rect 672354 709135 672410 709144
rect 672448 707260 672500 707266
rect 672448 707202 672500 707208
rect 672460 670177 672488 707202
rect 672446 670168 672502 670177
rect 672446 670103 672502 670112
rect 672446 669896 672502 669905
rect 672446 669831 672502 669840
rect 672170 661600 672226 661609
rect 672170 661535 672226 661544
rect 672170 638752 672226 638761
rect 672170 638687 672226 638696
rect 672184 630674 672212 638687
rect 672184 630646 672304 630674
rect 672000 618226 672120 618254
rect 672092 616729 672120 618226
rect 672078 616720 672134 616729
rect 672078 616655 672134 616664
rect 672078 614952 672134 614961
rect 672078 614887 672134 614896
rect 671896 612332 671948 612338
rect 671896 612274 671948 612280
rect 672092 608594 672120 614887
rect 672000 608566 672120 608594
rect 671710 578232 671766 578241
rect 671710 578167 671766 578176
rect 671712 578060 671764 578066
rect 671712 578002 671764 578008
rect 671724 576201 671752 578002
rect 671710 576192 671766 576201
rect 671710 576127 671766 576136
rect 671540 572686 671844 572714
rect 671816 567194 671844 572686
rect 671448 567166 671844 567194
rect 671448 534721 671476 567166
rect 671710 555248 671766 555257
rect 671710 555183 671766 555192
rect 671434 534712 671490 534721
rect 671434 534647 671490 534656
rect 671526 534440 671582 534449
rect 671526 534375 671582 534384
rect 671250 525736 671306 525745
rect 671250 525671 671306 525680
rect 671540 490929 671568 534375
rect 671526 490920 671582 490929
rect 671526 490855 671582 490864
rect 671066 489288 671122 489297
rect 671066 489223 671122 489232
rect 671724 486033 671752 555183
rect 671710 486024 671766 486033
rect 671710 485959 671766 485968
rect 672000 455433 672028 608566
rect 672276 601694 672304 630646
rect 672460 625161 672488 669831
rect 672644 662425 672672 736906
rect 672828 715329 672856 736906
rect 673012 728142 673040 736906
rect 673000 728136 673052 728142
rect 673000 728078 673052 728084
rect 672814 715320 672870 715329
rect 672814 715255 672870 715264
rect 672814 714912 672870 714921
rect 672814 714847 672870 714856
rect 672828 669497 672856 714847
rect 673196 714513 673224 759047
rect 673380 732873 673408 929455
rect 674852 928792 674880 953391
rect 675036 934289 675064 954479
rect 675220 954366 675418 954394
rect 675220 951425 675248 954366
rect 675404 953465 675432 953768
rect 675390 953456 675446 953465
rect 675390 953391 675446 953400
rect 675312 952530 675418 952558
rect 675312 951810 675340 952530
rect 675312 951782 675524 951810
rect 675496 951538 675524 951782
rect 677506 951552 677562 951561
rect 675496 951510 676076 951538
rect 675206 951416 675262 951425
rect 675206 951351 675262 951360
rect 675850 951416 675906 951425
rect 675850 951351 675906 951360
rect 675206 951144 675262 951153
rect 675206 951079 675262 951088
rect 675022 934280 675078 934289
rect 675022 934215 675078 934224
rect 675220 933881 675248 951079
rect 675864 949482 675892 951351
rect 675852 949476 675904 949482
rect 675852 949418 675904 949424
rect 676048 948054 676076 951510
rect 677506 951487 677562 951496
rect 676036 948048 676088 948054
rect 676036 947990 676088 947996
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676494 938088 676550 938097
rect 676048 938046 676494 938074
rect 676048 937825 676076 938046
rect 676494 938023 676550 938032
rect 676034 937816 676090 937825
rect 676034 937751 676090 937760
rect 675206 933872 675262 933881
rect 675206 933807 675262 933816
rect 677520 931161 677548 951487
rect 678242 950736 678298 950745
rect 678242 950671 678298 950680
rect 678256 935649 678284 950671
rect 682384 949476 682436 949482
rect 682384 949418 682436 949424
rect 681004 948048 681056 948054
rect 681004 947990 681056 947996
rect 678242 935640 678298 935649
rect 678242 935575 678298 935584
rect 681016 933609 681044 947990
rect 682396 935241 682424 949418
rect 683118 947336 683174 947345
rect 683118 947271 683174 947280
rect 683132 939729 683160 947271
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683118 939720 683174 939729
rect 683118 939655 683174 939664
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 681002 933600 681058 933609
rect 681002 933535 681058 933544
rect 677506 931152 677562 931161
rect 677506 931087 677562 931096
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 675298 879200 675354 879209
rect 675298 879135 675354 879144
rect 675312 877418 675340 879135
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675312 876982 675432 877010
rect 675312 876874 675340 876982
rect 674944 876846 675340 876874
rect 675404 876860 675432 876982
rect 674944 870913 674972 876846
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675404 873633 675432 873868
rect 675390 873624 675446 873633
rect 675390 873559 675446 873568
rect 675114 873216 675170 873225
rect 675170 873174 675418 873202
rect 675114 873151 675170 873160
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 674930 870904 674986 870913
rect 674930 870839 674986 870848
rect 675114 870088 675170 870097
rect 675170 870046 675418 870074
rect 675114 870023 675170 870032
rect 674116 869502 675418 869530
rect 673918 864920 673974 864929
rect 673918 864855 673974 864864
rect 673734 779240 673790 779249
rect 673734 779175 673790 779184
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673366 732864 673422 732873
rect 673366 732799 673422 732808
rect 673564 732154 673592 777407
rect 673748 756254 673776 779175
rect 673932 772041 673960 864855
rect 673918 772032 673974 772041
rect 673918 771967 673974 771976
rect 674116 756254 674144 869502
rect 674668 868861 675340 868889
rect 674470 788080 674526 788089
rect 674470 788015 674526 788024
rect 674286 779920 674342 779929
rect 674286 779855 674342 779864
rect 673656 756226 673776 756254
rect 673932 756226 674144 756254
rect 673656 736930 673684 756226
rect 673932 752185 673960 756226
rect 673918 752176 673974 752185
rect 673918 752111 673974 752120
rect 673656 736902 673776 736930
rect 673552 732148 673604 732154
rect 673552 732090 673604 732096
rect 673366 730144 673422 730153
rect 673366 730079 673422 730088
rect 673380 728634 673408 730079
rect 673748 728770 673776 736902
rect 674012 732148 674064 732154
rect 674012 732090 674064 732096
rect 673656 728742 673776 728770
rect 673380 728606 673592 728634
rect 673366 728512 673422 728521
rect 673366 728447 673368 728456
rect 673420 728447 673422 728456
rect 673368 728418 673420 728424
rect 673564 728362 673592 728606
rect 673380 728334 673592 728362
rect 673182 714504 673238 714513
rect 673182 714439 673238 714448
rect 672998 714096 673054 714105
rect 672998 714031 673054 714040
rect 673012 707266 673040 714031
rect 673000 707260 673052 707266
rect 673000 707202 673052 707208
rect 673182 698320 673238 698329
rect 673182 698255 673238 698264
rect 672998 685808 673054 685817
rect 672998 685743 673054 685752
rect 672814 669488 672870 669497
rect 672814 669423 672870 669432
rect 672814 668944 672870 668953
rect 672814 668879 672870 668888
rect 672630 662416 672686 662425
rect 672630 662351 672686 662360
rect 672630 661192 672686 661201
rect 672630 661127 672686 661136
rect 672446 625152 672502 625161
rect 672446 625087 672502 625096
rect 672446 604344 672502 604353
rect 672446 604279 672502 604288
rect 672184 601666 672304 601694
rect 672184 574569 672212 601666
rect 672170 574560 672226 574569
rect 672170 574495 672226 574504
rect 672264 572008 672316 572014
rect 672264 571950 672316 571956
rect 672276 532681 672304 571950
rect 672262 532672 672318 532681
rect 672262 532607 672318 532616
rect 672264 532024 672316 532030
rect 672264 531966 672316 531972
rect 672276 524414 672304 531966
rect 672460 529009 672488 604279
rect 672644 546281 672672 661127
rect 672828 635497 672856 668879
rect 672814 635488 672870 635497
rect 672814 635423 672870 635432
rect 672814 622296 672870 622305
rect 672814 622231 672870 622240
rect 672828 577425 672856 622231
rect 673012 615777 673040 685743
rect 673196 620945 673224 698255
rect 673380 666505 673408 728334
rect 673656 727274 673684 728742
rect 673828 728612 673880 728618
rect 673828 728554 673880 728560
rect 673840 728249 673868 728554
rect 673826 728240 673882 728249
rect 673826 728175 673882 728184
rect 673826 727696 673882 727705
rect 673826 727631 673882 727640
rect 673840 727274 673868 727631
rect 673564 727246 673684 727274
rect 673748 727246 673868 727274
rect 673564 724169 673592 727246
rect 673748 725778 673776 727246
rect 674024 726617 674052 732090
rect 674150 728136 674202 728142
rect 674150 728078 674202 728084
rect 674162 727977 674190 728078
rect 674148 727968 674204 727977
rect 674148 727903 674204 727912
rect 674300 726889 674328 779855
rect 674484 736934 674512 788015
rect 674668 757217 674696 868861
rect 675312 868850 675340 868861
rect 675404 868850 675432 868875
rect 675312 868822 675432 868850
rect 675298 868456 675354 868465
rect 675298 868391 675354 868400
rect 674838 868184 674894 868193
rect 674838 868119 674894 868128
rect 674852 867513 674880 868119
rect 674838 867504 674894 867513
rect 674838 867439 674894 867448
rect 675312 866266 675340 868391
rect 675496 867921 675524 868224
rect 675482 867912 675538 867921
rect 675482 867847 675538 867856
rect 675482 867504 675538 867513
rect 675482 867439 675538 867448
rect 675496 867035 675524 867439
rect 675312 866238 675432 866266
rect 675404 865844 675432 866238
rect 675404 864929 675432 865195
rect 675390 864920 675446 864929
rect 675390 864855 675446 864864
rect 675496 864249 675524 864552
rect 675482 864240 675538 864249
rect 675482 864175 675538 864184
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 674930 789440 674986 789449
rect 674930 789375 674986 789384
rect 674944 787545 674972 789375
rect 675128 788066 675156 863314
rect 675298 863152 675354 863161
rect 675298 863087 675354 863096
rect 675312 859754 675340 863087
rect 675220 859726 675340 859754
rect 675220 856994 675248 859726
rect 675220 856966 675340 856994
rect 675036 788038 675156 788066
rect 675036 787794 675064 788038
rect 675036 787766 675156 787794
rect 674930 787536 674986 787545
rect 674930 787471 674986 787480
rect 674838 787264 674894 787273
rect 674838 787199 674894 787208
rect 674852 768233 674880 787199
rect 675128 782474 675156 787766
rect 675312 787386 675340 856966
rect 675496 788089 675524 788324
rect 675482 788080 675538 788089
rect 675482 788015 675538 788024
rect 675496 787545 675524 787679
rect 675482 787536 675538 787545
rect 675482 787471 675538 787480
rect 675220 787358 675340 787386
rect 675220 785346 675248 787358
rect 675390 787264 675446 787273
rect 675390 787199 675446 787208
rect 675404 787032 675432 787199
rect 675482 786720 675538 786729
rect 675312 786678 675482 786706
rect 675312 785754 675340 786678
rect 675482 786655 675538 786664
rect 675312 785726 675432 785754
rect 675220 785318 675340 785346
rect 675312 785234 675340 785318
rect 674944 782446 675156 782474
rect 675220 785206 675340 785234
rect 674944 775574 674972 782446
rect 675220 781266 675248 785206
rect 675404 785196 675432 785726
rect 675496 784417 675524 784652
rect 675482 784408 675538 784417
rect 675482 784343 675538 784352
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 783057 675524 783360
rect 675482 783048 675538 783057
rect 675482 782983 675538 782992
rect 675128 781238 675248 781266
rect 674944 775546 675064 775574
rect 675036 774625 675064 775546
rect 675128 774738 675156 781238
rect 675298 781144 675354 781153
rect 675298 781079 675354 781088
rect 675312 779090 675340 781079
rect 675496 780609 675524 780844
rect 675482 780600 675538 780609
rect 675482 780535 675538 780544
rect 675496 779929 675524 780300
rect 675482 779920 675538 779929
rect 675482 779855 675538 779864
rect 675496 779249 675524 779688
rect 675482 779240 675538 779249
rect 675482 779175 675538 779184
rect 675312 779062 675432 779090
rect 675404 779008 675432 779062
rect 675482 778832 675538 778841
rect 675220 778790 675482 778818
rect 675220 776642 675248 778790
rect 675482 778767 675538 778776
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675220 776614 675418 776642
rect 675574 775704 675630 775713
rect 675574 775639 675630 775648
rect 675588 775574 675616 775639
rect 675772 775577 675800 776016
rect 675496 775546 675616 775574
rect 675758 775568 675814 775577
rect 675496 775336 675524 775546
rect 675758 775503 675814 775512
rect 675128 774710 675340 774738
rect 675022 774616 675078 774625
rect 675022 774551 675078 774560
rect 675114 774344 675170 774353
rect 675114 774279 675170 774288
rect 674838 768224 674894 768233
rect 674838 768159 674894 768168
rect 675128 766601 675156 774279
rect 675312 773922 675340 774710
rect 675220 773894 675340 773922
rect 675220 770794 675248 773894
rect 675404 773809 675432 774180
rect 675390 773800 675446 773809
rect 675390 773735 675446 773744
rect 682382 772712 682438 772721
rect 682382 772647 682438 772656
rect 675220 770766 675616 770794
rect 675114 766592 675170 766601
rect 675114 766527 675170 766536
rect 675588 765914 675616 770766
rect 675588 765886 675892 765914
rect 674654 757208 674710 757217
rect 674654 757143 674710 757152
rect 675864 755857 675892 765886
rect 676034 763056 676090 763065
rect 676034 762991 676090 763000
rect 676048 760753 676076 762991
rect 677046 761968 677102 761977
rect 677046 761903 677102 761912
rect 676770 761832 676826 761841
rect 676770 761767 676826 761776
rect 676034 760744 676090 760753
rect 676034 760679 676090 760688
rect 676034 757208 676090 757217
rect 676034 757143 676036 757152
rect 676088 757143 676090 757152
rect 676036 757114 676088 757120
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 676784 754633 676812 761767
rect 677060 755041 677088 761903
rect 682396 757081 682424 772647
rect 683210 772032 683266 772041
rect 683210 771967 683266 771976
rect 683224 770054 683252 771967
rect 683394 770944 683450 770953
rect 683394 770879 683450 770888
rect 683224 770026 683344 770054
rect 683120 757172 683172 757178
rect 683120 757114 683172 757120
rect 682382 757072 682438 757081
rect 682382 757007 682438 757016
rect 677046 755032 677102 755041
rect 677046 754967 677102 754976
rect 676770 754624 676826 754633
rect 676770 754559 676826 754568
rect 683132 753001 683160 757114
rect 683316 756673 683344 770026
rect 683408 759370 683436 770879
rect 683578 770672 683634 770681
rect 683578 770607 683634 770616
rect 683592 759529 683620 770607
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683578 759520 683634 759529
rect 683578 759455 683634 759464
rect 683408 759342 683528 759370
rect 683302 756664 683358 756673
rect 683302 756599 683358 756608
rect 683500 753817 683528 759342
rect 683486 753808 683542 753817
rect 683486 753743 683542 753752
rect 683118 752992 683174 753001
rect 683118 752927 683174 752936
rect 675128 743294 675418 743322
rect 675128 743209 675156 743294
rect 675114 743200 675170 743209
rect 675114 743135 675170 743144
rect 674930 742792 674986 742801
rect 674930 742727 674986 742736
rect 674944 741418 674972 742727
rect 675404 742529 675432 742696
rect 675390 742520 675446 742529
rect 675390 742455 675446 742464
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 741577 675156 742002
rect 675114 741568 675170 741577
rect 675114 741503 675170 741512
rect 674944 741390 675156 741418
rect 674930 741160 674986 741169
rect 674930 741095 674986 741104
rect 674944 739038 674972 741095
rect 675128 740194 675156 741390
rect 675128 740166 675418 740194
rect 675114 739664 675170 739673
rect 675170 739622 675418 739650
rect 675114 739599 675170 739608
rect 674944 739010 675340 739038
rect 675312 738970 675340 739010
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675022 738576 675078 738585
rect 675022 738511 675078 738520
rect 675036 738154 675064 738511
rect 675206 738372 675262 738381
rect 675262 738330 675418 738358
rect 675206 738307 675262 738316
rect 675036 738126 675340 738154
rect 675114 737080 675170 737089
rect 675114 737015 675170 737024
rect 674484 736906 674604 736934
rect 674286 726880 674342 726889
rect 674286 726815 674342 726824
rect 674576 726617 674604 736906
rect 675128 735333 675156 737015
rect 675312 735842 675340 738126
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675128 735305 675418 735333
rect 674760 734658 675418 734686
rect 674760 727705 674788 734658
rect 674930 734360 674986 734369
rect 674930 734295 674986 734304
rect 674944 731626 674972 734295
rect 675128 734017 675418 734045
rect 675128 733961 675156 734017
rect 675114 733952 675170 733961
rect 675114 733887 675170 733896
rect 675114 733680 675170 733689
rect 675114 733615 675170 733624
rect 675128 732850 675156 733615
rect 675128 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674944 731598 675340 731626
rect 675404 731612 675432 731734
rect 675114 731504 675170 731513
rect 675114 731439 675170 731448
rect 675128 729178 675156 731439
rect 675312 730986 675418 731014
rect 675312 730153 675340 730986
rect 675482 730552 675538 730561
rect 675482 730487 675538 730496
rect 675496 730351 675524 730487
rect 675298 730144 675354 730153
rect 675298 730079 675354 730088
rect 675128 729150 675418 729178
rect 674746 727696 674802 727705
rect 674746 727631 674802 727640
rect 683486 726880 683542 726889
rect 683486 726815 683542 726824
rect 674010 726608 674066 726617
rect 674010 726543 674066 726552
rect 674562 726608 674618 726617
rect 674562 726543 674618 726552
rect 673656 725750 673776 725778
rect 682382 725792 682438 725801
rect 673656 725506 673684 725750
rect 682382 725727 682438 725736
rect 673656 725478 673776 725506
rect 673550 724160 673606 724169
rect 673550 724095 673606 724104
rect 673550 689616 673606 689625
rect 673550 689551 673606 689560
rect 673366 666496 673422 666505
rect 673366 666431 673422 666440
rect 673368 666256 673420 666262
rect 673368 666198 673420 666204
rect 673380 660793 673408 666198
rect 673366 660784 673422 660793
rect 673366 660719 673422 660728
rect 673366 659968 673422 659977
rect 673366 659903 673422 659912
rect 673182 620936 673238 620945
rect 673182 620871 673238 620880
rect 672998 615768 673054 615777
rect 672998 615703 673054 615712
rect 673090 604616 673146 604625
rect 673090 604551 673146 604560
rect 672814 577416 672870 577425
rect 672814 577351 672870 577360
rect 672814 577008 672870 577017
rect 672814 576943 672870 576952
rect 672828 572014 672856 576943
rect 672816 572008 672868 572014
rect 672816 571950 672868 571956
rect 672906 559464 672962 559473
rect 672906 559399 672962 559408
rect 672920 557534 672948 559399
rect 672920 557506 673040 557534
rect 672814 548448 672870 548457
rect 672814 548383 672870 548392
rect 672630 546272 672686 546281
rect 672630 546207 672686 546216
rect 672630 533896 672686 533905
rect 672630 533831 672686 533840
rect 672644 532030 672672 533831
rect 672632 532024 672684 532030
rect 672632 531966 672684 531972
rect 672446 529000 672502 529009
rect 672446 528935 672502 528944
rect 672276 524386 672764 524414
rect 672736 490113 672764 524386
rect 672828 495434 672856 548383
rect 673012 543734 673040 557506
rect 672920 543706 673040 543734
rect 672920 505094 672948 543706
rect 673104 538214 673132 604551
rect 673104 538186 673224 538214
rect 673196 530641 673224 538186
rect 673182 530632 673238 530641
rect 673182 530567 673238 530576
rect 673184 530460 673236 530466
rect 673184 530402 673236 530408
rect 672920 505066 673040 505094
rect 673012 495434 673040 505066
rect 672828 495406 672948 495434
rect 673012 495406 673132 495434
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672446 489696 672502 489705
rect 672446 489631 672502 489640
rect 671986 455424 672042 455433
rect 671986 455359 672042 455368
rect 670882 455152 670938 455161
rect 670882 455087 670938 455096
rect 671986 455152 672042 455161
rect 671986 455087 671988 455096
rect 672040 455087 672042 455096
rect 671988 455058 672040 455064
rect 672264 453960 672316 453966
rect 672264 453902 672316 453908
rect 672276 453801 672304 453902
rect 672262 453792 672318 453801
rect 672262 453727 672318 453736
rect 671344 430636 671396 430642
rect 671344 430578 671396 430584
rect 669962 403744 670018 403753
rect 669962 403679 670018 403688
rect 670606 393544 670662 393553
rect 670606 393479 670662 393488
rect 668766 360904 668822 360913
rect 668766 360839 668822 360848
rect 669962 347304 670018 347313
rect 669962 347239 670018 347248
rect 668582 312896 668638 312905
rect 668582 312831 668638 312840
rect 668306 302288 668362 302297
rect 668306 302223 668362 302232
rect 668320 238754 668348 302223
rect 667952 238726 668348 238754
rect 667952 229809 667980 238726
rect 668768 237380 668820 237386
rect 668768 237322 668820 237328
rect 668582 234560 668638 234569
rect 668582 234495 668638 234504
rect 668308 233232 668360 233238
rect 668308 233174 668360 233180
rect 668122 230888 668178 230897
rect 668122 230823 668124 230832
rect 668176 230823 668178 230832
rect 668124 230794 668176 230800
rect 668124 230240 668176 230246
rect 668124 230182 668176 230188
rect 667938 229800 667994 229809
rect 667938 229735 667994 229744
rect 668136 224954 668164 230182
rect 668320 229106 668348 233174
rect 667952 224926 668164 224954
rect 668228 229078 668348 229106
rect 667952 192545 667980 224926
rect 668228 219434 668256 229078
rect 668400 225480 668452 225486
rect 668400 225422 668452 225428
rect 668412 225049 668440 225422
rect 668398 225040 668454 225049
rect 668398 224975 668454 224984
rect 668400 224664 668452 224670
rect 668400 224606 668452 224612
rect 668412 223689 668440 224606
rect 668398 223680 668454 223689
rect 668398 223615 668454 223624
rect 668398 220416 668454 220425
rect 668398 220351 668454 220360
rect 668412 219881 668440 220351
rect 668398 219872 668454 219881
rect 668398 219807 668454 219816
rect 668400 219700 668452 219706
rect 668400 219642 668452 219648
rect 668412 219434 668440 219642
rect 668596 219434 668624 234495
rect 668136 219406 668256 219434
rect 668320 219406 668440 219434
rect 668504 219406 668624 219434
rect 667938 192536 667994 192545
rect 667938 192471 667994 192480
rect 667940 189304 667992 189310
rect 667938 189272 667940 189281
rect 667992 189272 667994 189281
rect 667938 189207 667994 189216
rect 668136 182753 668164 219406
rect 668122 182744 668178 182753
rect 668122 182679 668178 182688
rect 667754 178800 667810 178809
rect 667754 178735 667810 178744
rect 667940 174616 667992 174622
rect 667938 174584 667940 174593
rect 667992 174584 667994 174593
rect 667938 174519 667994 174528
rect 668032 169720 668084 169726
rect 668030 169688 668032 169697
rect 668084 169688 668086 169697
rect 668030 169623 668086 169632
rect 667940 164824 667992 164830
rect 667938 164792 667940 164801
rect 667992 164792 667994 164801
rect 667938 164727 667994 164736
rect 668320 163169 668348 219406
rect 668306 163160 668362 163169
rect 668306 163095 668362 163104
rect 668504 148481 668532 219406
rect 668780 153377 668808 237322
rect 668950 236736 669006 236745
rect 668950 236671 669006 236680
rect 668964 159905 668992 236671
rect 669780 234592 669832 234598
rect 669780 234534 669832 234540
rect 669596 234252 669648 234258
rect 669596 234194 669648 234200
rect 669136 234116 669188 234122
rect 669136 234058 669188 234064
rect 669148 197441 669176 234058
rect 669410 230888 669466 230897
rect 669410 230823 669412 230832
rect 669464 230823 669466 230832
rect 669412 230794 669464 230800
rect 669320 229220 669372 229226
rect 669320 229162 669372 229168
rect 669332 229094 669360 229162
rect 669240 229066 669360 229094
rect 669240 219722 669268 229066
rect 669412 226636 669464 226642
rect 669412 226578 669464 226584
rect 669424 226409 669452 226578
rect 669410 226400 669466 226409
rect 669410 226335 669466 226344
rect 669410 225720 669466 225729
rect 669410 225655 669466 225664
rect 669424 225078 669452 225655
rect 669412 225072 669464 225078
rect 669412 225014 669464 225020
rect 669412 224868 669464 224874
rect 669412 224810 669464 224816
rect 669424 224754 669452 224810
rect 669424 224726 669544 224754
rect 669240 219706 669360 219722
rect 669240 219700 669372 219706
rect 669240 219694 669320 219700
rect 669320 219642 669372 219648
rect 669516 217002 669544 224726
rect 669424 216974 669544 217002
rect 669424 216481 669452 216974
rect 669410 216472 669466 216481
rect 669410 216407 669466 216416
rect 669410 214160 669466 214169
rect 669410 214095 669466 214104
rect 669424 205634 669452 214095
rect 669424 205606 669544 205634
rect 669320 199096 669372 199102
rect 669318 199064 669320 199073
rect 669372 199064 669374 199073
rect 669318 198999 669374 199008
rect 669516 198914 669544 205606
rect 669424 198886 669544 198914
rect 669134 197432 669190 197441
rect 669134 197367 669190 197376
rect 669424 197169 669452 198886
rect 669410 197160 669466 197169
rect 669410 197095 669466 197104
rect 669226 196072 669282 196081
rect 669226 196007 669282 196016
rect 669240 187649 669268 196007
rect 669412 194200 669464 194206
rect 669410 194168 669412 194177
rect 669464 194168 669466 194177
rect 669410 194103 669466 194112
rect 669608 190454 669636 234194
rect 669424 190426 669636 190454
rect 669226 187640 669282 187649
rect 669226 187575 669282 187584
rect 669226 184376 669282 184385
rect 669424 184362 669452 190426
rect 669282 184334 669452 184362
rect 669226 184311 669282 184320
rect 669792 174622 669820 234534
rect 669780 174616 669832 174622
rect 669780 174558 669832 174564
rect 669778 168192 669834 168201
rect 669778 168127 669834 168136
rect 669134 164248 669190 164257
rect 669134 164183 669190 164192
rect 668950 159896 669006 159905
rect 668950 159831 669006 159840
rect 668766 153368 668822 153377
rect 668766 153303 668822 153312
rect 668766 149152 668822 149161
rect 668766 149087 668822 149096
rect 668490 148472 668546 148481
rect 668490 148407 668546 148416
rect 668492 146056 668544 146062
rect 668492 145998 668544 146004
rect 668504 145217 668532 145998
rect 668490 145208 668546 145217
rect 668490 145143 668546 145152
rect 668032 136332 668084 136338
rect 668032 136274 668084 136280
rect 667570 135960 667626 135969
rect 667570 135895 667626 135904
rect 668044 135425 668072 136274
rect 668030 135416 668086 135425
rect 668030 135351 668086 135360
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 667018 133104 667074 133113
rect 667018 133039 667074 133048
rect 668780 125633 668808 149087
rect 669148 138689 669176 164183
rect 669134 138680 669190 138689
rect 669134 138615 669190 138624
rect 668950 128344 669006 128353
rect 668950 128279 669006 128288
rect 668766 125624 668822 125633
rect 668766 125559 668822 125568
rect 668216 125180 668268 125186
rect 668216 125122 668268 125128
rect 668228 119105 668256 125122
rect 668964 120737 668992 128279
rect 669792 125186 669820 168127
rect 669976 136338 670004 347239
rect 670422 257680 670478 257689
rect 670422 257615 670478 257624
rect 670436 235929 670464 257615
rect 670422 235920 670478 235929
rect 670422 235855 670478 235864
rect 670332 235748 670384 235754
rect 670332 235690 670384 235696
rect 670146 232928 670202 232937
rect 670146 232863 670202 232872
rect 670160 164830 670188 232863
rect 670344 169726 670372 235690
rect 670620 224954 670648 393479
rect 671356 269793 671384 430578
rect 672460 401713 672488 489631
rect 672630 488064 672686 488073
rect 672630 487999 672686 488008
rect 672446 401704 672502 401713
rect 672446 401639 672502 401648
rect 672446 400480 672502 400489
rect 672446 400415 672502 400424
rect 672460 355881 672488 400415
rect 672644 400081 672672 487999
rect 672920 485625 672948 495406
rect 672906 485616 672962 485625
rect 672906 485551 672962 485560
rect 673104 484809 673132 495406
rect 673196 488594 673224 530402
rect 673380 488714 673408 659903
rect 673564 636857 673592 689551
rect 673748 681057 673776 725478
rect 676034 718312 676090 718321
rect 676034 718247 676090 718256
rect 676048 715737 676076 718247
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 682396 711657 682424 725727
rect 683302 724160 683358 724169
rect 683302 724095 683358 724104
rect 682382 711648 682438 711657
rect 682382 711583 682438 711592
rect 683316 707985 683344 724095
rect 683302 707976 683358 707985
rect 683302 707911 683358 707920
rect 683500 707169 683528 726815
rect 683670 726472 683726 726481
rect 683670 726407 683726 726416
rect 683684 711249 683712 726407
rect 683854 725520 683910 725529
rect 683854 725455 683910 725464
rect 683670 711240 683726 711249
rect 683670 711175 683726 711184
rect 683868 708393 683896 725455
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683854 708384 683910 708393
rect 683854 708319 683910 708328
rect 683486 707160 683542 707169
rect 683486 707095 683542 707104
rect 674378 706344 674434 706353
rect 674378 706279 674434 706288
rect 674010 693560 674066 693569
rect 674010 693495 674066 693504
rect 673734 681048 673790 681057
rect 673734 680983 673790 680992
rect 673734 647864 673790 647873
rect 673734 647799 673790 647808
rect 673550 636848 673606 636857
rect 673550 636783 673606 636792
rect 673550 603528 673606 603537
rect 673550 603463 673606 603472
rect 673564 601694 673592 603463
rect 673472 601666 673592 601694
rect 673472 596174 673500 601666
rect 673748 598754 673776 647799
rect 674024 640334 674052 693495
rect 674194 690160 674250 690169
rect 674194 690095 674250 690104
rect 674208 683114 674236 690095
rect 674208 683086 674328 683114
rect 674300 649994 674328 683086
rect 674208 649966 674328 649994
rect 674208 642274 674236 649966
rect 674392 648938 674420 706279
rect 674930 699816 674986 699825
rect 674930 699751 674986 699760
rect 674944 697694 674972 699751
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 674944 697666 675418 697694
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695201 675418 695209
rect 675114 695192 675418 695201
rect 675170 695181 675418 695192
rect 675114 695127 675170 695136
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 675128 693994 675418 694022
rect 675128 693569 675156 693994
rect 675114 693560 675170 693569
rect 675114 693495 675170 693504
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 674668 693314 675340 693342
rect 675404 693328 675432 693382
rect 674668 656894 674696 693314
rect 675114 692880 675170 692889
rect 675114 692815 675170 692824
rect 675128 690894 675156 692815
rect 675128 690866 675418 690894
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675312 689710 675432 689738
rect 675312 689625 675340 689710
rect 675404 689656 675432 689710
rect 675298 689616 675354 689625
rect 675298 689551 675354 689560
rect 675128 689030 675418 689058
rect 674930 688936 674986 688945
rect 674930 688871 674986 688880
rect 674944 687154 674972 688871
rect 675128 688673 675156 689030
rect 675298 688936 675354 688945
rect 675298 688871 675354 688880
rect 675114 688664 675170 688673
rect 675114 688599 675170 688608
rect 674944 687126 675156 687154
rect 674838 686488 674894 686497
rect 674838 686423 674894 686432
rect 674852 683114 674880 686423
rect 675128 685998 675156 687126
rect 675312 687018 675340 688871
rect 675496 687449 675524 687820
rect 675482 687440 675538 687449
rect 675482 687375 675538 687384
rect 675312 686990 675524 687018
rect 675496 686664 675524 686990
rect 675128 685970 675418 685998
rect 675482 685808 675538 685817
rect 675482 685743 675538 685752
rect 675206 685536 675262 685545
rect 675206 685471 675262 685480
rect 675220 684570 675248 685471
rect 675496 685372 675524 685743
rect 675220 684542 675432 684570
rect 675404 684148 675432 684542
rect 674852 683086 675248 683114
rect 674838 670168 674894 670177
rect 674838 670103 674894 670112
rect 674852 669497 674880 670103
rect 674838 669488 674894 669497
rect 674838 669423 674894 669432
rect 674668 656866 674972 656894
rect 674300 648910 674420 648938
rect 674300 647234 674328 648910
rect 674944 648530 674972 656866
rect 675220 649777 675248 683086
rect 683210 682680 683266 682689
rect 683210 682615 683266 682624
rect 676494 673160 676550 673169
rect 676494 673095 676550 673104
rect 676508 671129 676536 673095
rect 676494 671120 676550 671129
rect 676494 671055 676550 671064
rect 676494 666224 676550 666233
rect 676494 666159 676550 666168
rect 676508 665417 676536 666159
rect 676494 665408 676550 665417
rect 676494 665343 676550 665352
rect 683224 664601 683252 682615
rect 683670 682408 683726 682417
rect 683670 682343 683726 682352
rect 683486 681048 683542 681057
rect 683486 680983 683542 680992
rect 683210 664592 683266 664601
rect 683210 664527 683266 664536
rect 683500 662969 683528 680983
rect 683684 667049 683712 682343
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683670 667040 683726 667049
rect 683670 666975 683726 666984
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 675390 654256 675446 654265
rect 675390 654191 675446 654200
rect 675404 654134 675432 654191
rect 675312 654106 675432 654134
rect 675312 653018 675340 654106
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675404 651545 675432 651848
rect 675390 651536 675446 651545
rect 675390 651471 675446 651480
rect 675206 649768 675262 649777
rect 675206 649703 675262 649712
rect 675404 649618 675432 650012
rect 675312 649590 675432 649618
rect 675312 649074 675340 649590
rect 675128 649046 675340 649074
rect 675128 648666 675156 649046
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675496 648689 675524 648788
rect 675482 648680 675538 648689
rect 675128 648638 675248 648666
rect 674944 648502 675064 648530
rect 675036 648258 675064 648502
rect 674944 648230 675064 648258
rect 674944 648190 674972 648230
rect 674760 648162 674972 648190
rect 674760 647850 674788 648162
rect 674668 647822 674788 647850
rect 674470 647592 674526 647601
rect 674470 647527 674526 647536
rect 674484 647234 674512 647527
rect 674300 647206 674420 647234
rect 674484 647206 674604 647234
rect 674392 645153 674420 647206
rect 674378 645144 674434 645153
rect 674378 645079 674434 645088
rect 674208 642246 674420 642274
rect 674194 641744 674250 641753
rect 674194 641679 674250 641688
rect 674208 640334 674236 641679
rect 673932 640306 674052 640334
rect 674116 640306 674236 640334
rect 673932 618633 673960 640306
rect 674116 630674 674144 640306
rect 674116 630646 674236 630674
rect 673918 618624 673974 618633
rect 673918 618559 673974 618568
rect 674010 599176 674066 599185
rect 674010 599111 674066 599120
rect 673564 598726 673776 598754
rect 673564 598346 673592 598726
rect 673826 598496 673882 598505
rect 673826 598431 673882 598440
rect 673564 598318 673776 598346
rect 673472 596146 673684 596174
rect 673656 592034 673684 596146
rect 673564 592006 673684 592034
rect 673564 582374 673592 592006
rect 673748 591161 673776 598318
rect 673840 592034 673868 598431
rect 674024 592034 674052 599111
rect 674208 592929 674236 630646
rect 674392 624889 674420 642246
rect 674576 640334 674604 647206
rect 674484 640306 674604 640334
rect 674668 640334 674696 647822
rect 674838 647592 674894 647601
rect 674838 647527 674894 647536
rect 674852 640801 674880 647527
rect 675022 647320 675078 647329
rect 675022 647255 675078 647264
rect 675036 641186 675064 647255
rect 675220 644065 675248 648638
rect 675482 648615 675538 648624
rect 675496 647873 675524 648176
rect 675482 647864 675538 647873
rect 675482 647799 675538 647808
rect 675496 645425 675524 645660
rect 675482 645416 675538 645425
rect 675482 645351 675538 645360
rect 675404 644881 675432 645116
rect 675390 644872 675446 644881
rect 675390 644807 675446 644816
rect 675772 644337 675800 644475
rect 675758 644328 675814 644337
rect 675758 644263 675814 644272
rect 675206 644056 675262 644065
rect 675206 643991 675262 644000
rect 675206 643784 675262 643793
rect 675206 643719 675262 643728
rect 675220 642649 675248 643719
rect 675496 643521 675524 643824
rect 675482 643512 675538 643521
rect 675482 643447 675538 643456
rect 675128 642621 675248 642649
rect 675312 642621 675418 642649
rect 675128 641458 675156 642621
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675036 641158 675248 641186
rect 674838 640792 674894 640801
rect 674838 640727 674894 640736
rect 674668 640306 674788 640334
rect 674484 630674 674512 640306
rect 674484 630646 674604 630674
rect 674378 624880 674434 624889
rect 674378 624815 674434 624824
rect 674378 606520 674434 606529
rect 674378 606455 674434 606464
rect 674194 592920 674250 592929
rect 674194 592855 674250 592864
rect 673840 592006 673960 592034
rect 674024 592006 674144 592034
rect 673734 591152 673790 591161
rect 673734 591087 673790 591096
rect 673932 582374 673960 592006
rect 674116 582374 674144 592006
rect 673564 582346 673684 582374
rect 673656 538214 673684 582346
rect 673840 582346 673960 582374
rect 674024 582346 674144 582374
rect 673656 538186 673776 538214
rect 673748 534074 673776 538186
rect 673656 534046 673776 534074
rect 673656 528465 673684 534046
rect 673840 532273 673868 582346
rect 674024 545737 674052 582346
rect 674194 552120 674250 552129
rect 674194 552055 674250 552064
rect 674010 545728 674066 545737
rect 674010 545663 674066 545672
rect 674010 535392 674066 535401
rect 674010 535327 674066 535336
rect 674024 534177 674052 535327
rect 674010 534168 674066 534177
rect 674010 534103 674066 534112
rect 673826 532264 673882 532273
rect 673826 532199 673882 532208
rect 673826 531856 673882 531865
rect 673826 531791 673882 531800
rect 673840 530466 673868 531791
rect 673828 530460 673880 530466
rect 673828 530402 673880 530408
rect 673642 528456 673698 528465
rect 673642 528391 673698 528400
rect 673368 488708 673420 488714
rect 673368 488650 673420 488656
rect 673196 488566 673408 488594
rect 673380 488481 673408 488566
rect 673366 488472 673422 488481
rect 673366 488407 673422 488416
rect 673368 488300 673420 488306
rect 673368 488242 673420 488248
rect 673090 484800 673146 484809
rect 673090 484735 673146 484744
rect 673380 455954 673408 488242
rect 674208 483993 674236 552055
rect 674392 547097 674420 606455
rect 674576 592657 674604 630646
rect 674760 617409 674788 640306
rect 675220 640166 675248 641158
rect 675404 640529 675432 640795
rect 675390 640520 675446 640529
rect 675390 640455 675446 640464
rect 674944 640138 675248 640166
rect 674944 631417 674972 640138
rect 675404 639826 675432 640152
rect 675220 639798 675432 639826
rect 674930 631408 674986 631417
rect 674930 631343 674986 631352
rect 674746 617400 674802 617409
rect 674746 617335 674802 617344
rect 674838 603256 674894 603265
rect 674838 603191 674894 603200
rect 674852 601089 674880 603191
rect 675022 601760 675078 601769
rect 675022 601695 675078 601704
rect 674838 601080 674894 601089
rect 674838 601015 674894 601024
rect 675036 600545 675064 601695
rect 675022 600536 675078 600545
rect 675022 600471 675078 600480
rect 675022 599720 675078 599729
rect 675022 599655 675078 599664
rect 674838 598904 674894 598913
rect 674838 598839 674894 598848
rect 674852 598097 674880 598839
rect 674838 598088 674894 598097
rect 674838 598023 674894 598032
rect 675036 596873 675064 599655
rect 675022 596864 675078 596873
rect 675022 596799 675078 596808
rect 675220 596174 675248 639798
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675390 638072 675446 638081
rect 675390 638007 675446 638016
rect 675404 637574 675432 638007
rect 677506 637936 677562 637945
rect 677506 637871 677562 637880
rect 675758 637664 675814 637673
rect 675758 637599 675814 637608
rect 675128 596146 675248 596174
rect 675312 637546 675432 637574
rect 674930 595504 674986 595513
rect 674930 595439 674986 595448
rect 674562 592648 674618 592657
rect 674562 592583 674618 592592
rect 674944 592034 674972 595439
rect 675128 592498 675156 596146
rect 675312 595898 675340 637546
rect 675772 631417 675800 637599
rect 675758 631408 675814 631417
rect 675758 631343 675814 631352
rect 675850 627872 675906 627881
rect 675850 627807 675906 627816
rect 675864 626618 675892 627807
rect 675852 626612 675904 626618
rect 675852 626554 675904 626560
rect 676496 626612 676548 626618
rect 676496 626554 676548 626560
rect 676508 625705 676536 626554
rect 676494 625696 676550 625705
rect 676494 625631 676550 625640
rect 677520 622033 677548 637871
rect 683302 636848 683358 636857
rect 683302 636783 683358 636792
rect 683118 624880 683174 624889
rect 683118 624815 683174 624824
rect 677506 622024 677562 622033
rect 677506 621959 677562 621968
rect 683132 617137 683160 624815
rect 683316 617953 683344 636783
rect 683670 635488 683726 635497
rect 683670 635423 683726 635432
rect 683684 624481 683712 635423
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683670 624472 683726 624481
rect 683670 624407 683726 624416
rect 683302 617944 683358 617953
rect 683302 617879 683358 617888
rect 683118 617128 683174 617137
rect 683118 617063 683174 617072
rect 675496 607753 675524 608124
rect 675482 607744 675538 607753
rect 675482 607679 675538 607688
rect 675496 607345 675524 607479
rect 675482 607336 675538 607345
rect 675482 607271 675538 607280
rect 675496 606529 675524 606832
rect 675482 606520 675538 606529
rect 675482 606455 675538 606464
rect 675496 604625 675524 604996
rect 675482 604616 675538 604625
rect 675482 604551 675538 604560
rect 675496 604353 675524 604452
rect 675482 604344 675538 604353
rect 675482 604279 675538 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675496 602993 675524 603160
rect 675482 602984 675538 602993
rect 675482 602919 675538 602928
rect 675482 601080 675538 601089
rect 675482 601015 675538 601024
rect 675496 600644 675524 601015
rect 675482 600536 675538 600545
rect 675482 600471 675538 600480
rect 675496 600100 675524 600471
rect 675496 599185 675524 599488
rect 675482 599176 675538 599185
rect 675482 599111 675538 599120
rect 675496 598505 675524 598808
rect 675482 598496 675538 598505
rect 675482 598431 675538 598440
rect 675482 598088 675538 598097
rect 675482 598023 675538 598032
rect 675496 597652 675524 598023
rect 675482 596864 675538 596873
rect 675482 596799 675538 596808
rect 675496 596428 675524 596799
rect 675220 595870 675340 595898
rect 675220 592634 675248 595870
rect 675404 595513 675432 595816
rect 675390 595504 675446 595513
rect 675390 595439 675446 595448
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593745 675432 593980
rect 675390 593736 675446 593745
rect 675390 593671 675446 593680
rect 683302 592920 683358 592929
rect 683302 592855 683358 592864
rect 683118 592648 683174 592657
rect 675220 592606 676168 592634
rect 675128 592470 675984 592498
rect 675758 592376 675814 592385
rect 675758 592311 675814 592320
rect 675574 592104 675630 592113
rect 675574 592039 675630 592048
rect 674944 592006 675064 592034
rect 674654 558376 674710 558385
rect 674654 558311 674710 558320
rect 674378 547088 674434 547097
rect 674378 547023 674434 547032
rect 674470 535120 674526 535129
rect 674470 535055 674526 535064
rect 674484 534177 674512 535055
rect 674470 534168 674526 534177
rect 674470 534103 674526 534112
rect 674668 484401 674696 558311
rect 674838 556200 674894 556209
rect 674838 556135 674894 556144
rect 674852 554849 674880 556135
rect 674838 554840 674894 554849
rect 674838 554775 674894 554784
rect 675036 554554 675064 592006
rect 675588 586265 675616 592039
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 675772 576609 675800 592311
rect 675956 591394 675984 592470
rect 675944 591388 675996 591394
rect 675944 591330 675996 591336
rect 676140 591258 676168 592606
rect 683118 592583 683174 592592
rect 679624 591388 679676 591394
rect 679624 591330 679676 591336
rect 676128 591252 676180 591258
rect 676128 591194 676180 591200
rect 676034 582992 676090 583001
rect 676034 582927 676090 582936
rect 676048 580281 676076 582927
rect 676034 580272 676090 580281
rect 676034 580207 676090 580216
rect 675758 576600 675814 576609
rect 675758 576535 675814 576544
rect 679636 571334 679664 591330
rect 682384 591252 682436 591258
rect 682384 591194 682436 591200
rect 682396 575657 682424 591194
rect 682382 575648 682438 575657
rect 682382 575583 682438 575592
rect 683132 574025 683160 592583
rect 683118 574016 683174 574025
rect 683118 573951 683174 573960
rect 683316 573209 683344 592855
rect 683486 591152 683542 591161
rect 683486 591087 683542 591096
rect 683302 573200 683358 573209
rect 683302 573135 683358 573144
rect 683500 572393 683528 591087
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683486 572384 683542 572393
rect 683486 572319 683542 572328
rect 679624 571328 679676 571334
rect 679624 571270 679676 571276
rect 683120 571328 683172 571334
rect 683120 571270 683172 571276
rect 683132 570761 683160 571270
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 675206 564496 675262 564505
rect 675206 564431 675262 564440
rect 675220 562306 675248 564431
rect 675390 563136 675446 563145
rect 675390 563071 675446 563080
rect 675404 562904 675432 563071
rect 675220 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 674852 554526 675064 554554
rect 675128 559762 675340 559790
rect 675404 559776 675432 559830
rect 674852 547641 674880 554526
rect 675128 554418 675156 559762
rect 675298 559464 675354 559473
rect 675298 559399 675354 559408
rect 675312 559246 675340 559399
rect 675312 559218 675418 559246
rect 675298 559056 675354 559065
rect 675298 558991 675354 559000
rect 675312 558906 675340 558991
rect 675220 558878 675340 558906
rect 675220 557954 675248 558878
rect 675404 558385 675432 558620
rect 675390 558376 675446 558385
rect 675390 558311 675446 558320
rect 675220 557926 675418 557954
rect 675298 557560 675354 557569
rect 675298 557495 675354 557504
rect 675312 556186 675340 557495
rect 675220 556158 675340 556186
rect 675220 554933 675248 556158
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675220 554905 675418 554933
rect 675298 554840 675354 554849
rect 675298 554775 675354 554784
rect 675128 554390 675248 554418
rect 675220 554146 675248 554390
rect 675312 554282 675340 554775
rect 675312 554254 675418 554282
rect 675128 554118 675248 554146
rect 675128 550634 675156 554118
rect 675298 554024 675354 554033
rect 675298 553959 675354 553968
rect 675312 553874 675340 553959
rect 675220 553846 675340 553874
rect 675220 551253 675248 553846
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 675220 551225 675418 551253
rect 675758 550760 675814 550769
rect 675758 550695 675814 550704
rect 675128 550606 675340 550634
rect 675114 549672 675170 549681
rect 675114 549607 675170 549616
rect 674838 547632 674894 547641
rect 674838 547567 674894 547576
rect 674838 546000 674894 546009
rect 674838 545935 674894 545944
rect 674852 540974 674880 545935
rect 675128 540974 675156 549607
rect 675312 547584 675340 550606
rect 675772 550596 675800 550695
rect 675496 549681 675524 549951
rect 675482 549672 675538 549681
rect 675482 549607 675538 549616
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675850 547632 675906 547641
rect 675312 547556 675524 547584
rect 675850 547567 675852 547576
rect 675298 546544 675354 546553
rect 675298 546479 675354 546488
rect 675312 542994 675340 546479
rect 674852 540946 674972 540974
rect 674944 503849 674972 540946
rect 675036 540946 675156 540974
rect 675220 542966 675340 542994
rect 675036 538214 675064 540946
rect 675036 538186 675156 538214
rect 674930 503840 674986 503849
rect 674930 503775 674986 503784
rect 675128 503690 675156 538186
rect 675220 503826 675248 542966
rect 675496 524414 675524 547556
rect 675904 547567 675906 547576
rect 678244 547596 678296 547602
rect 675852 547538 675904 547544
rect 678244 547538 678296 547544
rect 676402 546272 676458 546281
rect 676402 546207 676458 546216
rect 676034 537840 676090 537849
rect 676034 537775 676090 537784
rect 676048 535741 676076 537775
rect 676034 535732 676090 535741
rect 676034 535667 676090 535676
rect 675758 529680 675814 529689
rect 675758 529615 675814 529624
rect 675772 529213 675800 529615
rect 675758 529204 675814 529213
rect 675758 529139 675814 529148
rect 675312 524386 675524 524414
rect 675312 511994 675340 524386
rect 675852 518832 675904 518838
rect 675852 518774 675904 518780
rect 675864 511994 675892 518774
rect 675312 511966 675432 511994
rect 675220 503798 675340 503826
rect 675036 503662 675156 503690
rect 675036 503577 675064 503662
rect 675022 503568 675078 503577
rect 675022 503503 675078 503512
rect 675312 503418 675340 503798
rect 675036 503390 675340 503418
rect 675036 503305 675064 503390
rect 675022 503296 675078 503305
rect 675022 503231 675078 503240
rect 675404 502334 675432 511966
rect 675588 511966 675892 511994
rect 675588 502334 675616 511966
rect 675850 503840 675906 503849
rect 675850 503775 675906 503784
rect 675864 503674 675892 503775
rect 675852 503668 675904 503674
rect 675852 503610 675904 503616
rect 676034 503568 676090 503577
rect 676034 503503 676036 503512
rect 676088 503503 676090 503512
rect 676036 503474 676088 503480
rect 676034 503296 676090 503305
rect 676034 503231 676090 503240
rect 675312 502306 675432 502334
rect 675496 502306 675616 502334
rect 675852 502376 675904 502382
rect 675852 502318 675904 502324
rect 674930 500984 674986 500993
rect 674930 500919 674986 500928
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674194 483984 674250 483993
rect 674194 483919 674250 483928
rect 674746 464808 674802 464817
rect 674746 464743 674802 464752
rect 674760 456929 674788 464743
rect 673826 456920 673882 456929
rect 673826 456855 673882 456864
rect 674746 456920 674802 456929
rect 674746 456855 674802 456864
rect 673840 456074 673868 456855
rect 673946 456240 674002 456249
rect 673946 456175 673948 456184
rect 674000 456175 674002 456184
rect 673948 456146 674000 456152
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673380 455926 673500 455954
rect 673472 455870 673500 455926
rect 673460 455864 673512 455870
rect 673460 455806 673512 455812
rect 673596 455696 673652 455705
rect 673596 455631 673598 455640
rect 673650 455631 673652 455640
rect 673598 455602 673650 455608
rect 673504 455424 673560 455433
rect 673504 455359 673506 455368
rect 673558 455359 673560 455368
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673386 455152 673388 455161
rect 673440 455152 673442 455161
rect 673386 455087 673442 455096
rect 674944 454889 674972 500919
rect 675312 486441 675340 502306
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 673162 454880 673218 454889
rect 673162 454815 673164 454824
rect 673216 454815 673218 454824
rect 674930 454880 674986 454889
rect 674930 454815 674986 454824
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 675496 454617 675524 502306
rect 675864 485774 675892 502318
rect 676048 500954 676076 503231
rect 676036 500948 676088 500954
rect 676036 500890 676088 500896
rect 676416 495434 676444 546207
rect 678256 531457 678284 547538
rect 683210 547088 683266 547097
rect 683210 547023 683266 547032
rect 679622 546544 679678 546553
rect 679622 546479 679678 546488
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 679636 531049 679664 546479
rect 683224 531865 683252 547023
rect 683394 545728 683450 545737
rect 683394 545663 683450 545672
rect 683210 531856 683266 531865
rect 683210 531791 683266 531800
rect 679622 531040 679678 531049
rect 679622 530975 679678 530984
rect 683408 527785 683436 545663
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683578 532264 683634 532273
rect 683578 532199 683634 532208
rect 683394 527776 683450 527785
rect 683394 527711 683450 527720
rect 683592 526561 683620 532199
rect 683578 526552 683634 526561
rect 683578 526487 683634 526496
rect 676862 525736 676918 525745
rect 676862 525671 676918 525680
rect 676876 502382 676904 525671
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 677888 518838 677916 524447
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683210 503704 683266 503713
rect 679624 503668 679676 503674
rect 683210 503639 683266 503648
rect 679624 503610 679676 503616
rect 676864 502376 676916 502382
rect 676864 502318 676916 502324
rect 676416 495406 676812 495434
rect 676034 494048 676090 494057
rect 676034 493983 676090 493992
rect 676048 492726 676076 493983
rect 676036 492720 676088 492726
rect 676036 492662 676088 492668
rect 675680 485746 675892 485774
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 675482 454608 675538 454617
rect 675482 454543 675538 454552
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 675680 454345 675708 485746
rect 675850 481944 675906 481953
rect 675850 481879 675906 481888
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 675666 454336 675722 454345
rect 675666 454271 675722 454280
rect 672816 454096 672868 454102
rect 672814 454064 672816 454073
rect 672868 454064 672870 454073
rect 672814 453999 672870 454008
rect 675864 453801 675892 481879
rect 676034 480720 676090 480729
rect 676034 480655 676090 480664
rect 676048 454073 676076 480655
rect 676784 455705 676812 495406
rect 677322 492416 677378 492425
rect 677322 492351 677378 492360
rect 677336 487257 677364 492351
rect 677322 487248 677378 487257
rect 677322 487183 677378 487192
rect 679636 486849 679664 503610
rect 682384 503532 682436 503538
rect 682384 503474 682436 503480
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 681016 487665 681044 500890
rect 681002 487656 681058 487665
rect 681002 487591 681058 487600
rect 679622 486840 679678 486849
rect 679622 486775 679678 486784
rect 682396 481545 682424 503474
rect 683224 482769 683252 503639
rect 683578 494728 683634 494737
rect 683578 494663 683634 494672
rect 683396 492720 683448 492726
rect 683396 492662 683448 492668
rect 683408 491745 683436 492662
rect 683394 491736 683450 491745
rect 683394 491671 683450 491680
rect 683592 491337 683620 494663
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 491328 683634 491337
rect 683578 491263 683634 491272
rect 683210 482760 683266 482769
rect 683210 482695 683266 482704
rect 682382 481536 682438 481545
rect 682382 481471 682438 481480
rect 676770 455696 676826 455705
rect 676770 455631 676826 455640
rect 676034 454064 676090 454073
rect 676034 453999 676090 454008
rect 675850 453792 675906 453801
rect 675850 453727 675906 453736
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 676034 405648 676090 405657
rect 676034 405583 676090 405592
rect 676048 403481 676076 405583
rect 676034 403472 676090 403481
rect 676034 403407 676090 403416
rect 683132 403345 683160 406263
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 674654 402248 674710 402257
rect 674654 402183 674710 402192
rect 674194 401432 674250 401441
rect 674194 401367 674250 401376
rect 672630 400072 672686 400081
rect 672630 400007 672686 400016
rect 673182 398848 673238 398857
rect 673182 398783 673238 398792
rect 672998 397216 673054 397225
rect 672998 397151 673054 397160
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 672644 376281 672672 393887
rect 672814 392592 672870 392601
rect 672814 392527 672870 392536
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672446 355872 672502 355881
rect 672446 355807 672502 355816
rect 672446 355464 672502 355473
rect 672446 355399 672502 355408
rect 672262 351384 672318 351393
rect 672262 351319 672318 351328
rect 671986 348936 672042 348945
rect 671986 348871 672042 348880
rect 672000 332353 672028 348871
rect 672276 335345 672304 351319
rect 672262 335336 672318 335345
rect 672262 335271 672318 335280
rect 671986 332344 672042 332353
rect 671986 332279 672042 332288
rect 672460 310865 672488 355399
rect 672630 348528 672686 348537
rect 672630 348463 672686 348472
rect 672446 310856 672502 310865
rect 672446 310791 672502 310800
rect 671986 302016 672042 302025
rect 671986 301951 672042 301960
rect 671342 269784 671398 269793
rect 671342 269719 671398 269728
rect 671526 264072 671582 264081
rect 671526 264007 671582 264016
rect 671342 262168 671398 262177
rect 671342 262103 671398 262112
rect 671356 244769 671384 262103
rect 671342 244760 671398 244769
rect 671342 244695 671398 244704
rect 671540 238241 671568 264007
rect 671802 258904 671858 258913
rect 671802 258839 671858 258848
rect 671816 241505 671844 258839
rect 671802 241496 671858 241505
rect 671802 241431 671858 241440
rect 671526 238232 671582 238241
rect 671526 238167 671582 238176
rect 671344 237652 671396 237658
rect 671344 237594 671396 237600
rect 671356 234614 671384 237594
rect 671528 237244 671580 237250
rect 671528 237186 671580 237192
rect 671540 237130 671568 237186
rect 671264 234586 671384 234614
rect 671448 237102 671568 237130
rect 670792 233640 670844 233646
rect 670792 233582 670844 233588
rect 670804 233186 670832 233582
rect 671068 233504 671120 233510
rect 671068 233446 671120 233452
rect 670712 233158 670832 233186
rect 670712 225060 670740 233158
rect 670884 233096 670936 233102
rect 670884 233038 670936 233044
rect 670896 231854 670924 233038
rect 670896 231826 671016 231854
rect 670988 228970 671016 231826
rect 670896 228942 671016 228970
rect 670896 225162 670924 228942
rect 671080 227225 671108 233446
rect 671066 227216 671122 227225
rect 671066 227151 671122 227160
rect 671068 227044 671120 227050
rect 671068 226986 671120 226992
rect 671080 226681 671108 226986
rect 671066 226672 671122 226681
rect 671066 226607 671122 226616
rect 671068 226296 671120 226302
rect 671068 226238 671120 226244
rect 671080 225729 671108 226238
rect 671066 225720 671122 225729
rect 671066 225655 671122 225664
rect 671066 225448 671122 225457
rect 671066 225383 671122 225392
rect 671080 225282 671108 225383
rect 671068 225276 671120 225282
rect 671068 225218 671120 225224
rect 670896 225134 671200 225162
rect 670712 225032 671108 225060
rect 670528 224926 670648 224954
rect 670528 215294 670556 224926
rect 670928 224496 670984 224505
rect 670928 224431 670984 224440
rect 670942 224330 670970 224431
rect 670930 224324 670982 224330
rect 670930 224266 670982 224272
rect 670882 224088 670938 224097
rect 670882 224023 670938 224032
rect 670700 223984 670752 223990
rect 670698 223952 670700 223961
rect 670752 223952 670754 223961
rect 670698 223887 670754 223896
rect 670698 220416 670754 220425
rect 670698 220351 670754 220360
rect 670712 219881 670740 220351
rect 670698 219872 670754 219881
rect 670698 219807 670754 219816
rect 670896 215294 670924 224023
rect 671080 215294 671108 225032
rect 670528 215266 670648 215294
rect 670620 211177 670648 215266
rect 670804 215266 670924 215294
rect 670988 215266 671108 215294
rect 670606 211168 670662 211177
rect 670606 211103 670662 211112
rect 670606 210896 670662 210905
rect 670606 210831 670662 210840
rect 670620 190369 670648 210831
rect 670804 199102 670832 215266
rect 670792 199096 670844 199102
rect 670792 199038 670844 199044
rect 670988 194290 671016 215266
rect 670804 194262 671016 194290
rect 670804 194206 670832 194262
rect 670792 194200 670844 194206
rect 670792 194142 670844 194148
rect 671172 190454 671200 225134
rect 671264 224954 671292 234586
rect 671448 224954 671476 237102
rect 671620 237040 671672 237046
rect 671620 236982 671672 236988
rect 671632 234614 671660 236982
rect 671540 234586 671660 234614
rect 671540 225162 671568 234586
rect 671804 230444 671856 230450
rect 671804 230386 671856 230392
rect 671816 229537 671844 230386
rect 671802 229528 671858 229537
rect 671802 229463 671858 229472
rect 671804 228268 671856 228274
rect 671804 228210 671856 228216
rect 671816 226001 671844 228210
rect 672000 226409 672028 301951
rect 672644 263594 672672 348463
rect 672644 263566 672764 263594
rect 672736 260834 672764 263566
rect 672368 260806 672764 260834
rect 672368 251174 672396 260806
rect 672630 257000 672686 257009
rect 672630 256935 672686 256944
rect 672644 251174 672672 256935
rect 672368 251146 672580 251174
rect 672644 251146 672764 251174
rect 672552 249098 672580 251146
rect 672552 249070 672672 249098
rect 672172 237856 672224 237862
rect 672172 237798 672224 237804
rect 672184 234569 672212 237798
rect 672448 235748 672500 235754
rect 672448 235690 672500 235696
rect 672170 234560 672226 234569
rect 672170 234495 672226 234504
rect 672264 234388 672316 234394
rect 672264 234330 672316 234336
rect 672276 231606 672304 234330
rect 672264 231600 672316 231606
rect 672264 231542 672316 231548
rect 672170 231432 672226 231441
rect 672170 231367 672226 231376
rect 672184 228478 672212 231367
rect 672172 228472 672224 228478
rect 672172 228414 672224 228420
rect 672264 227248 672316 227254
rect 672264 227190 672316 227196
rect 672276 227089 672304 227190
rect 672262 227080 672318 227089
rect 672262 227015 672318 227024
rect 672264 226908 672316 226914
rect 672264 226850 672316 226856
rect 672276 226545 672304 226850
rect 672262 226536 672318 226545
rect 672262 226471 672318 226480
rect 671986 226400 672042 226409
rect 671986 226335 672042 226344
rect 671802 225992 671858 226001
rect 671802 225927 671858 225936
rect 671820 225752 671872 225758
rect 671820 225694 671872 225700
rect 671712 225548 671764 225554
rect 671832 225536 671860 225694
rect 671832 225508 672304 225536
rect 671712 225490 671764 225496
rect 671724 225264 671752 225490
rect 671724 225236 671844 225264
rect 671540 225134 671752 225162
rect 671724 224954 671752 225134
rect 671264 224926 671384 224954
rect 671448 224926 671568 224954
rect 670804 190426 671200 190454
rect 670606 190360 670662 190369
rect 670606 190295 670662 190304
rect 670804 189310 670832 190426
rect 670792 189304 670844 189310
rect 670792 189246 670844 189252
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670332 169720 670384 169726
rect 670332 169662 670384 169668
rect 670330 165608 670386 165617
rect 670330 165543 670386 165552
rect 670148 164824 670200 164830
rect 670148 164766 670200 164772
rect 669964 136332 670016 136338
rect 669964 136274 670016 136280
rect 669780 125180 669832 125186
rect 669780 125122 669832 125128
rect 669594 122768 669650 122777
rect 669594 122703 669650 122712
rect 669226 121408 669282 121417
rect 669226 121343 669282 121352
rect 668950 120728 669006 120737
rect 668950 120663 669006 120672
rect 668214 119096 668270 119105
rect 668214 119031 668270 119040
rect 668032 117700 668084 117706
rect 668032 117642 668084 117648
rect 668044 117473 668072 117642
rect 668030 117464 668086 117473
rect 668030 117399 668086 117408
rect 591304 114436 591356 114442
rect 591304 114378 591356 114384
rect 668216 114300 668268 114306
rect 668216 114242 668268 114248
rect 668228 112577 668256 114242
rect 669240 114209 669268 121343
rect 669608 114306 669636 122703
rect 670344 117706 670372 165543
rect 670620 147665 670648 170303
rect 671356 147674 671384 224926
rect 671540 150113 671568 224926
rect 671632 224926 671752 224954
rect 671632 215294 671660 224926
rect 671816 221785 671844 225236
rect 672276 225049 672304 225508
rect 671986 225040 672042 225049
rect 671986 224975 672042 224984
rect 672262 225040 672318 225049
rect 672262 224975 672318 224984
rect 671802 221776 671858 221785
rect 671802 221711 671858 221720
rect 671802 220960 671858 220969
rect 672000 220946 672028 224975
rect 672262 224768 672318 224777
rect 672262 224703 672318 224712
rect 672276 224210 672304 224703
rect 671858 220918 672028 220946
rect 672092 224182 672304 224210
rect 671802 220895 671858 220904
rect 672092 220814 672120 224182
rect 672262 224088 672318 224097
rect 672262 224023 672318 224032
rect 672276 222194 672304 224023
rect 672276 222166 672396 222194
rect 672092 220786 672304 220814
rect 671986 219872 672042 219881
rect 671986 219807 672042 219816
rect 672000 215294 672028 219807
rect 671632 215266 671752 215294
rect 671724 158273 671752 215266
rect 671908 215266 672028 215294
rect 671908 176497 671936 215266
rect 672276 214962 672304 220786
rect 672184 214934 672304 214962
rect 672184 214849 672212 214934
rect 672170 214840 672226 214849
rect 672170 214775 672226 214784
rect 672078 213752 672134 213761
rect 672078 213687 672134 213696
rect 672092 200705 672120 213687
rect 672368 205634 672396 222166
rect 672276 205606 672396 205634
rect 672078 200696 672134 200705
rect 672078 200631 672134 200640
rect 672276 196081 672304 205606
rect 672262 196072 672318 196081
rect 672262 196007 672318 196016
rect 672078 183560 672134 183569
rect 672078 183495 672134 183504
rect 671894 176488 671950 176497
rect 671894 176423 671950 176432
rect 671894 166968 671950 166977
rect 671894 166903 671950 166912
rect 671710 158264 671766 158273
rect 671710 158199 671766 158208
rect 671526 150104 671582 150113
rect 671526 150039 671582 150048
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670988 147646 671384 147674
rect 670988 146146 671016 147646
rect 670804 146118 671016 146146
rect 670804 146062 670832 146118
rect 670792 146056 670844 146062
rect 670792 145998 670844 146004
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670332 117700 670384 117706
rect 670332 117642 670384 117648
rect 669596 114300 669648 114306
rect 669596 114242 669648 114248
rect 669226 114200 669282 114209
rect 669226 114135 669282 114144
rect 671356 113174 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670712 113146 671384 113174
rect 668214 112568 668270 112577
rect 668214 112503 668270 112512
rect 668306 111888 668362 111897
rect 668306 111823 668362 111832
rect 668030 109304 668086 109313
rect 668030 109239 668086 109248
rect 667204 106208 667256 106214
rect 667204 106150 667256 106156
rect 667216 106049 667244 106150
rect 666650 106040 666706 106049
rect 666650 105975 666706 105984
rect 667202 106040 667258 106049
rect 667202 105975 667258 105984
rect 590106 103592 590162 103601
rect 590106 103527 590162 103536
rect 589924 102808 589976 102814
rect 589924 102750 589976 102756
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100774 589504 101895
rect 589464 100768 589516 100774
rect 589464 100710 589516 100716
rect 588728 93832 588780 93838
rect 588728 93774 588780 93780
rect 590120 93158 590148 103527
rect 613272 100150 613608 100178
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596468 100014 597080 100042
rect 595272 99346 595300 100014
rect 595260 99340 595312 99346
rect 595260 99282 595312 99288
rect 595272 93854 595300 99282
rect 595272 93826 595484 93854
rect 590108 93152 590160 93158
rect 590108 93094 590160 93100
rect 588544 82816 588596 82822
rect 588544 82758 588596 82764
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 585968 80096 586020 80102
rect 585968 80038 586020 80044
rect 585782 77888 585838 77897
rect 585782 77823 585838 77832
rect 585796 55078 585824 77823
rect 589924 77308 589976 77314
rect 589924 77250 589976 77256
rect 588544 74860 588596 74866
rect 588544 74802 588596 74808
rect 588556 56574 588584 74802
rect 588544 56568 588596 56574
rect 588544 56510 588596 56516
rect 585784 55072 585836 55078
rect 585784 55014 585836 55020
rect 589936 54806 589964 77250
rect 596192 56030 596220 100014
rect 596468 56166 596496 100014
rect 597802 99770 597830 100028
rect 598216 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 597802 99742 597876 99770
rect 597652 96960 597704 96966
rect 597652 96902 597704 96908
rect 596456 56160 596508 56166
rect 596456 56102 596508 56108
rect 596180 56024 596232 56030
rect 596180 55966 596232 55972
rect 589924 54800 589976 54806
rect 584402 54768 584458 54777
rect 589924 54742 589976 54748
rect 584402 54703 584458 54712
rect 597664 54534 597692 96902
rect 597848 54670 597876 99742
rect 598216 96966 598244 100014
rect 598204 96960 598256 96966
rect 598204 96902 598256 96908
rect 598952 95946 598980 100014
rect 598940 95940 598992 95946
rect 598940 95882 598992 95888
rect 599504 84194 599532 100014
rect 600424 96082 600452 100014
rect 600412 96076 600464 96082
rect 600412 96018 600464 96024
rect 600884 84194 600912 100014
rect 601896 94518 601924 100014
rect 601884 94512 601936 94518
rect 601884 94454 601936 94460
rect 602356 84194 602384 100014
rect 599136 84166 599532 84194
rect 600516 84166 600912 84194
rect 601896 84166 602384 84194
rect 599136 55894 599164 84166
rect 600516 58682 600544 84166
rect 601896 62830 601924 84166
rect 603092 65550 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 607168 100042
rect 607384 100014 607720 100042
rect 608120 100014 608456 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 604426 99742 604500 99770
rect 603080 65544 603132 65550
rect 603080 65486 603132 65492
rect 601884 62824 601936 62830
rect 601884 62766 601936 62772
rect 600504 58676 600556 58682
rect 600504 58618 600556 58624
rect 599124 55888 599176 55894
rect 599124 55830 599176 55836
rect 597836 54664 597888 54670
rect 597836 54606 597888 54612
rect 597652 54528 597704 54534
rect 604472 54505 604500 99742
rect 605484 97986 605512 100014
rect 605472 97980 605524 97986
rect 605472 97922 605524 97928
rect 606220 96762 606248 100014
rect 606484 97980 606536 97986
rect 606484 97922 606536 97928
rect 606208 96756 606260 96762
rect 606208 96698 606260 96704
rect 606496 76566 606524 97922
rect 607140 93854 607168 100014
rect 607692 96082 607720 100014
rect 607680 96076 607732 96082
rect 607680 96018 607732 96024
rect 608428 94518 608456 100014
rect 609164 96354 609192 100014
rect 609152 96348 609204 96354
rect 609152 96290 609204 96296
rect 608416 94512 608468 94518
rect 608416 94454 608468 94460
rect 607140 93826 607260 93854
rect 607232 88330 607260 93826
rect 607220 88324 607272 88330
rect 607220 88266 607272 88272
rect 609900 85542 609928 100014
rect 610636 96218 610664 100014
rect 610624 96212 610676 96218
rect 610624 96154 610676 96160
rect 611280 91050 611308 100014
rect 612108 96898 612136 100014
rect 612660 97306 612688 100014
rect 613384 100020 613436 100026
rect 613384 99962 613436 99968
rect 612648 97300 612700 97306
rect 612648 97242 612700 97248
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 612004 96756 612056 96762
rect 612004 96698 612056 96704
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 612016 76702 612044 96698
rect 612660 77994 612688 96834
rect 612648 77988 612700 77994
rect 612648 77930 612700 77936
rect 612004 76696 612056 76702
rect 612004 76638 612056 76644
rect 606484 76560 606536 76566
rect 606484 76502 606536 76508
rect 605840 66292 605892 66298
rect 605840 66234 605892 66240
rect 605852 58682 605880 66234
rect 613396 64870 613424 99962
rect 613580 95946 613608 100150
rect 615224 100156 615276 100162
rect 615224 100098 615276 100104
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 613994 99742 614068 99770
rect 613568 95940 613620 95946
rect 613568 95882 613620 95888
rect 614040 80850 614068 99742
rect 615052 97578 615080 100014
rect 615040 97572 615092 97578
rect 615040 97514 615092 97520
rect 615236 84194 615264 100098
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620140 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 615788 96966 615816 100014
rect 616144 97572 616196 97578
rect 616144 97514 616196 97520
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 614868 84166 615264 84194
rect 614028 80844 614080 80850
rect 614028 80786 614080 80792
rect 613384 64864 613436 64870
rect 613384 64806 613436 64812
rect 614868 60722 614896 84166
rect 616156 79354 616184 97514
rect 616524 94654 616552 100014
rect 617260 96762 617288 100014
rect 617248 96756 617300 96762
rect 617248 96698 617300 96704
rect 616512 94648 616564 94654
rect 616512 94590 616564 94596
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618904 96960 618956 96966
rect 618904 96902 618956 96908
rect 618168 96756 618220 96762
rect 618168 96698 618220 96704
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96698
rect 617340 91044 617392 91050
rect 617340 90986 617392 90992
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 617352 88194 617380 90986
rect 617340 88188 617392 88194
rect 617340 88130 617392 88136
rect 616144 79348 616196 79354
rect 616144 79290 616196 79296
rect 618916 75206 618944 96902
rect 619560 93838 619588 100014
rect 620112 97170 620140 100014
rect 620284 97300 620336 97306
rect 620284 97242 620336 97248
rect 620100 97164 620152 97170
rect 620100 97106 620152 97112
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 620296 76838 620324 97242
rect 620940 96082 620968 100014
rect 621676 97578 621704 100014
rect 622320 98802 622348 100014
rect 622308 98796 622360 98802
rect 622308 98738 622360 98744
rect 623148 97714 623176 100014
rect 623700 98666 623728 100014
rect 624620 99346 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628236 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 631916 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635504 100042
rect 625034 99742 625108 99770
rect 624608 99340 624660 99346
rect 624608 99282 624660 99288
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 623688 98660 623740 98666
rect 623688 98602 623740 98608
rect 625620 97980 625672 97986
rect 625620 97922 625672 97928
rect 623136 97708 623188 97714
rect 623136 97650 623188 97656
rect 621664 97572 621716 97578
rect 621664 97514 621716 97520
rect 621664 96348 621716 96354
rect 621664 96290 621716 96296
rect 620468 96076 620520 96082
rect 620468 96018 620520 96024
rect 620928 96076 620980 96082
rect 620928 96018 620980 96024
rect 620480 89690 620508 96018
rect 620468 89684 620520 89690
rect 620468 89626 620520 89632
rect 621676 84182 621704 96290
rect 623044 96212 623096 96218
rect 623044 96154 623096 96160
rect 623056 86494 623084 96154
rect 625344 94648 625396 94654
rect 625344 94590 625396 94596
rect 624424 94512 624476 94518
rect 624424 94454 624476 94460
rect 623044 86488 623096 86494
rect 623044 86430 623096 86436
rect 621664 84176 621716 84182
rect 621664 84118 621716 84124
rect 624436 82929 624464 94454
rect 625356 93854 625384 94590
rect 625264 93826 625384 93854
rect 625264 89729 625292 93826
rect 625632 92585 625660 97922
rect 626092 96898 626120 100014
rect 626828 99210 626856 100014
rect 626816 99204 626868 99210
rect 626816 99146 626868 99152
rect 627564 97442 627592 100014
rect 627552 97436 627604 97442
rect 627552 97378 627604 97384
rect 628208 97306 628236 100014
rect 629036 97986 629064 100014
rect 629772 98938 629800 100014
rect 629760 98932 629812 98938
rect 629760 98874 629812 98880
rect 630508 98802 630536 100014
rect 629484 98796 629536 98802
rect 629484 98738 629536 98744
rect 630496 98796 630548 98802
rect 630496 98738 630548 98744
rect 629024 97980 629076 97986
rect 629024 97922 629076 97928
rect 628380 97572 628432 97578
rect 628380 97514 628432 97520
rect 628196 97300 628248 97306
rect 628196 97242 628248 97248
rect 626264 97164 626316 97170
rect 626264 97106 626316 97112
rect 626080 96892 626132 96898
rect 626080 96834 626132 96840
rect 626276 94489 626304 97106
rect 626448 96076 626500 96082
rect 626448 96018 626500 96024
rect 626460 95441 626488 96018
rect 628392 95826 628420 97514
rect 629496 95826 629524 98738
rect 630864 97708 630916 97714
rect 630864 97650 630916 97656
rect 630876 95826 630904 97650
rect 631244 96626 631272 100014
rect 631888 97578 631916 100014
rect 632152 98660 632204 98666
rect 632152 98602 632204 98608
rect 631876 97572 631928 97578
rect 631876 97514 631928 97520
rect 631232 96620 631284 96626
rect 631232 96562 631284 96568
rect 632164 95826 632192 98602
rect 632716 97850 632744 100014
rect 632980 99340 633032 99346
rect 632980 99282 633032 99288
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 628392 95798 628728 95826
rect 629496 95798 629832 95826
rect 630876 95798 631028 95826
rect 632132 95798 632192 95826
rect 632992 95826 633020 99282
rect 633360 97714 633388 100014
rect 634188 99374 634216 100014
rect 634188 99346 634308 99374
rect 634084 99068 634136 99074
rect 634084 99010 634136 99016
rect 633348 97708 633400 97714
rect 633348 97650 633400 97656
rect 634096 95826 634124 99010
rect 634280 97170 634308 99346
rect 634268 97164 634320 97170
rect 634268 97106 634320 97112
rect 634740 97034 634768 100014
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635280 96892 635332 96898
rect 635280 96834 635332 96840
rect 635292 95826 635320 96834
rect 635476 95946 635504 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 637560 100014 637896 100042
rect 638296 100014 638448 100042
rect 639032 100014 639368 100042
rect 639768 100014 640104 100042
rect 640504 100014 640840 100042
rect 641240 100014 641576 100042
rect 641976 100014 642312 100042
rect 642712 100014 643048 100042
rect 643448 100014 643784 100042
rect 644184 100014 644336 100042
rect 644920 100014 645256 100042
rect 645656 100014 645808 100042
rect 646392 100014 646728 100042
rect 635752 96665 635780 100014
rect 636384 99204 636436 99210
rect 636384 99146 636436 99152
rect 635738 96656 635794 96665
rect 635738 96591 635794 96600
rect 635464 95940 635516 95946
rect 635464 95882 635516 95888
rect 636396 95826 636424 99146
rect 637040 96665 637068 100014
rect 637868 98666 637896 100014
rect 638420 99374 638448 100014
rect 638328 99346 638448 99374
rect 637856 98660 637908 98666
rect 637856 98602 637908 98608
rect 637580 97436 637632 97442
rect 637580 97378 637632 97384
rect 637026 96656 637082 96665
rect 637026 96591 637082 96600
rect 637592 95826 637620 97378
rect 632992 95798 633328 95826
rect 634096 95798 634432 95826
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 638328 95674 638356 99346
rect 639052 97300 639104 97306
rect 639052 97242 639104 97248
rect 639064 95826 639092 97242
rect 639340 95946 639368 100014
rect 639880 97980 639932 97986
rect 639880 97922 639932 97928
rect 639328 95940 639380 95946
rect 639328 95882 639380 95888
rect 639032 95798 639092 95826
rect 639892 95826 639920 97922
rect 640076 96354 640104 100014
rect 640064 96348 640116 96354
rect 640064 96290 640116 96296
rect 640812 96218 640840 100014
rect 640984 98932 641036 98938
rect 640984 98874 641036 98880
rect 640800 96212 640852 96218
rect 640800 96154 640852 96160
rect 640996 95826 641024 98874
rect 641548 96082 641576 100014
rect 642284 96490 642312 100014
rect 642548 98796 642600 98802
rect 642548 98738 642600 98744
rect 642272 96484 642324 96490
rect 642272 96426 642324 96432
rect 641536 96076 641588 96082
rect 641536 96018 641588 96024
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 642560 95690 642588 98738
rect 643020 97986 643048 100014
rect 643008 97980 643060 97986
rect 643008 97922 643060 97928
rect 643284 97844 643336 97850
rect 643284 97786 643336 97792
rect 643296 97594 643324 97786
rect 643468 97708 643520 97714
rect 643468 97650 643520 97656
rect 643296 97566 643416 97594
rect 643192 96620 643244 96626
rect 643192 96562 643244 96568
rect 638132 95668 638184 95674
rect 638132 95610 638184 95616
rect 638316 95668 638368 95674
rect 638316 95610 638368 95616
rect 638592 95668 638644 95674
rect 642528 95662 642588 95690
rect 638592 95610 638644 95616
rect 638144 95554 638172 95610
rect 638604 95554 638632 95610
rect 638144 95526 638632 95554
rect 626446 95432 626502 95441
rect 626446 95367 626502 95376
rect 643204 95169 643232 96562
rect 643190 95160 643246 95169
rect 643190 95095 643246 95104
rect 626262 94480 626318 94489
rect 626262 94415 626318 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 93537 626488 93774
rect 626446 93528 626502 93537
rect 626446 93463 626502 93472
rect 625618 92576 625674 92585
rect 625618 92511 625674 92520
rect 625436 92472 625488 92478
rect 625436 92414 625488 92420
rect 625448 91633 625476 92414
rect 625434 91624 625490 91633
rect 625434 91559 625490 91568
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90681 626488 90986
rect 626446 90672 626502 90681
rect 626446 90607 626502 90616
rect 643388 89729 643416 97566
rect 643480 93854 643508 97650
rect 643756 97306 643784 100014
rect 644308 97442 644336 100014
rect 644940 97572 644992 97578
rect 644940 97514 644992 97520
rect 644296 97436 644348 97442
rect 644296 97378 644348 97384
rect 643744 97300 643796 97306
rect 643744 97242 643796 97248
rect 644756 97164 644808 97170
rect 644756 97106 644808 97112
rect 643744 97028 643796 97034
rect 643744 96970 643796 96976
rect 643480 93826 643600 93854
rect 625250 89720 625306 89729
rect 643374 89720 643430 89729
rect 625250 89655 625306 89664
rect 626448 89684 626500 89690
rect 643374 89655 643430 89664
rect 626448 89626 626500 89632
rect 626460 88913 626488 89626
rect 626446 88904 626502 88913
rect 626446 88839 626502 88848
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 625620 88188 625672 88194
rect 625620 88130 625672 88136
rect 625632 87009 625660 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 643572 87145 643600 93826
rect 643558 87136 643614 87145
rect 643558 87071 643614 87080
rect 625618 87000 625674 87009
rect 625618 86935 625674 86944
rect 626448 86488 626500 86494
rect 626448 86430 626500 86436
rect 626460 86057 626488 86430
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 625620 84176 625672 84182
rect 625618 84144 625620 84153
rect 625672 84144 625674 84153
rect 625618 84079 625674 84088
rect 624422 82920 624478 82929
rect 624422 82855 624478 82864
rect 643756 82793 643784 96970
rect 644480 96620 644532 96626
rect 644480 96562 644532 96568
rect 643928 96348 643980 96354
rect 643928 96290 643980 96296
rect 643940 95946 643968 96290
rect 643928 95940 643980 95946
rect 643928 95882 643980 95888
rect 644492 93838 644520 96562
rect 644480 93832 644532 93838
rect 644480 93774 644532 93780
rect 644768 84697 644796 97106
rect 644952 92177 644980 97514
rect 645228 96966 645256 100014
rect 645216 96960 645268 96966
rect 645216 96902 645268 96908
rect 644938 92168 644994 92177
rect 644938 92103 644994 92112
rect 645780 88806 645808 100014
rect 646700 96762 646728 100014
rect 647114 99770 647142 100028
rect 647864 100014 648200 100042
rect 648600 100014 648936 100042
rect 649336 100014 649672 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 647114 99742 647188 99770
rect 647160 97714 647188 99742
rect 647148 97708 647200 97714
rect 647148 97650 647200 97656
rect 646688 96756 646740 96762
rect 646688 96698 646740 96704
rect 647884 96756 647936 96762
rect 647884 96698 647936 96704
rect 647700 96484 647752 96490
rect 647700 96426 647752 96432
rect 647712 95946 647740 96426
rect 647700 95940 647752 95946
rect 647700 95882 647752 95888
rect 646044 95804 646096 95810
rect 646044 95746 646096 95752
rect 645768 88800 645820 88806
rect 645768 88742 645820 88748
rect 644754 84688 644810 84697
rect 644754 84623 644810 84632
rect 643742 82784 643798 82793
rect 643742 82719 643798 82728
rect 628654 81696 628710 81705
rect 628654 81631 628710 81640
rect 628668 80986 628696 81631
rect 628656 80980 628708 80986
rect 628656 80922 628708 80928
rect 631520 80974 631856 81002
rect 639064 80974 639308 81002
rect 642456 80980 642508 80986
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 629220 79490 629248 80815
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 628196 77580 628248 77586
rect 628196 77522 628248 77528
rect 628208 77314 628236 77522
rect 631060 77450 631088 78066
rect 631048 77444 631100 77450
rect 631048 77386 631100 77392
rect 628196 77308 628248 77314
rect 628196 77250 628248 77256
rect 628380 77308 628432 77314
rect 628380 77250 628432 77256
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 628392 75290 628420 77250
rect 631060 75290 631088 77386
rect 631520 77314 631548 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 80472 633954 80481
rect 633898 80407 633954 80416
rect 633912 77586 633940 80407
rect 633900 77580 633952 77586
rect 633900 77522 633952 77528
rect 631508 77308 631560 77314
rect 631508 77250 631560 77256
rect 633912 75290 633940 77522
rect 636120 77294 636148 80650
rect 638868 79484 638920 79490
rect 638868 79426 638920 79432
rect 638880 78334 638908 79426
rect 638868 78328 638920 78334
rect 638868 78270 638920 78276
rect 639064 78130 639092 80974
rect 642456 80922 642508 80928
rect 639052 78124 639104 78130
rect 639052 78066 639104 78072
rect 639602 77888 639658 77897
rect 639602 77823 639658 77832
rect 636120 77266 636332 77294
rect 628176 75276 628420 75290
rect 628162 75262 628420 75276
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 618904 75200 618956 75206
rect 618904 75142 618956 75148
rect 628162 74882 628190 75262
rect 636304 75154 636332 77266
rect 639616 75290 639644 77823
rect 642468 75290 642496 80922
rect 645308 78328 645360 78334
rect 645308 78270 645360 78276
rect 645320 75290 645348 78270
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 628024 74868 628190 74882
rect 628024 74866 628176 74868
rect 628012 74860 628176 74866
rect 628064 74854 628176 74860
rect 628012 74802 628064 74808
rect 624424 67652 624476 67658
rect 624424 67594 624476 67600
rect 614856 60716 614908 60722
rect 614856 60658 614908 60664
rect 605840 58676 605892 58682
rect 605840 58618 605892 58624
rect 624436 55894 624464 67594
rect 646056 64874 646084 95746
rect 646228 95668 646280 95674
rect 646228 95610 646280 95616
rect 646240 68921 646268 95610
rect 647896 87174 647924 96698
rect 648172 96490 648200 100014
rect 648160 96484 648212 96490
rect 648160 96426 648212 96432
rect 648908 95810 648936 100014
rect 649264 96960 649316 96966
rect 649264 96902 649316 96908
rect 648896 95804 648948 95810
rect 648896 95746 648948 95752
rect 648528 95532 648580 95538
rect 648528 95474 648580 95480
rect 648540 92478 648568 95474
rect 648528 92472 648580 92478
rect 648528 92414 648580 92420
rect 647884 87168 647936 87174
rect 647884 87110 647936 87116
rect 649276 86902 649304 96902
rect 649644 96626 649672 100014
rect 650380 97170 650408 100014
rect 651116 97306 651144 100014
rect 650828 97300 650880 97306
rect 650828 97242 650880 97248
rect 651104 97300 651156 97306
rect 651104 97242 651156 97248
rect 650368 97164 650420 97170
rect 650368 97106 650420 97112
rect 649632 96620 649684 96626
rect 649632 96562 649684 96568
rect 650644 96620 650696 96626
rect 650644 96562 650696 96568
rect 649264 86896 649316 86902
rect 649264 86838 649316 86844
rect 650656 86766 650684 96562
rect 650840 87038 650868 97242
rect 651852 97034 651880 100014
rect 651840 97028 651892 97034
rect 651840 96970 651892 96976
rect 652588 96626 652616 100014
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 650828 87032 650880 87038
rect 650828 86974 650880 86980
rect 650644 86760 650696 86766
rect 650644 86702 650696 86708
rect 652036 86630 652064 96426
rect 653324 96354 653352 100014
rect 653968 96830 653996 100014
rect 654600 97436 654652 97442
rect 654600 97378 654652 97384
rect 654612 97034 654640 97378
rect 654600 97028 654652 97034
rect 654600 96970 654652 96976
rect 654796 96966 654824 100014
rect 655440 97714 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97708 655480 97714
rect 655428 97650 655480 97656
rect 655060 97300 655112 97306
rect 655060 97242 655112 97248
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 653956 96824 654008 96830
rect 653956 96766 654008 96772
rect 653864 96484 653916 96490
rect 653864 96426 653916 96432
rect 653312 96348 653364 96354
rect 653312 96290 653364 96296
rect 653404 95940 653456 95946
rect 653404 95882 653456 95888
rect 652024 86624 652076 86630
rect 652024 86566 652076 86572
rect 653416 86494 653444 95882
rect 653876 90794 653904 96426
rect 654876 93832 654928 93838
rect 654876 93774 654928 93780
rect 654888 92585 654916 93774
rect 655072 93401 655100 97242
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655244 96824 655296 96830
rect 655244 96766 655296 96772
rect 655256 94217 655284 96766
rect 655242 94208 655298 94217
rect 655242 94143 655298 94152
rect 655058 93392 655114 93401
rect 655058 93327 655114 93336
rect 655440 92698 655468 96902
rect 655072 92670 655468 92698
rect 654874 92576 654930 92585
rect 654874 92511 654930 92520
rect 653876 90766 654180 90794
rect 654152 90681 654180 90766
rect 654138 90672 654194 90681
rect 654138 90607 654194 90616
rect 655072 88330 655100 92670
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655808 89865 655836 100014
rect 656820 97306 656848 100014
rect 657544 97844 657596 97850
rect 657544 97786 657596 97792
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 657556 96830 657584 97786
rect 657544 96824 657596 96830
rect 657544 96766 657596 96772
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97986 658228 99742
rect 658188 97980 658240 97986
rect 658188 97922 658240 97928
rect 659212 97714 659240 100014
rect 659948 97850 659976 100014
rect 660396 98660 660448 98666
rect 660396 98602 660448 98608
rect 659752 97844 659804 97850
rect 659752 97786 659804 97792
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659200 97708 659252 97714
rect 659200 97650 659252 97656
rect 658832 97572 658884 97578
rect 658832 97514 658884 97520
rect 658280 97164 658332 97170
rect 658280 97106 658332 97112
rect 658292 95132 658320 97106
rect 658844 95132 658872 97514
rect 659568 97436 659620 97442
rect 659568 97378 659620 97384
rect 659580 95132 659608 97378
rect 659764 95146 659792 97786
rect 660408 95146 660436 98602
rect 660684 96966 660712 100014
rect 663064 97980 663116 97986
rect 663064 97922 663116 97928
rect 662512 97572 662564 97578
rect 662512 97514 662564 97520
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660672 96960 660724 96966
rect 660672 96902 660724 96908
rect 659764 95118 660146 95146
rect 660408 95118 660698 95146
rect 661420 95132 661448 97242
rect 661960 96824 662012 96830
rect 661960 96766 662012 96772
rect 661972 95132 662000 96766
rect 662524 95132 662552 97514
rect 663076 95132 663104 97922
rect 665180 97844 665232 97850
rect 665180 97786 665232 97792
rect 663892 97708 663944 97714
rect 663892 97650 663944 97656
rect 663432 96960 663484 96966
rect 663432 96902 663484 96908
rect 663248 96076 663300 96082
rect 663248 96018 663300 96024
rect 663260 93129 663288 96018
rect 663246 93120 663302 93129
rect 663246 93055 663302 93064
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 657452 88800 657504 88806
rect 662328 88800 662380 88806
rect 657504 88748 657754 88754
rect 657452 88742 657754 88748
rect 657464 88726 657754 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 655060 88324 655112 88330
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 655060 88266 655112 88272
rect 658464 88266 658516 88272
rect 657188 87174 657216 88196
rect 657176 87168 657228 87174
rect 657176 87110 657228 87116
rect 658844 86766 658872 88196
rect 659580 86766 659608 88196
rect 658832 86760 658884 86766
rect 658832 86702 658884 86708
rect 659568 86760 659620 86766
rect 659568 86702 659620 86708
rect 660132 86494 660160 88196
rect 660684 86902 660712 88196
rect 661420 87038 661448 88196
rect 661408 87032 661460 87038
rect 661408 86974 661460 86980
rect 660672 86896 660724 86902
rect 660672 86838 660724 86844
rect 662524 86630 662552 88196
rect 663444 86766 663472 96902
rect 663708 96212 663760 96218
rect 663708 96154 663760 96160
rect 663720 96098 663748 96154
rect 663720 96070 663840 96098
rect 663812 92154 663840 96070
rect 663720 92126 663840 92154
rect 663720 92041 663748 92126
rect 663706 92032 663762 92041
rect 663706 91967 663762 91976
rect 663904 88806 663932 97650
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89049 664208 96290
rect 664628 95940 664680 95946
rect 664628 95882 664680 95888
rect 664444 92540 664496 92546
rect 664444 92482 664496 92488
rect 664166 89040 664222 89049
rect 664166 88975 664222 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663432 86760 663484 86766
rect 663432 86702 663484 86708
rect 662512 86624 662564 86630
rect 662512 86566 662564 86572
rect 653404 86488 653456 86494
rect 653404 86430 653456 86436
rect 660120 86488 660172 86494
rect 660120 86430 660172 86436
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 647056 76696 647108 76702
rect 647056 76638 647108 76644
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646884 73001 646912 75142
rect 647068 74497 647096 76638
rect 647054 74488 647110 74497
rect 647054 74423 647110 74432
rect 646870 72992 646926 73001
rect 646870 72927 646926 72936
rect 647344 70009 647372 80786
rect 648988 79348 649040 79354
rect 648988 79290 649040 79296
rect 647516 77988 647568 77994
rect 647516 77930 647568 77936
rect 647330 70000 647386 70009
rect 647330 69935 647386 69944
rect 646226 68912 646282 68921
rect 646226 68847 646282 68856
rect 647528 65521 647556 77930
rect 649000 71505 649028 79290
rect 649172 76832 649224 76838
rect 649172 76774 649224 76780
rect 648986 71496 649042 71505
rect 648986 71431 649042 71440
rect 649184 67017 649212 76774
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 649170 67008 649226 67017
rect 649170 66943 649226 66952
rect 647514 65512 647570 65521
rect 647514 65447 647570 65456
rect 646056 64846 646176 64874
rect 646148 64433 646176 64846
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 624424 55888 624476 55894
rect 624424 55830 624476 55836
rect 597652 54470 597704 54476
rect 604458 54496 604514 54505
rect 604458 54431 604514 54440
rect 579068 54198 579120 54204
rect 580262 54224 580318 54233
rect 580262 54159 580318 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459468 53644 459520 53650
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 462594 53615 462650 53624
rect 465172 53644 465224 53650
rect 459468 53586 459520 53592
rect 129004 53372 129056 53378
rect 129004 53314 129056 53320
rect 127164 51876 127216 51882
rect 127164 51818 127216 51824
rect 127176 50794 127204 51818
rect 127164 50788 127216 50794
rect 127164 50730 127216 50736
rect 129016 50674 129044 53314
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 129464 51740 129516 51746
rect 129464 51682 129516 51688
rect 129280 50788 129332 50794
rect 129280 50730 129332 50736
rect 129016 50646 129228 50674
rect 128636 50516 128688 50522
rect 128636 50458 128688 50464
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 128452 49156 128504 49162
rect 128452 49098 128504 49104
rect 47584 49020 47636 49026
rect 47584 48962 47636 48968
rect 128464 44810 128492 49098
rect 128648 47870 128676 50458
rect 129004 50380 129056 50386
rect 129004 50322 129056 50328
rect 128636 47864 128688 47870
rect 128636 47806 128688 47812
rect 128452 44804 128504 44810
rect 128452 44746 128504 44752
rect 129016 44198 129044 50322
rect 129200 44470 129228 50646
rect 129292 48314 129320 50730
rect 129292 48286 129412 48314
rect 129384 44606 129412 48286
rect 129476 47274 129504 51682
rect 129648 49020 129700 49026
rect 129648 48962 129700 48968
rect 129660 48314 129688 48962
rect 129660 48286 129780 48314
rect 129476 47246 129596 47274
rect 129568 45082 129596 47246
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129752 44946 129780 48286
rect 129740 44940 129792 44946
rect 129740 44882 129792 44888
rect 129372 44600 129424 44606
rect 129372 44542 129424 44548
rect 129188 44464 129240 44470
rect 129188 44406 129240 44412
rect 129004 44192 129056 44198
rect 129004 44134 129056 44140
rect 130396 43926 130424 53178
rect 312360 53168 312412 53174
rect 130568 53100 130620 53106
rect 130568 53042 130620 53048
rect 130580 44062 130608 53042
rect 306024 52494 306052 53108
rect 145380 52488 145432 52494
rect 145380 52430 145432 52436
rect 306012 52488 306064 52494
rect 306012 52430 306064 52436
rect 130752 52012 130804 52018
rect 130752 51954 130804 51960
rect 130764 44334 130792 51954
rect 145392 50810 145420 52430
rect 145084 50782 145420 50810
rect 308048 50289 308076 53108
rect 309704 53094 310040 53122
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 309704 49745 309732 53094
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53586
rect 459848 52578 459876 53615
rect 460066 52828 460118 52834
rect 460066 52770 460118 52776
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460078 52564 460106 52770
rect 460768 52578 460796 53615
rect 461308 53508 461360 53514
rect 461308 53450 461360 53456
rect 461320 52578 461348 53450
rect 461688 52578 461716 53615
rect 461904 52864 461960 52873
rect 461904 52799 461960 52808
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461918 52564 461946 52799
rect 462608 52578 462636 53615
rect 465172 53586 465224 53592
rect 465724 53644 465776 53650
rect 465724 53586 465776 53592
rect 465908 53644 465960 53650
rect 465908 53586 465960 53592
rect 469956 53644 470008 53650
rect 469956 53586 470008 53592
rect 470140 53644 470192 53650
rect 470140 53586 470192 53592
rect 470416 53644 470468 53650
rect 470416 53586 470468 53592
rect 477960 53644 478012 53650
rect 477960 53586 478012 53592
rect 481732 53644 481784 53650
rect 481732 53586 481784 53592
rect 482008 53644 482060 53650
rect 482008 53586 482060 53592
rect 463608 53372 463660 53378
rect 463608 53314 463660 53320
rect 463148 53236 463200 53242
rect 463148 53178 463200 53184
rect 463160 52578 463188 53178
rect 463620 52578 463648 53314
rect 464896 53100 464948 53106
rect 464896 53042 464948 53048
rect 464068 52964 464120 52970
rect 464068 52906 464120 52912
rect 464080 52578 464108 52906
rect 464206 52828 464258 52834
rect 464206 52770 464258 52776
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463772 52550 464108 52578
rect 464218 52564 464246 52770
rect 464908 52578 464936 53042
rect 464692 52550 464936 52578
rect 465184 52442 465212 53586
rect 465736 52873 465764 53586
rect 465722 52864 465778 52873
rect 465722 52799 465778 52808
rect 465920 52578 465948 53586
rect 469968 52834 469996 53586
rect 470152 53378 470180 53586
rect 470140 53372 470192 53378
rect 470140 53314 470192 53320
rect 469956 52828 470008 52834
rect 469956 52770 470008 52776
rect 470428 52698 470456 53586
rect 477972 53242 478000 53586
rect 477960 53236 478012 53242
rect 477960 53178 478012 53184
rect 481744 53106 481772 53586
rect 481732 53100 481784 53106
rect 481732 53042 481784 53048
rect 482020 52970 482048 53586
rect 482008 52964 482060 52970
rect 482008 52906 482060 52912
rect 470416 52692 470468 52698
rect 470416 52634 470468 52640
rect 465612 52550 465948 52578
rect 465152 52414 465212 52442
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 309690 49736 309746 49745
rect 309690 49671 309746 49680
rect 132132 47864 132184 47870
rect 132132 47806 132184 47812
rect 132144 44506 132172 47806
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132132 44500 132184 44506
rect 132132 44442 132184 44448
rect 132408 44464 132460 44470
rect 132236 44412 132408 44418
rect 132236 44406 132460 44412
rect 132236 44390 132448 44406
rect 130752 44328 130804 44334
rect 130752 44270 130804 44276
rect 132236 44198 132264 44390
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 132224 44192 132276 44198
rect 132224 44134 132276 44140
rect 310426 44160 310482 44169
rect 310426 44095 310482 44104
rect 364890 44160 364946 44169
rect 364890 44095 364946 44104
rect 130568 44056 130620 44062
rect 130568 43998 130620 44004
rect 130384 43920 130436 43926
rect 130384 43862 130436 43868
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 43444 42832 43496 42838
rect 43444 42774 43496 42780
rect 187344 42092 187372 43522
rect 308954 42800 309010 42809
rect 307300 42764 307352 42770
rect 308954 42735 309010 42744
rect 307300 42706 307352 42712
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 42706
rect 308968 42231 308996 42735
rect 308956 42225 309008 42231
rect 308956 42167 309008 42173
rect 310440 42106 310468 44095
rect 361764 42492 361816 42498
rect 361764 42434 361816 42440
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 42434
rect 364904 42092 364932 44095
rect 431236 43654 431264 44775
rect 431224 43648 431276 43654
rect 431224 43590 431276 43596
rect 369400 42764 369452 42770
rect 369400 42706 369452 42712
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 369412 42498 369440 42706
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 369400 42492 369452 42498
rect 369400 42434 369452 42440
rect 416594 42392 416650 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 416594 42327 416650 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 194322 42055 194378 42064
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415766 42120 415822 42129
rect 405200 42078 405582 42106
rect 415426 42078 415766 42106
rect 416608 42092 416636 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 415766 42055 415822 42064
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42090 427124 42570
rect 431236 42090 431264 42706
rect 455880 42628 455932 42634
rect 455880 42570 455932 42576
rect 443550 42256 443606 42265
rect 443550 42191 443606 42200
rect 427084 42084 427136 42090
rect 427084 42026 427136 42032
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 443564 41585 443592 42191
rect 455892 41954 455920 42570
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 455880 41948 455932 41954
rect 455880 41890 455932 41896
rect 443550 41576 443606 41585
rect 443550 41511 443606 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460860 43489 460888 47654
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461964 44441 461992 47654
rect 462378 47410 462406 47668
rect 462332 47382 462406 47410
rect 462516 47654 462852 47682
rect 462976 47654 463312 47682
rect 461950 44432 462006 44441
rect 461950 44367 462006 44376
rect 462332 43217 462360 47382
rect 462516 44441 462544 47654
rect 462502 44432 462558 44441
rect 462502 44367 462558 44376
rect 462976 43897 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463988 47654 464232 47682
rect 464356 47654 464692 47682
rect 463712 44169 463740 47382
rect 463698 44160 463754 44169
rect 463698 44095 463754 44104
rect 462962 43888 463018 43897
rect 462962 43823 463018 43832
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 463698 42936 463754 42945
rect 463698 42871 463754 42880
rect 463712 42378 463740 42871
rect 463988 42634 464016 47654
rect 464356 42770 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 544028 47569 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 544014 47560 544070 47569
rect 544014 47495 544070 47504
rect 545684 47297 545712 53094
rect 547892 47841 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 48113 552060 53108
rect 553688 53094 554024 53122
rect 553688 50289 553716 53094
rect 553674 50280 553730 50289
rect 553674 50215 553730 50224
rect 552018 48104 552074 48113
rect 552018 48039 552074 48048
rect 547878 47832 547934 47841
rect 547878 47767 547934 47776
rect 662432 47433 662460 76502
rect 664456 62082 664484 92482
rect 664640 89865 664668 95882
rect 665192 93401 665220 97786
rect 665364 96620 665416 96626
rect 665364 96562 665416 96568
rect 665178 93392 665234 93401
rect 665178 93327 665234 93336
rect 665376 90681 665404 96562
rect 665362 90672 665418 90681
rect 665362 90607 665418 90616
rect 664626 89856 664682 89865
rect 664626 89791 664682 89800
rect 666664 84194 666692 105975
rect 668044 100162 668072 109239
rect 668320 104417 668348 111823
rect 670712 106214 670740 113146
rect 671540 107681 671568 130863
rect 671908 115841 671936 166903
rect 672092 140321 672120 183495
rect 672460 177857 672488 235690
rect 672644 230353 672672 249070
rect 672602 230344 672672 230353
rect 672658 230302 672672 230344
rect 672602 230279 672658 230288
rect 672736 227576 672764 251146
rect 672828 229094 672856 392527
rect 673012 378049 673040 397151
rect 672998 378040 673054 378049
rect 672998 377975 673054 377984
rect 673196 355065 673224 398783
rect 673366 396400 673422 396409
rect 673366 396335 673422 396344
rect 673380 382265 673408 396335
rect 673826 396128 673882 396137
rect 673826 396063 673882 396072
rect 673366 382256 673422 382265
rect 673366 382191 673422 382200
rect 673840 381449 673868 396063
rect 674010 395720 674066 395729
rect 674010 395655 674066 395664
rect 673826 381440 673882 381449
rect 673826 381375 673882 381384
rect 674024 375465 674052 395655
rect 674010 375456 674066 375465
rect 674010 375391 674066 375400
rect 674208 356697 674236 401367
rect 674470 394496 674526 394505
rect 674470 394431 674526 394440
rect 674484 377777 674512 394431
rect 674470 377768 674526 377777
rect 674470 377703 674526 377712
rect 674668 357513 674696 402183
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675114 377768 675170 377777
rect 675170 377726 675340 377754
rect 675114 377703 675170 377712
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675206 377496 675262 377505
rect 675206 377431 675262 377440
rect 675220 373994 675248 377431
rect 675758 377224 675814 377233
rect 675758 377159 675814 377168
rect 675772 377060 675800 377159
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675390 375456 675446 375465
rect 675390 375391 675446 375400
rect 675404 375224 675432 375391
rect 675220 373966 675340 373994
rect 675312 373402 675340 373966
rect 675312 373374 675418 373402
rect 675758 373008 675814 373017
rect 675758 372943 675814 372952
rect 675772 372776 675800 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 357504 674710 357513
rect 674654 357439 674710 357448
rect 674654 357096 674710 357105
rect 674654 357031 674710 357040
rect 674194 356688 674250 356697
rect 674194 356623 674250 356632
rect 674102 356280 674158 356289
rect 674102 356215 674158 356224
rect 673182 355056 673238 355065
rect 673182 354991 673238 355000
rect 672998 354648 673054 354657
rect 672998 354583 673054 354592
rect 673012 310049 673040 354583
rect 673182 353424 673238 353433
rect 673182 353359 673238 353368
rect 673196 340785 673224 353359
rect 673918 352608 673974 352617
rect 673918 352543 673974 352552
rect 673550 352200 673606 352209
rect 673550 352135 673606 352144
rect 673366 349752 673422 349761
rect 673366 349687 673422 349696
rect 673182 340776 673238 340785
rect 673182 340711 673238 340720
rect 673380 335889 673408 349687
rect 673366 335880 673422 335889
rect 673366 335815 673422 335824
rect 673564 325689 673592 352135
rect 673734 350568 673790 350577
rect 673734 350503 673790 350512
rect 673748 331129 673776 350503
rect 673932 336705 673960 352543
rect 673918 336696 673974 336705
rect 673918 336631 673974 336640
rect 673734 331120 673790 331129
rect 673734 331055 673790 331064
rect 673550 325680 673606 325689
rect 673550 325615 673606 325624
rect 673918 312080 673974 312089
rect 673918 312015 673974 312024
rect 673182 311264 673238 311273
rect 673182 311199 673238 311208
rect 672998 310040 673054 310049
rect 672998 309975 673054 309984
rect 672998 304328 673054 304337
rect 672998 304263 673054 304272
rect 673012 287881 673040 304263
rect 672998 287872 673054 287881
rect 672998 287807 673054 287816
rect 673196 266529 673224 311199
rect 673734 305552 673790 305561
rect 673734 305487 673790 305496
rect 673366 304736 673422 304745
rect 673366 304671 673422 304680
rect 673380 290057 673408 304671
rect 673366 290048 673422 290057
rect 673366 289983 673422 289992
rect 673748 285569 673776 305487
rect 673734 285560 673790 285569
rect 673734 285495 673790 285504
rect 673932 267481 673960 312015
rect 674116 311681 674144 356215
rect 674470 349480 674526 349489
rect 674470 349415 674526 349424
rect 674286 347712 674342 347721
rect 674286 347647 674342 347656
rect 674300 327593 674328 347647
rect 674484 332897 674512 349415
rect 674668 340874 674696 357031
rect 676034 353832 676090 353841
rect 676090 353790 676260 353818
rect 676034 353767 676090 353776
rect 675942 349208 675998 349217
rect 676232 349194 676260 353790
rect 675998 349166 676260 349194
rect 675942 349143 675998 349152
rect 674576 340846 674696 340874
rect 674576 338114 674604 340846
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675404 339017 675432 339252
rect 675390 339008 675446 339017
rect 675390 338943 675446 338952
rect 674576 338086 674696 338114
rect 674470 332888 674526 332897
rect 674470 332823 674526 332832
rect 674286 327584 674342 327593
rect 674286 327519 674342 327528
rect 674668 312497 674696 338086
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675312 336829 675418 336857
rect 675114 336696 675170 336705
rect 675114 336631 675170 336640
rect 675128 333078 675156 336631
rect 675312 335345 675340 336829
rect 675758 336696 675814 336705
rect 675758 336631 675814 336640
rect 675772 336192 675800 336631
rect 675482 335880 675538 335889
rect 675482 335815 675538 335824
rect 675496 335580 675524 335815
rect 675298 335336 675354 335345
rect 675298 335271 675354 335280
rect 675128 333050 675418 333078
rect 675390 332888 675446 332897
rect 675390 332823 675446 332832
rect 675404 332520 675432 332823
rect 675114 332344 675170 332353
rect 675114 332279 675170 332288
rect 675128 331242 675156 332279
rect 675758 332208 675814 332217
rect 675758 332143 675814 332152
rect 675772 331875 675800 332143
rect 675128 331214 675418 331242
rect 675114 331120 675170 331129
rect 675114 331055 675170 331064
rect 675128 330049 675156 331055
rect 675128 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675114 327584 675170 327593
rect 675170 327542 675418 327570
rect 675114 327519 675170 327528
rect 675312 326454 675432 326482
rect 675312 326346 675340 326454
rect 675128 326318 675340 326346
rect 675404 326332 675432 326454
rect 675128 325689 675156 326318
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 312488 674710 312497
rect 674654 312423 674710 312432
rect 674102 311672 674158 311681
rect 674102 311607 674158 311616
rect 674470 310448 674526 310457
rect 674470 310383 674526 310392
rect 674194 309632 674250 309641
rect 674194 309567 674250 309576
rect 673918 267472 673974 267481
rect 673918 267407 673974 267416
rect 673182 266520 673238 266529
rect 673182 266455 673238 266464
rect 674010 266248 674066 266257
rect 674010 266183 674066 266192
rect 673182 263800 673238 263809
rect 673182 263735 673238 263744
rect 672998 260128 673054 260137
rect 672998 260063 673054 260072
rect 673012 245041 673040 260063
rect 672998 245032 673054 245041
rect 672998 244967 673054 244976
rect 673196 244274 673224 263735
rect 674024 263594 674052 266183
rect 674208 265033 674236 309567
rect 674484 265849 674512 310383
rect 674838 309224 674894 309233
rect 674838 309159 674894 309168
rect 674654 303920 674710 303929
rect 674654 303855 674710 303864
rect 674668 286226 674696 303855
rect 674852 298081 674880 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675022 308000 675078 308009
rect 675022 307935 675078 307944
rect 675036 302234 675064 307935
rect 676232 304994 676260 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 676402 305960 676458 305969
rect 676402 305895 676458 305904
rect 675864 304966 676260 304994
rect 675864 302234 675892 304966
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 675036 302206 675248 302234
rect 675220 299474 675248 302206
rect 675128 299446 675248 299474
rect 675772 302206 675892 302234
rect 674838 298072 674894 298081
rect 674838 298007 674894 298016
rect 675128 297922 675156 299446
rect 675298 298072 675354 298081
rect 675298 298007 675354 298016
rect 675128 297894 675248 297922
rect 674838 296848 674894 296857
rect 674838 296783 674894 296792
rect 674852 288062 674880 296783
rect 675022 296576 675078 296585
rect 675022 296511 675078 296520
rect 675036 292574 675064 296511
rect 675036 292546 675156 292574
rect 675128 291870 675156 292546
rect 675220 292414 675248 297894
rect 675312 294250 675340 298007
rect 675772 296313 675800 302206
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676416 301617 676444 305895
rect 676678 305144 676734 305153
rect 676678 305079 676734 305088
rect 676402 301608 676458 301617
rect 676402 301543 676458 301552
rect 676692 301481 676720 305079
rect 676678 301472 676734 301481
rect 676678 301407 676734 301416
rect 675944 298104 675996 298110
rect 675944 298046 675996 298052
rect 675956 296585 675984 298046
rect 676128 297900 676180 297906
rect 676128 297842 676180 297848
rect 676140 296857 676168 297842
rect 678256 297401 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 681016 297906 681044 307527
rect 681004 297900 681056 297906
rect 681004 297842 681056 297848
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 676126 296848 676182 296857
rect 676126 296783 676182 296792
rect 675942 296576 675998 296585
rect 675942 296511 675998 296520
rect 675758 296304 675814 296313
rect 675758 296239 675814 296248
rect 675758 295896 675814 295905
rect 675758 295831 675814 295840
rect 675772 295528 675800 295831
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675312 294222 675418 294250
rect 675220 292386 675418 292414
rect 675128 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675128 290550 675418 290578
rect 675128 290057 675156 290550
rect 675114 290048 675170 290057
rect 675114 289983 675170 289992
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675312 286334 675432 286362
rect 675312 286226 675340 286334
rect 674668 286198 675340 286226
rect 675404 286212 675432 286334
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 676034 269784 676090 269793
rect 676034 269719 676090 269728
rect 676048 268297 676076 269719
rect 676034 268288 676090 268297
rect 676034 268223 676090 268232
rect 683132 268161 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 674654 267064 674710 267073
rect 674654 266999 674710 267008
rect 674470 265840 674526 265849
rect 674470 265775 674526 265784
rect 674378 265432 674434 265441
rect 674378 265367 674434 265376
rect 674194 265024 674250 265033
rect 674194 264959 674250 264968
rect 674392 263594 674420 265367
rect 674024 263566 674144 263594
rect 674392 263566 674512 263594
rect 673734 259720 673790 259729
rect 673734 259655 673790 259664
rect 673366 259312 673422 259321
rect 673366 259247 673422 259256
rect 673012 244246 673224 244274
rect 673012 233986 673040 244246
rect 673380 242865 673408 259247
rect 673748 245585 673776 259655
rect 673918 258496 673974 258505
rect 673918 258431 673974 258440
rect 673734 245576 673790 245585
rect 673734 245511 673790 245520
rect 673366 242856 673422 242865
rect 673366 242791 673422 242800
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673184 236768 673236 236774
rect 673184 236710 673236 236716
rect 673000 233980 673052 233986
rect 673000 233922 673052 233928
rect 673196 233209 673224 236710
rect 673426 236450 673454 236846
rect 673526 236736 673582 236745
rect 673526 236671 673528 236680
rect 673580 236671 673582 236680
rect 673528 236642 673580 236648
rect 673644 236564 673696 236570
rect 673644 236506 673696 236512
rect 673426 236422 673592 236450
rect 673368 236292 673420 236298
rect 673368 236234 673420 236240
rect 673380 236178 673408 236234
rect 673380 236150 673500 236178
rect 673304 236088 673356 236094
rect 673288 236036 673304 236042
rect 673288 236030 673356 236036
rect 673288 236014 673344 236030
rect 673288 234614 673316 236014
rect 673288 234586 673408 234614
rect 673182 233200 673238 233209
rect 673182 233135 673238 233144
rect 673380 233050 673408 234586
rect 672920 233022 673408 233050
rect 672920 231792 672948 233022
rect 673182 232928 673238 232937
rect 673472 232914 673500 236150
rect 673238 232886 673500 232914
rect 673182 232863 673238 232872
rect 672920 231764 673040 231792
rect 673012 231441 673040 231764
rect 673368 231600 673420 231606
rect 673368 231542 673420 231548
rect 672998 231432 673054 231441
rect 672998 231367 673054 231376
rect 673092 230852 673144 230858
rect 673092 230794 673144 230800
rect 673104 229809 673132 230794
rect 673380 230353 673408 231542
rect 673366 230344 673422 230353
rect 673366 230279 673422 230288
rect 673564 230194 673592 236422
rect 673288 230166 673592 230194
rect 673090 229800 673146 229809
rect 673090 229735 673146 229744
rect 673090 229528 673146 229537
rect 673090 229463 673146 229472
rect 673104 229362 673132 229463
rect 673092 229356 673144 229362
rect 673092 229298 673144 229304
rect 673288 229226 673316 230166
rect 673458 230072 673514 230081
rect 673458 230007 673514 230016
rect 673472 229498 673500 230007
rect 673460 229492 673512 229498
rect 673460 229434 673512 229440
rect 673276 229220 673328 229226
rect 673276 229162 673328 229168
rect 673458 229120 673514 229129
rect 672828 229066 672948 229094
rect 672920 228721 672948 229066
rect 673458 229055 673460 229064
rect 673512 229055 673514 229064
rect 673460 229026 673512 229032
rect 673506 228880 673558 228886
rect 673504 228848 673506 228857
rect 673558 228848 673560 228857
rect 673504 228783 673560 228792
rect 672906 228712 672962 228721
rect 672906 228647 672962 228656
rect 673386 228576 673442 228585
rect 673386 228511 673388 228520
rect 673440 228511 673442 228520
rect 673388 228482 673440 228488
rect 673046 227928 673098 227934
rect 673098 227876 673316 227882
rect 673046 227870 673316 227876
rect 673058 227854 673316 227870
rect 673288 227780 673316 227854
rect 673288 227752 673500 227780
rect 672954 227724 673006 227730
rect 672954 227666 673006 227672
rect 672966 227610 672994 227666
rect 672966 227582 673224 227610
rect 672552 227548 672764 227576
rect 672552 209774 672580 227548
rect 672816 227520 672868 227526
rect 672816 227462 672868 227468
rect 673196 227474 673224 227582
rect 672828 227372 672856 227462
rect 673196 227446 673316 227474
rect 672828 227344 672948 227372
rect 672724 227316 672776 227322
rect 672724 227258 672776 227264
rect 672736 224618 672764 227258
rect 672920 224754 672948 227344
rect 673288 227236 673316 227446
rect 673196 227208 673316 227236
rect 673196 226817 673224 227208
rect 673472 226896 673500 227752
rect 673472 226868 673546 226896
rect 673182 226808 673238 226817
rect 673182 226743 673238 226752
rect 673518 226658 673546 226868
rect 673380 226630 673546 226658
rect 673182 225176 673238 225185
rect 673182 225111 673238 225120
rect 672920 224726 673132 224754
rect 672906 224632 672962 224641
rect 672736 224590 672906 224618
rect 672906 224567 672962 224576
rect 672722 224360 672778 224369
rect 672722 224295 672778 224304
rect 672736 222194 672764 224295
rect 673104 222194 673132 224726
rect 672644 222166 672764 222194
rect 672828 222166 673132 222194
rect 672644 219434 672672 222166
rect 672828 220425 672856 222166
rect 672814 220416 672870 220425
rect 672814 220351 672870 220360
rect 672644 219406 672764 219434
rect 672736 214713 672764 219406
rect 673196 215294 673224 225111
rect 673380 222194 673408 226630
rect 673504 225448 673560 225457
rect 673504 225383 673560 225392
rect 673518 225298 673546 225383
rect 673518 225270 673592 225298
rect 673380 222166 673500 222194
rect 673472 216322 673500 222166
rect 673564 220810 673592 225270
rect 673656 222194 673684 236506
rect 673932 230466 673960 258431
rect 674116 235249 674144 263566
rect 674286 260944 674342 260953
rect 674286 260879 674342 260888
rect 674300 246945 674328 260879
rect 674286 246936 674342 246945
rect 674286 246871 674342 246880
rect 674102 235240 674158 235249
rect 674102 235175 674158 235184
rect 674196 235000 674248 235006
rect 674484 234977 674512 263566
rect 674196 234942 674248 234948
rect 674470 234968 674526 234977
rect 674208 233238 674236 234942
rect 674470 234903 674526 234912
rect 674380 234796 674432 234802
rect 674380 234738 674432 234744
rect 674196 233232 674248 233238
rect 674196 233174 674248 233180
rect 673840 230438 673960 230466
rect 673840 223689 673868 230438
rect 674392 230330 674420 234738
rect 674668 234433 674696 266999
rect 674838 264480 674894 264489
rect 674838 264415 674894 264424
rect 674852 263809 674880 264415
rect 676494 264072 676550 264081
rect 676494 264007 676550 264016
rect 674838 263800 674894 263809
rect 674838 263735 674894 263744
rect 676508 263673 676536 264007
rect 676494 263664 676550 263673
rect 676494 263599 676550 263608
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259570 676260 262783
rect 675496 259542 676260 259570
rect 675496 252362 675524 259542
rect 675220 252334 675524 252362
rect 674930 251560 674986 251569
rect 674930 251495 674986 251504
rect 674944 251174 674972 251495
rect 674944 251146 675156 251174
rect 674930 249384 674986 249393
rect 674930 249319 674986 249328
rect 674944 245426 674972 249319
rect 675128 247058 675156 251146
rect 675220 247398 675248 252334
rect 678256 252278 678284 263191
rect 678426 261216 678482 261225
rect 678426 261151 678482 261160
rect 675852 252272 675904 252278
rect 675312 252220 675852 252226
rect 675312 252214 675904 252220
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 675312 252198 675892 252214
rect 675312 250526 675340 252198
rect 678440 251598 678468 261151
rect 675852 251592 675904 251598
rect 675850 251560 675852 251569
rect 678428 251592 678480 251598
rect 675904 251560 675906 251569
rect 678428 251534 678480 251540
rect 675850 251495 675906 251504
rect 675312 250498 675418 250526
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249656 675446 249665
rect 675390 249591 675446 249600
rect 675404 249220 675432 249591
rect 675220 247370 675418 247398
rect 675128 247030 675340 247058
rect 675114 246936 675170 246945
rect 675114 246871 675170 246880
rect 675128 246213 675156 246871
rect 675312 246854 675340 247030
rect 675312 246826 675418 246854
rect 675128 246185 675418 246213
rect 675114 245576 675170 245585
rect 675170 245534 675418 245562
rect 675114 245511 675170 245520
rect 674944 245398 675156 245426
rect 674838 245304 674894 245313
rect 674838 245239 674894 245248
rect 674852 241890 674880 245239
rect 675128 243085 675156 245398
rect 675128 243057 675418 243085
rect 675114 242856 675170 242865
rect 675114 242791 675170 242800
rect 675128 242533 675156 242791
rect 675128 242505 675418 242533
rect 674852 241862 675418 241890
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675206 240272 675262 240281
rect 675206 240207 675262 240216
rect 675220 240054 675248 240207
rect 675220 240026 675418 240054
rect 675114 238232 675170 238241
rect 675170 238190 675418 238218
rect 675114 238167 675170 238176
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 675128 237510 675340 237538
rect 675404 237524 675432 237646
rect 675128 235929 675156 237510
rect 675390 236872 675446 236881
rect 675390 236807 675446 236816
rect 675404 236368 675432 236807
rect 675114 235920 675170 235929
rect 675114 235855 675170 235864
rect 675666 235240 675722 235249
rect 675666 235175 675722 235184
rect 674654 234424 674710 234433
rect 674654 234359 674710 234368
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 675680 234274 675708 235175
rect 675850 234968 675906 234977
rect 675850 234903 675906 234912
rect 675864 234598 675892 234903
rect 675852 234592 675904 234598
rect 675852 234534 675904 234540
rect 679624 234592 679676 234598
rect 679624 234534 679676 234540
rect 675850 234424 675906 234433
rect 675850 234359 675852 234368
rect 675904 234359 675906 234368
rect 675852 234330 675904 234336
rect 674564 234252 674616 234258
rect 674564 234194 674616 234200
rect 674576 230602 674604 234194
rect 674898 234104 674926 234262
rect 675680 234258 675892 234274
rect 675680 234252 675904 234258
rect 675680 234246 675852 234252
rect 675852 234194 675904 234200
rect 674760 234076 674926 234104
rect 674760 233102 674788 234076
rect 674944 233986 675892 234002
rect 674932 233980 675904 233986
rect 674984 233974 675852 233980
rect 674932 233922 674984 233928
rect 675852 233922 675904 233928
rect 675236 233708 675288 233714
rect 675236 233650 675288 233656
rect 675248 233594 675276 233650
rect 675248 233578 675892 233594
rect 675248 233572 675904 233578
rect 675248 233566 675852 233572
rect 675852 233514 675904 233520
rect 677784 233572 677836 233578
rect 677784 233514 677836 233520
rect 674748 233096 674800 233102
rect 674748 233038 674800 233044
rect 675496 232626 675892 232642
rect 675484 232620 675892 232626
rect 675536 232614 675892 232620
rect 675484 232562 675536 232568
rect 675864 232558 675892 232614
rect 675852 232552 675904 232558
rect 675852 232494 675904 232500
rect 675346 232348 675398 232354
rect 675346 232290 675398 232296
rect 675358 232082 675386 232290
rect 675346 232076 675398 232082
rect 675346 232018 675398 232024
rect 675178 231840 675234 231849
rect 675178 231775 675180 231784
rect 675232 231775 675234 231784
rect 675180 231746 675232 231752
rect 675070 231532 675122 231538
rect 675070 231474 675122 231480
rect 674956 231328 675008 231334
rect 674954 231296 674956 231305
rect 675008 231296 675010 231305
rect 674954 231231 675010 231240
rect 674840 231192 674892 231198
rect 674838 231160 674840 231169
rect 674892 231160 674894 231169
rect 675082 231146 675110 231474
rect 675850 231296 675906 231305
rect 675850 231231 675852 231240
rect 675904 231231 675906 231240
rect 677600 231260 677652 231266
rect 675852 231202 675904 231208
rect 677600 231202 677652 231208
rect 674838 231095 674894 231104
rect 675036 231118 675110 231146
rect 674732 230920 674784 230926
rect 674730 230888 674732 230897
rect 674784 230888 674786 230897
rect 674730 230823 674786 230832
rect 675036 230625 675064 231118
rect 675022 230616 675078 230625
rect 674576 230574 674696 230602
rect 674518 230512 674570 230518
rect 674518 230454 674570 230460
rect 674530 230353 674558 230454
rect 673932 230302 674420 230330
rect 674516 230344 674572 230353
rect 673932 229786 673960 230302
rect 674516 230279 674572 230288
rect 674104 230240 674156 230246
rect 674668 230194 674696 230574
rect 675022 230551 675078 230560
rect 676770 230344 676826 230353
rect 676770 230279 676826 230288
rect 674156 230188 674696 230194
rect 674104 230182 674696 230188
rect 674116 230166 674696 230182
rect 674288 230104 674340 230110
rect 674056 230072 674112 230081
rect 675114 230072 675170 230081
rect 674340 230052 674604 230058
rect 674288 230046 674604 230052
rect 674300 230030 674604 230046
rect 674056 230007 674112 230016
rect 674070 229906 674098 230007
rect 674172 229968 674224 229974
rect 674576 229922 674604 230030
rect 675170 230042 675892 230058
rect 675170 230036 675904 230042
rect 675170 230030 675852 230036
rect 675114 230007 675170 230016
rect 675852 229978 675904 229984
rect 676588 230036 676640 230042
rect 676588 229978 676640 229984
rect 674224 229916 674512 229922
rect 674172 229910 674512 229916
rect 674058 229900 674110 229906
rect 674184 229894 674512 229910
rect 674576 229906 675892 229922
rect 674576 229900 675904 229906
rect 674576 229894 675852 229900
rect 674058 229842 674110 229848
rect 674484 229786 674512 229894
rect 675852 229842 675904 229848
rect 673932 229758 674144 229786
rect 674484 229770 675892 229786
rect 674484 229764 675904 229770
rect 674484 229758 675852 229764
rect 673948 229560 674000 229566
rect 673932 229508 673948 229514
rect 673932 229502 674000 229508
rect 673932 229486 673988 229502
rect 673932 224954 673960 229486
rect 673932 224926 674052 224954
rect 673826 223680 673882 223689
rect 673826 223615 673882 223624
rect 674024 223394 674052 224926
rect 673932 223366 674052 223394
rect 673932 222873 673960 223366
rect 673918 222864 673974 222873
rect 673918 222799 673974 222808
rect 673656 222166 673960 222194
rect 673564 220782 673776 220810
rect 673748 220697 673776 220782
rect 673734 220688 673790 220697
rect 673734 220623 673790 220632
rect 673472 216294 673592 216322
rect 673366 216200 673422 216209
rect 673366 216135 673422 216144
rect 673104 215266 673224 215294
rect 672722 214704 672778 214713
rect 672722 214639 672778 214648
rect 672906 209944 672962 209953
rect 672906 209879 672962 209888
rect 672552 209746 672672 209774
rect 672644 205634 672672 209746
rect 672644 205606 672764 205634
rect 672446 177848 672502 177857
rect 672446 177783 672502 177792
rect 672538 175264 672594 175273
rect 672538 175199 672594 175208
rect 672354 169144 672410 169153
rect 672354 169079 672410 169088
rect 672368 153105 672396 169079
rect 672354 153096 672410 153105
rect 672354 153031 672410 153040
rect 672078 140312 672134 140321
rect 672078 140247 672134 140256
rect 672552 130529 672580 175199
rect 672736 149161 672764 205606
rect 672722 149152 672778 149161
rect 672722 149087 672778 149096
rect 672538 130520 672594 130529
rect 672538 130455 672594 130464
rect 672354 124400 672410 124409
rect 672354 124335 672410 124344
rect 671894 115832 671950 115841
rect 671894 115767 671950 115776
rect 672368 110265 672396 124335
rect 672920 124001 672948 209879
rect 673104 172961 673132 215266
rect 673380 201929 673408 216135
rect 673564 212945 673592 216294
rect 673550 212936 673606 212945
rect 673550 212871 673606 212880
rect 673932 212534 673960 222166
rect 673748 212506 673960 212534
rect 673550 206952 673606 206961
rect 673550 206887 673606 206896
rect 673366 201920 673422 201929
rect 673366 201855 673422 201864
rect 673564 201657 673592 206887
rect 673550 201648 673606 201657
rect 673550 201583 673606 201592
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 673090 172952 673146 172961
rect 673090 172887 673146 172896
rect 673182 169960 673238 169969
rect 673182 169895 673238 169904
rect 673196 151745 673224 169895
rect 673182 151736 673238 151745
rect 673182 151671 673238 151680
rect 673380 129713 673408 174383
rect 673748 168473 673776 212506
rect 673918 209672 673974 209681
rect 673918 209607 673974 209616
rect 673932 203289 673960 209607
rect 673918 203280 673974 203289
rect 673918 203215 673974 203224
rect 674116 179489 674144 229758
rect 675852 229706 675904 229712
rect 675114 229528 675170 229537
rect 675170 229486 675892 229514
rect 675114 229463 675170 229472
rect 675864 229226 675892 229486
rect 675852 229220 675904 229226
rect 675852 229162 675904 229168
rect 675114 229120 675170 229129
rect 675170 229090 675892 229106
rect 675170 229084 675904 229090
rect 675170 229078 675852 229084
rect 675114 229055 675170 229064
rect 675852 229026 675904 229032
rect 675114 228848 675170 228857
rect 675170 228818 675892 228834
rect 675170 228812 675904 228818
rect 675170 228806 675852 228812
rect 675114 228783 675170 228792
rect 675852 228754 675904 228760
rect 676220 228812 676272 228818
rect 676220 228754 676272 228760
rect 675022 227080 675078 227089
rect 675022 227015 675078 227024
rect 674286 225720 674342 225729
rect 674286 225655 674342 225664
rect 674300 224954 674328 225655
rect 674300 224926 674788 224954
rect 674562 221912 674618 221921
rect 674562 221847 674618 221856
rect 674378 220280 674434 220289
rect 674378 220215 674434 220224
rect 674102 179480 674158 179489
rect 674102 179415 674158 179424
rect 674194 176896 674250 176905
rect 674194 176831 674250 176840
rect 674010 168736 674066 168745
rect 674010 168671 674066 168680
rect 673734 168464 673790 168473
rect 673734 168399 673790 168408
rect 674024 151065 674052 168671
rect 674010 151056 674066 151065
rect 674010 150991 674066 151000
rect 674208 132161 674236 176831
rect 674392 175681 674420 220215
rect 674576 177313 674604 221847
rect 674760 218657 674788 224926
rect 675036 221513 675064 227015
rect 675206 226128 675262 226137
rect 675206 226063 675262 226072
rect 675022 221504 675078 221513
rect 675022 221439 675078 221448
rect 674930 220552 674986 220561
rect 674930 220487 674986 220496
rect 674746 218648 674802 218657
rect 674746 218583 674802 218592
rect 674944 217569 674972 220487
rect 675220 219314 675248 226063
rect 675390 224904 675446 224913
rect 675390 224839 675446 224848
rect 675404 222193 675432 224839
rect 675850 224632 675906 224641
rect 675850 224567 675906 224576
rect 675390 222184 675446 222193
rect 675390 222119 675446 222128
rect 675864 220561 675892 224567
rect 675850 220552 675906 220561
rect 675850 220487 675906 220496
rect 676036 220040 676088 220046
rect 676034 220008 676036 220017
rect 676088 220008 676090 220017
rect 676034 219943 676090 219952
rect 676036 219768 676088 219774
rect 676034 219736 676036 219745
rect 676088 219736 676090 219745
rect 676034 219671 676090 219680
rect 676232 219586 676260 228754
rect 675128 219286 675248 219314
rect 675312 219558 676260 219586
rect 674930 217560 674986 217569
rect 674930 217495 674986 217504
rect 674930 216880 674986 216889
rect 674930 216815 674986 216824
rect 674746 216608 674802 216617
rect 674746 216543 674802 216552
rect 674760 205057 674788 216543
rect 674944 215937 674972 216815
rect 674930 215928 674986 215937
rect 674930 215863 674986 215872
rect 675128 215665 675156 219286
rect 675312 219201 675340 219558
rect 676220 219428 676272 219434
rect 676220 219370 676272 219376
rect 675298 219192 675354 219201
rect 675298 219127 675354 219136
rect 675666 219056 675722 219065
rect 675666 218991 675722 219000
rect 675298 215792 675354 215801
rect 675298 215727 675354 215736
rect 675114 215656 675170 215665
rect 675114 215591 675170 215600
rect 675312 214146 675340 215727
rect 675312 214118 675432 214146
rect 675022 212936 675078 212945
rect 675022 212871 675078 212880
rect 674746 205048 674802 205057
rect 674746 204983 674802 204992
rect 675036 204762 675064 212871
rect 675404 212534 675432 214118
rect 675680 213874 675708 218991
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675852 215144 675904 215150
rect 675850 215112 675852 215121
rect 675904 215112 675906 215121
rect 675850 215047 675906 215056
rect 674852 204734 675064 204762
rect 675128 212506 675432 212534
rect 675496 213846 675708 213874
rect 674852 202745 674880 204734
rect 675128 202874 675156 212506
rect 675496 208298 675524 213846
rect 676048 213602 676076 217767
rect 675680 213574 676076 213602
rect 675680 212945 675708 213574
rect 675850 213480 675906 213489
rect 676232 213466 676260 219370
rect 676600 215294 676628 229978
rect 676784 215294 676812 230279
rect 677232 229900 677284 229906
rect 677232 229842 677284 229848
rect 676956 229764 677008 229770
rect 676956 229706 677008 229712
rect 676968 229242 676996 229706
rect 675906 213438 676260 213466
rect 676324 215266 676628 215294
rect 676692 215266 676812 215294
rect 676876 229214 676996 229242
rect 675850 213415 675906 213424
rect 676324 213330 676352 215266
rect 676140 213302 676352 213330
rect 675852 213240 675904 213246
rect 675850 213208 675852 213217
rect 675904 213208 675906 213217
rect 675850 213143 675906 213152
rect 675666 212936 675722 212945
rect 675666 212871 675722 212880
rect 676140 210338 676168 213302
rect 676692 213246 676720 215266
rect 676680 213240 676732 213246
rect 676680 213182 676732 213188
rect 676140 210310 676260 210338
rect 676232 210066 676260 210310
rect 675312 208270 675524 208298
rect 676140 210038 676260 210066
rect 675312 204049 675340 208270
rect 676140 207233 676168 210038
rect 676876 209681 676904 229214
rect 677048 229084 677100 229090
rect 677048 229026 677100 229032
rect 677060 220046 677088 229026
rect 677048 220040 677100 220046
rect 677048 219982 677100 219988
rect 677244 215150 677272 229842
rect 677416 229084 677468 229090
rect 677416 229026 677468 229032
rect 677428 219774 677456 229026
rect 677416 219768 677468 219774
rect 677416 219710 677468 219716
rect 677612 219434 677640 231202
rect 677600 219428 677652 219434
rect 677600 219370 677652 219376
rect 677232 215144 677284 215150
rect 677232 215086 677284 215092
rect 676862 209672 676918 209681
rect 676862 209607 676918 209616
rect 676126 207224 676182 207233
rect 676126 207159 676182 207168
rect 677796 206961 677824 233514
rect 679254 223816 679310 223825
rect 679254 223751 679310 223760
rect 679268 223582 679296 223751
rect 679256 223576 679308 223582
rect 679256 223518 679308 223524
rect 679636 220697 679664 234534
rect 679992 234388 680044 234394
rect 679992 234330 680044 234336
rect 679808 234252 679860 234258
rect 679808 234194 679860 234200
rect 679820 221513 679848 234194
rect 680004 222329 680032 234330
rect 683854 234152 683910 234161
rect 683854 234087 683910 234096
rect 683488 233980 683540 233986
rect 683488 233922 683540 233928
rect 683302 233880 683358 233889
rect 683302 233815 683358 233824
rect 680176 232552 680228 232558
rect 680176 232494 680228 232500
rect 680188 223582 680216 232494
rect 680176 223576 680228 223582
rect 680176 223518 680228 223524
rect 683316 223145 683344 233815
rect 683302 223136 683358 223145
rect 683302 223071 683358 223080
rect 679990 222320 680046 222329
rect 679990 222255 680046 222264
rect 679806 221504 679862 221513
rect 679806 221439 679862 221448
rect 679622 220688 679678 220697
rect 679622 220623 679678 220632
rect 683500 219881 683528 233922
rect 683868 222737 683896 234087
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683854 222728 683910 222737
rect 683854 222663 683910 222672
rect 683486 219872 683542 219881
rect 683486 219807 683542 219816
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 677782 206952 677838 206961
rect 677782 206887 677838 206896
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675482 205048 675538 205057
rect 675482 204983 675538 204992
rect 675496 204680 675524 204983
rect 675312 204021 675418 204049
rect 675128 202846 675248 202874
rect 674838 202736 674894 202745
rect 674838 202671 674894 202680
rect 675220 201022 675248 202846
rect 675390 202736 675446 202745
rect 675390 202671 675446 202680
rect 675404 202195 675432 202671
rect 675482 201920 675538 201929
rect 675482 201855 675538 201864
rect 675496 201620 675524 201855
rect 675220 200994 675418 201022
rect 675022 200968 675078 200977
rect 675022 200903 675078 200912
rect 675036 194834 675064 200903
rect 675206 200696 675262 200705
rect 675206 200631 675262 200640
rect 675758 200696 675814 200705
rect 675758 200631 675814 200640
rect 675220 196058 675248 200631
rect 675772 200328 675800 200631
rect 675574 198248 675630 198257
rect 675574 198183 675630 198192
rect 675588 197880 675616 198183
rect 675404 197169 675432 197336
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675220 196030 675418 196058
rect 675036 194806 675418 194834
rect 675666 193216 675722 193225
rect 675666 193151 675722 193160
rect 675680 192984 675708 193151
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190369 675340 191950
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675298 190360 675354 190369
rect 675298 190295 675354 190304
rect 683118 186960 683174 186969
rect 683118 186895 683174 186904
rect 676494 181384 676550 181393
rect 676494 181319 676550 181328
rect 676034 178120 676090 178129
rect 676508 178106 676536 181319
rect 683132 178809 683160 186895
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 178800 683174 178809
rect 683118 178735 683174 178744
rect 676090 178078 676536 178106
rect 676034 178055 676090 178064
rect 674562 177304 674618 177313
rect 674562 177239 674618 177248
rect 674654 176080 674710 176089
rect 674654 176015 674710 176024
rect 674378 175672 674434 175681
rect 674378 175607 674434 175616
rect 674378 169552 674434 169561
rect 674378 169487 674434 169496
rect 674392 155417 674420 169487
rect 674378 155408 674434 155417
rect 674378 155343 674434 155352
rect 674194 132152 674250 132161
rect 674194 132087 674250 132096
rect 674668 131345 674696 176015
rect 678242 173224 678298 173233
rect 678242 173159 678298 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674852 157593 674880 172751
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 676048 165617 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162858 678284 173159
rect 681002 171592 681058 171601
rect 681002 171527 681058 171536
rect 679622 171184 679678 171193
rect 679622 171119 679678 171128
rect 676128 162852 676180 162858
rect 676128 162794 676180 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675944 162648 675996 162654
rect 675944 162590 675996 162596
rect 675956 161945 675984 162590
rect 675942 161936 675998 161945
rect 675942 161871 675998 161880
rect 675852 161764 675904 161770
rect 675852 161706 675904 161712
rect 675864 161242 675892 161706
rect 676140 161401 676168 162794
rect 679636 162654 679664 171119
rect 679624 162648 679676 162654
rect 679624 162590 679676 162596
rect 681016 161770 681044 171527
rect 681004 161764 681056 161770
rect 681004 161706 681056 161712
rect 676126 161392 676182 161401
rect 676126 161327 676182 161336
rect 675312 161214 675892 161242
rect 675312 159678 675340 161214
rect 675758 160712 675814 160721
rect 675758 160647 675814 160656
rect 675772 160344 675800 160647
rect 675312 159650 675418 159678
rect 675758 159352 675814 159361
rect 675758 159287 675814 159296
rect 675772 159052 675800 159287
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675390 157040 675446 157049
rect 675390 156975 675446 156984
rect 675404 156643 675432 156975
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675114 155408 675170 155417
rect 675170 155366 675340 155394
rect 675114 155343 675170 155352
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675312 155230 675432 155258
rect 675114 153096 675170 153105
rect 675114 153031 675170 153040
rect 675758 153096 675814 153105
rect 675758 153031 675814 153040
rect 675128 152334 675156 153031
rect 675772 152864 675800 153031
rect 675128 152306 675418 152334
rect 675114 151736 675170 151745
rect 675170 151680 675418 151689
rect 675114 151671 675418 151680
rect 675128 151661 675418 151671
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675666 148472 675722 148481
rect 675666 148407 675722 148416
rect 675680 147968 675708 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675772 146033 675800 146132
rect 675758 146024 675814 146033
rect 675758 145959 675814 145968
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 683132 132705 683160 135895
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 675942 130112 675998 130121
rect 675942 130047 675998 130056
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 674102 129296 674158 129305
rect 674102 129231 674158 129240
rect 673274 126032 673330 126041
rect 673274 125967 673330 125976
rect 672906 123992 672962 124001
rect 672906 123927 672962 123936
rect 673090 123992 673146 124001
rect 673090 123927 673146 123936
rect 672814 123176 672870 123185
rect 672814 123111 672870 123120
rect 672828 121417 672856 123111
rect 672814 121408 672870 121417
rect 672814 121343 672870 121352
rect 673104 121258 673132 123927
rect 673288 123706 673316 125967
rect 672736 121230 673132 121258
rect 673196 123678 673316 123706
rect 672538 121136 672594 121145
rect 672538 121071 672594 121080
rect 672552 110945 672580 121071
rect 672736 117994 672764 121230
rect 673196 118694 673224 123678
rect 673366 123584 673422 123593
rect 673366 123519 673422 123528
rect 673104 118666 673224 118694
rect 672736 117966 672856 117994
rect 672538 110936 672594 110945
rect 672538 110871 672594 110880
rect 672354 110256 672410 110265
rect 672354 110191 672410 110200
rect 671526 107672 671582 107681
rect 671526 107607 671582 107616
rect 672828 106457 672856 117966
rect 673104 111489 673132 118666
rect 673090 111480 673146 111489
rect 673090 111415 673146 111424
rect 672814 106448 672870 106457
rect 672814 106383 672870 106392
rect 670700 106208 670752 106214
rect 670700 106150 670752 106156
rect 673380 105641 673408 123519
rect 674116 111897 674144 129231
rect 675956 128353 675984 130047
rect 674286 128344 674342 128353
rect 674286 128279 674342 128288
rect 675942 128344 675998 128353
rect 675942 128279 675998 128288
rect 674102 111888 674158 111897
rect 674102 111823 674158 111832
rect 673366 105632 673422 105641
rect 673366 105567 673422 105576
rect 668306 104408 668362 104417
rect 668306 104343 668362 104352
rect 668032 100156 668084 100162
rect 668032 100098 668084 100104
rect 668320 92546 668348 104343
rect 674300 102241 674328 128279
rect 682382 127800 682438 127809
rect 682382 127735 682438 127744
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 125624 674710 125633
rect 674654 125559 674710 125568
rect 674470 125216 674526 125225
rect 674470 125151 674526 125160
rect 674484 104666 674512 125151
rect 674668 110786 674696 125559
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 682396 117298 682424 127735
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 682384 117292 682436 117298
rect 682384 117234 682436 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 675114 111480 675170 111489
rect 675170 111438 675418 111466
rect 675114 111415 675170 111424
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 674668 110758 675340 110786
rect 675404 110772 675432 110894
rect 674654 110256 674710 110265
rect 674710 110214 674880 110242
rect 674654 110191 674710 110200
rect 674852 110174 674880 110214
rect 674852 110146 675418 110174
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106457 675156 107086
rect 675114 106448 675170 106457
rect 675114 106383 675170 106392
rect 675772 106185 675800 106488
rect 675758 106176 675814 106185
rect 675758 106111 675814 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 675128 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 105641 675156 105794
rect 675114 105632 675170 105641
rect 675114 105567 675170 105576
rect 674484 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 668490 102232 668546 102241
rect 668490 102167 668546 102176
rect 674286 102232 674342 102241
rect 674286 102167 674342 102176
rect 668504 100026 668532 102167
rect 675680 102136 675708 102575
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668492 100020 668544 100026
rect 668492 99962 668544 99968
rect 668308 92540 668360 92546
rect 668308 92482 668360 92488
rect 666572 84166 666692 84194
rect 664444 62076 664496 62082
rect 664444 62018 664496 62024
rect 663800 58676 663852 58682
rect 663800 58618 663852 58624
rect 663812 47841 663840 58618
rect 666572 57934 666600 84166
rect 666560 57928 666612 57934
rect 666560 57870 666612 57876
rect 663984 55888 664036 55894
rect 663984 55830 664036 55836
rect 663996 48521 664024 55830
rect 663982 48512 664038 48521
rect 663982 48447 664038 48456
rect 663798 47832 663854 47841
rect 663798 47767 663854 47776
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464344 42764 464396 42770
rect 464344 42706 464396 42712
rect 463976 42628 464028 42634
rect 463976 42570 464028 42576
rect 465828 42500 465856 43143
rect 463712 42350 464036 42378
rect 461122 42256 461178 42265
rect 461122 42191 461178 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42364 518848 42735
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40488 141754 40497
rect 141698 40423 141754 40432
rect 141712 39984 141740 40423
<< via2 >>
rect 106830 1007292 106832 1007312
rect 106832 1007292 106884 1007312
rect 106884 1007292 106886 1007312
rect 106830 1007256 106886 1007292
rect 101954 1006596 102010 1006632
rect 101954 1006576 101956 1006596
rect 101956 1006576 102008 1006596
rect 102008 1006576 102010 1006596
rect 84658 995696 84714 995752
rect 85210 995696 85266 995752
rect 86038 995696 86094 995752
rect 90270 995696 90326 995752
rect 88982 995560 89038 995616
rect 89534 995560 89590 995616
rect 77206 995288 77262 995344
rect 80150 995016 80206 995072
rect 81990 994744 82046 994800
rect 86314 994472 86370 994528
rect 92570 997192 92626 997248
rect 92938 996920 92994 996976
rect 92754 996240 92810 996296
rect 93122 994744 93178 994800
rect 93490 995696 93546 995752
rect 87878 994200 87934 994256
rect 104806 1006460 104862 1006496
rect 104806 1006440 104808 1006460
rect 104808 1006440 104860 1006460
rect 104860 1006440 104862 1006460
rect 100298 1006324 100354 1006360
rect 100298 1006304 100300 1006324
rect 100300 1006304 100352 1006324
rect 100352 1006304 100354 1006324
rect 98274 1006052 98330 1006088
rect 98274 1006032 98276 1006052
rect 98276 1006032 98328 1006052
rect 98328 1006032 98330 1006052
rect 95146 994200 95202 994256
rect 81070 993928 81126 993984
rect 94502 993928 94558 993984
rect 42154 967544 42210 967600
rect 42614 967544 42670 967600
rect 41786 967136 41842 967192
rect 42154 967136 42210 967192
rect 42430 964688 42486 964744
rect 42430 963872 42486 963928
rect 42430 963328 42486 963384
rect 42430 963056 42486 963112
rect 41786 962104 41842 962160
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42430 958704 42486 958760
rect 41786 957752 41842 957808
rect 41786 955440 41842 955496
rect 41786 954624 41842 954680
rect 41786 954352 41842 954408
rect 35162 952856 35218 952912
rect 31758 946600 31814 946656
rect 28722 942656 28778 942712
rect 33782 938168 33838 938224
rect 37922 952448 37978 952504
rect 35806 943064 35862 943120
rect 35806 941840 35862 941896
rect 35806 940208 35862 940264
rect 36542 938984 36598 939040
rect 39302 952176 39358 952232
rect 37922 938576 37978 938632
rect 35162 937760 35218 937816
rect 40038 951632 40094 951688
rect 39302 937352 39358 937408
rect 40038 934496 40094 934552
rect 42062 940616 42118 940672
rect 42062 939800 42118 939856
rect 42062 935720 42118 935776
rect 43442 967136 43498 967192
rect 43442 964688 43498 964744
rect 43258 963872 43314 963928
rect 43074 963328 43130 963384
rect 42798 936944 42854 937000
rect 43074 934904 43130 934960
rect 44270 963056 44326 963112
rect 43442 935312 43498 935368
rect 44454 958704 44510 958760
rect 46202 946600 46258 946656
rect 45558 943472 45614 943528
rect 44822 941432 44878 941488
rect 44638 941024 44694 941080
rect 44454 936128 44510 936184
rect 44270 934088 44326 934144
rect 43258 933680 43314 933736
rect 43350 933272 43406 933328
rect 42246 932864 42302 932920
rect 41694 911920 41750 911976
rect 41510 911648 41566 911704
rect 42936 892472 42992 892528
rect 43074 892254 43130 892256
rect 43074 892202 43076 892254
rect 43076 892202 43128 892254
rect 43128 892202 43130 892254
rect 43074 892200 43130 892202
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 35806 817264 35862 817320
rect 35806 816448 35862 816504
rect 35806 814816 35862 814872
rect 42062 884584 42118 884640
rect 41326 812776 41382 812832
rect 40958 812368 41014 812424
rect 35162 811552 35218 811608
rect 35898 811144 35954 811200
rect 40590 808288 40646 808344
rect 40774 805432 40830 805488
rect 41142 811960 41198 812016
rect 41786 809104 41842 809160
rect 42246 806656 42302 806712
rect 41142 805568 41198 805624
rect 40958 805296 41014 805352
rect 40590 805024 40646 805080
rect 41694 802460 41750 802496
rect 41694 802440 41696 802460
rect 41696 802440 41748 802460
rect 41748 802440 41750 802460
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 43166 810736 43222 810792
rect 42798 809920 42854 809976
rect 42522 802440 42578 802496
rect 42522 798904 42578 798960
rect 42154 796184 42210 796240
rect 42522 795368 42578 795424
rect 42062 794960 42118 795016
rect 41786 794144 41842 794200
rect 42246 792512 42302 792568
rect 42982 807472 43038 807528
rect 42154 789248 42210 789304
rect 41786 788568 41842 788624
rect 42246 788160 42302 788216
rect 41786 786800 41842 786856
rect 42706 788976 42762 789032
rect 42706 788568 42762 788624
rect 35806 773472 35862 773528
rect 35622 769392 35678 769448
rect 35438 768984 35494 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 31022 768168 31078 768224
rect 35530 767760 35586 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 37094 763292 37150 763328
rect 37094 763272 37096 763292
rect 37096 763272 37148 763292
rect 37148 763272 37150 763292
rect 41326 765720 41382 765776
rect 40038 764496 40094 764552
rect 36542 757696 36598 757752
rect 40682 758140 40684 758160
rect 40684 758140 40736 758160
rect 40736 758140 40738 758160
rect 40682 758104 40738 758140
rect 42706 765720 42762 765776
rect 39486 757288 39542 757344
rect 41786 756608 41842 756664
rect 42338 754160 42394 754216
rect 41970 754024 42026 754080
rect 42062 752936 42118 752992
rect 42154 751712 42210 751768
rect 42246 750488 42302 750544
rect 41786 750352 41842 750408
rect 41786 747360 41842 747416
rect 42154 746680 42210 746736
rect 42798 757832 42854 757888
rect 42798 750488 42854 750544
rect 42430 745048 42486 745104
rect 42246 744776 42302 744832
rect 41786 743688 41842 743744
rect 42614 743008 42670 743064
rect 42430 741648 42486 741704
rect 35622 731312 35678 731368
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 31022 725192 31078 725248
rect 36542 724784 36598 724840
rect 33046 723968 33102 724024
rect 33782 723152 33838 723208
rect 40682 724376 40738 724432
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41326 720296 41382 720352
rect 40682 714720 40738 714776
rect 41602 715808 41658 715864
rect 41878 715536 41934 715592
rect 42706 715808 42762 715864
rect 42614 715536 42670 715592
rect 41326 714176 41382 714232
rect 42062 714448 42118 714504
rect 41786 713904 41842 713960
rect 41786 713496 41842 713552
rect 42062 713224 42118 713280
rect 41786 712136 41842 712192
rect 42154 710776 42210 710832
rect 42706 711048 42762 711104
rect 41878 709824 41934 709880
rect 42154 708464 42210 708520
rect 42062 707648 42118 707704
rect 41786 707376 41842 707432
rect 42062 706696 42118 706752
rect 42706 708600 42762 708656
rect 42706 707376 42762 707432
rect 42522 706696 42578 706752
rect 42246 706424 42302 706480
rect 42062 703432 42118 703488
rect 42062 702752 42118 702808
rect 42706 702752 42762 702808
rect 42614 702344 42670 702400
rect 41786 700440 41842 700496
rect 42154 699896 42210 699952
rect 41694 697856 41750 697912
rect 35622 691328 35678 691384
rect 35806 687656 35862 687712
rect 35622 687248 35678 687304
rect 35806 683188 35862 683224
rect 35806 683168 35808 683188
rect 35808 683168 35860 683188
rect 35860 683168 35862 683188
rect 35438 682760 35494 682816
rect 35622 682352 35678 682408
rect 35806 681944 35862 682000
rect 35622 681536 35678 681592
rect 35162 680720 35218 680776
rect 35806 681128 35862 681184
rect 41786 680992 41842 681048
rect 39946 677048 40002 677104
rect 40498 672560 40554 672616
rect 42798 679904 42854 679960
rect 42062 673104 42118 673160
rect 42798 672832 42854 672888
rect 42798 672560 42854 672616
rect 41510 672288 41566 672344
rect 42246 672288 42302 672344
rect 37922 671200 37978 671256
rect 42062 668480 42118 668536
rect 42246 668208 42302 668264
rect 41970 667664 42026 667720
rect 42062 666576 42118 666632
rect 42246 664808 42302 664864
rect 41786 663992 41842 664048
rect 42430 663448 42486 663504
rect 42246 662632 42302 662688
rect 42062 659096 42118 659152
rect 42614 659640 42670 659696
rect 42430 658552 42486 658608
rect 42246 658280 42302 658336
rect 42062 657328 42118 657384
rect 42798 659096 42854 659152
rect 42614 657328 42670 657384
rect 35806 646720 35862 646776
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35806 639784 35862 639840
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35806 638560 35862 638616
rect 32402 638152 32458 638208
rect 41786 638152 41842 638208
rect 40038 637336 40094 637392
rect 41786 637540 41842 637596
rect 41418 627680 41474 627736
rect 42062 625776 42118 625832
rect 42522 633800 42578 633856
rect 42706 627680 42762 627736
rect 42522 625776 42578 625832
rect 42522 624960 42578 625016
rect 42246 624008 42302 624064
rect 41970 623328 42026 623384
rect 41786 622104 41842 622160
rect 42430 623328 42486 623384
rect 42522 620064 42578 620120
rect 42706 619792 42762 619848
rect 42430 618840 42486 618896
rect 42430 618432 42486 618488
rect 42062 615848 42118 615904
rect 42430 615440 42486 615496
rect 42062 615168 42118 615224
rect 41878 614080 41934 614136
rect 43166 788160 43222 788216
rect 43166 766264 43222 766320
rect 43166 752936 43222 752992
rect 43166 723560 43222 723616
rect 43166 703432 43222 703488
rect 43166 679088 43222 679144
rect 43166 662632 43222 662688
rect 43166 636248 43222 636304
rect 43166 624008 43222 624064
rect 43534 932048 43590 932104
rect 44086 892764 44142 892800
rect 44086 892744 44088 892764
rect 44088 892744 44140 892764
rect 44140 892744 44142 892764
rect 44086 891948 44142 891984
rect 44086 891928 44088 891948
rect 44088 891928 44140 891948
rect 44140 891928 44142 891948
rect 44454 816040 44510 816096
rect 44270 814408 44326 814464
rect 43902 809512 43958 809568
rect 43718 806248 43774 806304
rect 43902 796184 43958 796240
rect 48962 940072 49018 940128
rect 51722 942248 51778 942304
rect 50342 939800 50398 939856
rect 47582 891928 47638 891984
rect 44638 815632 44694 815688
rect 44822 815224 44878 815280
rect 44638 813592 44694 813648
rect 44454 773200 44510 773256
rect 44454 771976 44510 772032
rect 44270 771568 44326 771624
rect 44270 766672 44326 766728
rect 44270 746680 44326 746736
rect 44270 729680 44326 729736
rect 45006 810328 45062 810384
rect 45190 807880 45246 807936
rect 45190 794960 45246 795016
rect 45006 789248 45062 789304
rect 45098 772792 45154 772848
rect 44822 772384 44878 772440
rect 44730 771160 44786 771216
rect 44454 729272 44510 729328
rect 44178 722744 44234 722800
rect 43902 721520 43958 721576
rect 43902 711048 43958 711104
rect 44178 707648 44234 707704
rect 44546 728864 44602 728920
rect 44362 686840 44418 686896
rect 44362 686432 44418 686488
rect 44914 770752 44970 770808
rect 44914 770344 44970 770400
rect 44730 728456 44786 728512
rect 44730 728048 44786 728104
rect 45282 764768 45338 764824
rect 45558 764224 45614 764280
rect 45282 753480 45338 753536
rect 45098 730088 45154 730144
rect 44914 727640 44970 727696
rect 45098 727232 45154 727288
rect 44730 721112 44786 721168
rect 44546 686024 44602 686080
rect 44178 680312 44234 680368
rect 44362 679496 44418 679552
rect 44362 664808 44418 664864
rect 44178 663448 44234 663504
rect 44914 685208 44970 685264
rect 45374 685616 45430 685672
rect 45282 684800 45338 684856
rect 45098 684392 45154 684448
rect 44914 683984 44970 684040
rect 44730 653112 44786 653168
rect 44546 643592 44602 643648
rect 44730 643320 44786 643376
rect 44454 642504 44510 642560
rect 43902 635296 43958 635352
rect 44270 633392 44326 633448
rect 43902 623328 43958 623384
rect 43994 614080 44050 614136
rect 42982 612312 43038 612368
rect 43580 612332 43636 612368
rect 43580 612312 43582 612332
rect 43582 612312 43634 612332
rect 43634 612312 43636 612332
rect 42706 610952 42762 611008
rect 45374 643048 45430 643104
rect 45190 642232 45246 642288
rect 44914 641416 44970 641472
rect 45006 641144 45062 641200
rect 45374 640872 45430 640928
rect 45190 636520 45246 636576
rect 44914 635704 44970 635760
rect 44914 620064 44970 620120
rect 44822 610972 44878 611008
rect 44822 610952 44824 610972
rect 44824 610952 44876 610972
rect 44876 610952 44878 610972
rect 44730 600480 44786 600536
rect 44914 600072 44970 600128
rect 44454 599664 44510 599720
rect 44730 599256 44786 599312
rect 42982 596944 43038 597000
rect 41050 596808 41106 596864
rect 32402 595584 32458 595640
rect 36542 595176 36598 595232
rect 35162 594360 35218 594416
rect 37922 594768 37978 594824
rect 40682 593544 40738 593600
rect 39946 590688 40002 590744
rect 37922 585112 37978 585168
rect 40498 589600 40554 589656
rect 39946 584840 40002 584896
rect 41234 595992 41290 596048
rect 41326 593952 41382 594008
rect 41878 592728 41934 592784
rect 41694 586064 41750 586120
rect 41878 585792 41934 585848
rect 41510 585384 41566 585440
rect 40682 584568 40738 584624
rect 42522 586064 42578 586120
rect 42430 585792 42486 585848
rect 42154 584840 42210 584896
rect 42246 581440 42302 581496
rect 42246 580760 42302 580816
rect 41786 580216 41842 580272
rect 42430 580488 42486 580544
rect 41786 578176 41842 578232
rect 41786 577496 41842 577552
rect 42430 577360 42486 577416
rect 42246 576816 42302 576872
rect 42154 573824 42210 573880
rect 42706 573824 42762 573880
rect 42062 572600 42118 572656
rect 42246 572192 42302 572248
rect 42062 570968 42118 571024
rect 42614 571920 42670 571976
rect 42338 569200 42394 569256
rect 35806 558048 35862 558104
rect 42062 558456 42118 558512
rect 42062 557504 42118 557560
rect 44454 591912 44510 591968
rect 43442 590280 43498 590336
rect 35806 554804 35862 554840
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35622 553968 35678 554024
rect 35806 553580 35862 553616
rect 35806 553560 35808 553580
rect 35808 553560 35860 553580
rect 35860 553560 35862 553580
rect 40958 553352 41014 553408
rect 33782 551928 33838 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41694 553016 41750 553072
rect 41142 552744 41198 552800
rect 41326 552336 41382 552392
rect 41786 552064 41842 552120
rect 41694 551792 41750 551848
rect 41326 551112 41382 551168
rect 41786 550568 41842 550624
rect 42062 550160 42118 550216
rect 41326 548256 41382 548312
rect 41326 546352 41382 546408
rect 41786 549888 41842 549944
rect 41694 547712 41750 547768
rect 42062 545672 42118 545728
rect 41510 545400 41566 545456
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42982 552064 43038 552120
rect 42798 550568 42854 550624
rect 42614 540232 42670 540288
rect 42522 537512 42578 537568
rect 41786 536968 41842 537024
rect 42154 536968 42210 537024
rect 41786 535200 41842 535256
rect 42154 533840 42210 533896
rect 42246 533160 42302 533216
rect 42522 532752 42578 532808
rect 43166 549480 43222 549536
rect 42982 533840 43038 533896
rect 43166 533160 43222 533216
rect 42154 530032 42210 530088
rect 41878 529352 41934 529408
rect 42522 530576 42578 530632
rect 42706 530032 42762 530088
rect 42614 529624 42670 529680
rect 42890 529080 42946 529136
rect 41326 425992 41382 426048
rect 40958 425584 41014 425640
rect 36542 424360 36598 424416
rect 41326 423952 41382 424008
rect 41142 418784 41198 418840
rect 41970 422728 42026 422784
rect 41786 421912 41842 421968
rect 42430 419872 42486 419928
rect 41970 418512 42026 418568
rect 41786 418240 41842 418296
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42430 406952 42486 407008
rect 41786 406272 41842 406328
rect 42614 405592 42670 405648
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 42430 399744 42486 399800
rect 43074 423136 43130 423192
rect 43258 421096 43314 421152
rect 43258 407768 43314 407824
rect 43074 402872 43130 402928
rect 41786 398792 41842 398848
rect 41142 387116 41198 387152
rect 41142 387096 41144 387116
rect 41144 387096 41196 387116
rect 41196 387096 41198 387116
rect 41878 386960 41934 387016
rect 41326 386688 41382 386744
rect 41510 386688 41566 386744
rect 41326 382608 41382 382664
rect 40038 382200 40094 382256
rect 37922 381384 37978 381440
rect 33782 380160 33838 380216
rect 28538 376488 28594 376544
rect 28538 373224 28594 373280
rect 35806 379344 35862 379400
rect 35806 376080 35862 376136
rect 40222 380976 40278 381032
rect 40038 376896 40094 376952
rect 41694 375420 41750 375456
rect 41694 375400 41696 375420
rect 41696 375400 41748 375420
rect 41748 375400 41750 375420
rect 41694 373260 41696 373280
rect 41696 373260 41748 373280
rect 41748 373260 41750 373280
rect 41694 373224 41750 373260
rect 33782 371864 33838 371920
rect 41786 368464 41842 368520
rect 42614 373224 42670 373280
rect 42430 366968 42486 367024
rect 42338 365744 42394 365800
rect 42154 364928 42210 364984
rect 44454 581032 44510 581088
rect 45282 625232 45338 625288
rect 45098 598848 45154 598904
rect 45098 598440 45154 598496
rect 44914 557232 44970 557288
rect 44730 556416 44786 556472
rect 44638 556008 44694 556064
rect 44362 554376 44418 554432
rect 44178 549072 44234 549128
rect 43626 547712 43682 547768
rect 43810 547032 43866 547088
rect 43350 375400 43406 375456
rect 42798 365744 42854 365800
rect 42430 364248 42486 364304
rect 41786 363568 41842 363624
rect 41786 360032 41842 360088
rect 41786 359352 41842 359408
rect 41786 358672 41842 358728
rect 42430 357312 42486 357368
rect 42062 356904 42118 356960
rect 42430 356088 42486 356144
rect 43350 355816 43406 355872
rect 41878 355680 41934 355736
rect 44178 537512 44234 537568
rect 44178 428440 44234 428496
rect 43994 419464 44050 419520
rect 46386 763000 46442 763056
rect 46202 756336 46258 756392
rect 45742 676640 45798 676696
rect 46018 637744 46074 637800
rect 46202 637064 46258 637120
rect 46202 618432 46258 618488
rect 46018 615576 46074 615632
rect 46938 719888 46994 719944
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47582 712136 47638 712192
rect 47214 677864 47270 677920
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 97446 997192 97502 997248
rect 100298 1002516 100354 1002552
rect 100298 1002496 100300 1002516
rect 100300 1002496 100352 1002516
rect 100352 1002496 100354 1002516
rect 99102 1002380 99158 1002416
rect 99102 1002360 99104 1002380
rect 99104 1002360 99156 1002380
rect 99156 1002360 99158 1002380
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 99470 1002108 99526 1002144
rect 99470 1002088 99472 1002108
rect 99472 1002088 99524 1002108
rect 99524 1002088 99526 1002108
rect 101126 1001972 101182 1002008
rect 101126 1001952 101128 1001972
rect 101128 1001952 101180 1001972
rect 101180 1001952 101182 1001972
rect 98826 995832 98882 995888
rect 103978 1006188 104034 1006224
rect 103978 1006168 103980 1006188
rect 103980 1006168 104032 1006188
rect 104032 1006168 104034 1006188
rect 106002 1006188 106058 1006224
rect 106002 1006168 106004 1006188
rect 106004 1006168 106056 1006188
rect 106056 1006168 106058 1006188
rect 102322 1006052 102378 1006088
rect 102322 1006032 102324 1006052
rect 102324 1006032 102376 1006052
rect 102376 1006032 102378 1006052
rect 108486 1006052 108542 1006088
rect 108486 1006032 108488 1006052
rect 108488 1006032 108540 1006052
rect 108540 1006032 108542 1006052
rect 108854 1005252 108856 1005272
rect 108856 1005252 108908 1005272
rect 108908 1005252 108910 1005272
rect 101954 1002652 102010 1002688
rect 101954 1002632 101956 1002652
rect 101956 1002632 102008 1002652
rect 102008 1002632 102010 1002652
rect 101402 995288 101458 995344
rect 97262 994472 97318 994528
rect 108854 1005216 108910 1005252
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 103150 1003892 103152 1003912
rect 103152 1003892 103204 1003912
rect 103204 1003892 103206 1003912
rect 103150 1003856 103206 1003892
rect 105634 1002244 105690 1002280
rect 105634 1002224 105636 1002244
rect 105636 1002224 105688 1002244
rect 105688 1002224 105690 1002244
rect 103150 1002108 103206 1002144
rect 103150 1002088 103152 1002108
rect 103152 1002088 103204 1002108
rect 103204 1002088 103206 1002108
rect 104806 1001952 104862 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 107658 1002380 107714 1002416
rect 107658 1002360 107660 1002380
rect 107660 1002360 107712 1002380
rect 107712 1002360 107714 1002380
rect 108026 1002244 108082 1002280
rect 108026 1002224 108028 1002244
rect 108028 1002224 108080 1002244
rect 108080 1002224 108082 1002244
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 425518 1007140 425574 1007176
rect 425518 1007120 425520 1007140
rect 425520 1007120 425572 1007140
rect 425572 1007120 425574 1007140
rect 359738 1007004 359794 1007040
rect 359738 1006984 359740 1007004
rect 359740 1006984 359792 1007004
rect 359792 1006984 359794 1007004
rect 359370 1006868 359426 1006904
rect 359370 1006848 359372 1006868
rect 359372 1006848 359424 1006868
rect 359424 1006848 359426 1006868
rect 361394 1006732 361450 1006768
rect 361394 1006712 361396 1006732
rect 361396 1006712 361448 1006732
rect 361448 1006712 361450 1006732
rect 153750 1006596 153806 1006632
rect 153750 1006576 153752 1006596
rect 153752 1006576 153804 1006596
rect 153804 1006576 153806 1006596
rect 157430 1006596 157486 1006632
rect 157430 1006576 157432 1006596
rect 157432 1006576 157484 1006596
rect 157484 1006576 157486 1006596
rect 117134 997192 117190 997248
rect 116122 996920 116178 996976
rect 143814 997192 143870 997248
rect 126242 996240 126298 996296
rect 131854 995696 131910 995752
rect 132958 995696 133014 995752
rect 136730 995696 136786 995752
rect 140410 995696 140466 995752
rect 141790 995560 141846 995616
rect 124862 995016 124918 995072
rect 132406 995288 132462 995344
rect 132130 994744 132186 994800
rect 137374 995424 137430 995480
rect 135902 994336 135958 994392
rect 133142 994064 133198 994120
rect 137558 993828 137560 993848
rect 137560 993828 137612 993848
rect 137612 993828 137614 993848
rect 137558 993792 137614 993828
rect 139214 994064 139270 994120
rect 137742 993656 137798 993712
rect 139398 993928 139454 993984
rect 142158 994472 142214 994528
rect 141974 994336 142030 994392
rect 142158 994200 142214 994256
rect 142158 993656 142214 993712
rect 142342 993656 142398 993712
rect 144826 996920 144882 996976
rect 144642 996648 144698 996704
rect 144550 996240 144606 996296
rect 144274 995832 144330 995888
rect 152922 1006460 152978 1006496
rect 152922 1006440 152924 1006460
rect 152924 1006440 152976 1006460
rect 152976 1006440 152978 1006460
rect 158258 1006460 158314 1006496
rect 158258 1006440 158260 1006460
rect 158260 1006440 158312 1006460
rect 158312 1006440 158314 1006460
rect 145562 994744 145618 994800
rect 158626 1006324 158682 1006360
rect 158626 1006304 158628 1006324
rect 158628 1006304 158680 1006324
rect 158680 1006304 158682 1006324
rect 151266 1006188 151322 1006224
rect 151266 1006168 151268 1006188
rect 151268 1006168 151320 1006188
rect 151320 1006168 151322 1006188
rect 152094 1006188 152150 1006224
rect 152094 1006168 152096 1006188
rect 152096 1006168 152148 1006188
rect 152148 1006168 152150 1006188
rect 160282 1006188 160338 1006224
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 147126 1006032 147182 1006088
rect 148874 1006052 148930 1006088
rect 148874 1006032 148876 1006052
rect 148876 1006032 148928 1006052
rect 148928 1006032 148930 1006052
rect 145746 993928 145802 993984
rect 139214 993384 139270 993440
rect 143814 993384 143870 993440
rect 150070 1006052 150126 1006088
rect 150070 1006032 150072 1006052
rect 150072 1006032 150124 1006052
rect 150124 1006032 150126 1006052
rect 158258 1006052 158314 1006088
rect 158258 1006032 158260 1006052
rect 158260 1006032 158312 1006052
rect 158312 1006032 158314 1006052
rect 159454 1006052 159510 1006088
rect 159454 1006032 159456 1006052
rect 159456 1006032 159508 1006052
rect 159508 1006032 159510 1006052
rect 152922 1005100 152978 1005136
rect 152922 1005080 152924 1005100
rect 152924 1005080 152976 1005100
rect 152976 1005080 152978 1005100
rect 147126 995560 147182 995616
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 153750 1004964 153806 1005000
rect 153750 1004944 153752 1004964
rect 153752 1004944 153804 1004964
rect 153804 1004944 153806 1004964
rect 150898 1002380 150954 1002416
rect 150898 1002360 150900 1002380
rect 150900 1002360 150952 1002380
rect 150952 1002360 150954 1002380
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 148506 994200 148562 994256
rect 151726 1004828 151782 1004864
rect 151726 1004808 151728 1004828
rect 151728 1004808 151780 1004828
rect 151780 1004808 151782 1004828
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 154118 1004692 154174 1004728
rect 154118 1004672 154120 1004692
rect 154120 1004672 154172 1004692
rect 154172 1004672 154174 1004692
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 154578 1002108 154634 1002144
rect 154578 1002088 154580 1002108
rect 154580 1002088 154632 1002108
rect 154632 1002088 154634 1002108
rect 154302 995696 154358 995752
rect 154302 995016 154358 995072
rect 154946 1001952 155002 1002008
rect 155774 1001952 155830 1002008
rect 156602 1001972 156658 1002008
rect 156602 1001952 156604 1001972
rect 156604 1001952 156656 1001972
rect 156656 1001952 156658 1001972
rect 157798 1002108 157854 1002144
rect 157798 1002088 157800 1002108
rect 157800 1002088 157852 1002108
rect 157852 1002088 157854 1002108
rect 154578 994472 154634 994528
rect 152462 993656 152518 993712
rect 171046 995152 171102 995208
rect 171506 995165 171508 995208
rect 171508 995165 171560 995208
rect 171560 995165 171562 995208
rect 171506 995152 171562 995165
rect 256146 1006460 256202 1006496
rect 256146 1006440 256148 1006460
rect 256148 1006440 256200 1006460
rect 256200 1006440 256202 1006460
rect 307758 1006460 307814 1006496
rect 307758 1006440 307760 1006460
rect 307760 1006440 307812 1006460
rect 307812 1006440 307814 1006460
rect 360566 1006460 360622 1006496
rect 360566 1006440 360568 1006460
rect 360568 1006440 360620 1006460
rect 360620 1006440 360622 1006460
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 208398 1006052 208454 1006088
rect 208398 1006032 208400 1006052
rect 208400 1006032 208452 1006052
rect 208452 1006032 208454 1006052
rect 175922 995968 175978 996024
rect 195150 997056 195206 997112
rect 195058 996784 195114 996840
rect 188066 995696 188122 995752
rect 189446 995696 189502 995752
rect 191746 995696 191802 995752
rect 192482 995696 192538 995752
rect 192298 995560 192354 995616
rect 194322 995560 194378 995616
rect 195058 995560 195114 995616
rect 177302 995288 177358 995344
rect 173162 995016 173218 995072
rect 184846 994744 184902 994800
rect 186134 994356 186190 994392
rect 186134 994336 186136 994356
rect 186136 994336 186188 994356
rect 186188 994336 186190 994356
rect 186502 994336 186558 994392
rect 184294 993964 184296 993984
rect 184296 993964 184348 993984
rect 184348 993964 184350 993984
rect 184294 993928 184350 993964
rect 186272 993964 186274 993984
rect 186274 993964 186326 993984
rect 186326 993964 186328 993984
rect 186272 993928 186328 993964
rect 188802 994472 188858 994528
rect 187422 993812 187478 993848
rect 187422 993792 187424 993812
rect 187424 993792 187476 993812
rect 187476 993792 187478 993812
rect 195702 996104 195758 996160
rect 195518 995288 195574 995344
rect 195518 994744 195574 994800
rect 195242 993792 195298 993848
rect 196622 994200 196678 994256
rect 212078 1005252 212080 1005272
rect 212080 1005252 212132 1005272
rect 212132 1005252 212134 1005272
rect 202694 1001972 202750 1002008
rect 202694 1001952 202696 1001972
rect 202696 1001952 202748 1001972
rect 202748 1001952 202750 1001972
rect 200670 997908 200672 997928
rect 200672 997908 200724 997928
rect 200724 997908 200726 997928
rect 200670 997872 200726 997908
rect 198738 997736 198794 997792
rect 200026 997736 200082 997792
rect 202694 998180 202696 998200
rect 202696 998180 202748 998200
rect 202748 998180 202750 998200
rect 202694 998144 202750 998180
rect 201866 998044 201868 998064
rect 201868 998044 201920 998064
rect 201920 998044 201922 998064
rect 201866 998008 201922 998044
rect 198738 997056 198794 997112
rect 200210 996820 200212 996840
rect 200212 996820 200264 996840
rect 200264 996820 200266 996840
rect 200210 996784 200266 996820
rect 198186 996376 198242 996432
rect 203522 998572 203578 998608
rect 203522 998552 203524 998572
rect 203524 998552 203576 998572
rect 203576 998552 203578 998572
rect 203522 998316 203524 998336
rect 203524 998316 203576 998336
rect 203576 998316 203578 998336
rect 203522 998280 203578 998316
rect 202970 995868 202972 995888
rect 202972 995868 203024 995888
rect 203024 995868 203026 995888
rect 202970 995832 203026 995868
rect 203154 995832 203210 995888
rect 203154 995288 203210 995344
rect 200762 994472 200818 994528
rect 203890 1001172 203892 1001192
rect 203892 1001172 203944 1001192
rect 203944 1001172 203946 1001192
rect 203890 1001136 203946 1001172
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 204718 997908 204720 997928
rect 204720 997908 204772 997928
rect 204772 997908 204774 997928
rect 204718 997872 204774 997908
rect 212078 1005216 212134 1005252
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 211250 1004828 211306 1004864
rect 211250 1004808 211252 1004828
rect 211252 1004808 211304 1004828
rect 211304 1004808 211306 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002244 206430 1002280
rect 206374 1002224 206376 1002244
rect 206376 1002224 206428 1002244
rect 206428 1002224 206430 1002244
rect 206742 1002244 206798 1002280
rect 206742 1002224 206744 1002244
rect 206744 1002224 206796 1002244
rect 206796 1002224 206798 1002244
rect 207202 1002108 207258 1002144
rect 207202 1002088 207204 1002108
rect 207204 1002088 207256 1002108
rect 207256 1002088 207258 1002108
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 205546 998044 205548 998064
rect 205548 998044 205600 998064
rect 205600 998044 205602 998064
rect 205546 998008 205602 998044
rect 206742 1001952 206798 1002008
rect 207570 1001952 207626 1002008
rect 208398 995832 208454 995888
rect 210882 1002108 210938 1002144
rect 210882 1002088 210884 1002108
rect 210884 1002088 210936 1002108
rect 210936 1002088 210938 1002108
rect 212538 1001972 212594 1002008
rect 212538 1001952 212540 1001972
rect 212540 1001952 212592 1001972
rect 212592 1001952 212594 1001972
rect 208398 995016 208454 995072
rect 234526 995696 234582 995752
rect 238574 995696 238630 995752
rect 240046 995696 240102 995752
rect 243450 995696 243506 995752
rect 243818 995696 243874 995752
rect 244094 995696 244150 995752
rect 240874 995560 240930 995616
rect 243266 995560 243322 995616
rect 241886 995288 241942 995344
rect 242070 995288 242126 995344
rect 235906 995016 235962 995072
rect 239586 995016 239642 995072
rect 235262 994744 235318 994800
rect 246946 996920 247002 996976
rect 246762 995696 246818 995752
rect 247498 997192 247554 997248
rect 247314 995968 247370 996024
rect 246486 995016 246542 995072
rect 246670 995016 246726 995072
rect 241886 994472 241942 994528
rect 258998 1006324 259054 1006360
rect 258998 1006304 259000 1006324
rect 259000 1006304 259052 1006324
rect 259052 1006304 259054 1006324
rect 252466 1006032 252522 1006088
rect 249062 997192 249118 997248
rect 248050 996648 248106 996704
rect 247866 994472 247922 994528
rect 255318 1003892 255320 1003912
rect 255320 1003892 255372 1003912
rect 255372 1003892 255374 1003912
rect 255318 1003856 255374 1003892
rect 252466 997772 252468 997792
rect 252468 997772 252520 997792
rect 252520 997772 252522 997792
rect 252466 997736 252522 997772
rect 250626 995016 250682 995072
rect 254122 1002532 254124 1002552
rect 254124 1002532 254176 1002552
rect 254176 1002532 254178 1002552
rect 254122 1002496 254178 1002532
rect 254490 1002380 254546 1002416
rect 254490 1002360 254492 1002380
rect 254492 1002360 254544 1002380
rect 254544 1002360 254546 1002380
rect 253662 998164 253718 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 253662 997908 253664 997928
rect 253664 997908 253716 997928
rect 253716 997908 253718 997928
rect 253662 997872 253718 997908
rect 253386 995288 253442 995344
rect 255318 1002108 255374 1002144
rect 255318 1002088 255320 1002108
rect 255320 1002088 255372 1002108
rect 255372 1002088 255374 1002108
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 257342 1006052 257398 1006088
rect 257342 1006032 257344 1006052
rect 257344 1006032 257396 1006052
rect 257396 1006032 257398 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 256146 1002668 256148 1002688
rect 256148 1002668 256200 1002688
rect 256200 1002668 256202 1002688
rect 256146 1002632 256202 1002668
rect 256514 1002244 256570 1002280
rect 256514 1002224 256516 1002244
rect 256516 1002224 256568 1002244
rect 256568 1002224 256570 1002244
rect 256974 1001972 257030 1002008
rect 256974 1001952 256976 1001972
rect 256976 1001952 257028 1001972
rect 257028 1001952 257030 1001972
rect 258170 1005080 258226 1005136
rect 263046 1004964 263102 1005000
rect 263046 1004944 263048 1004964
rect 263048 1004944 263100 1004964
rect 263100 1004944 263102 1004964
rect 258170 1004828 258226 1004864
rect 258170 1004808 258172 1004828
rect 258172 1004808 258224 1004828
rect 258224 1004808 258226 1004828
rect 253110 994744 253166 994800
rect 258998 1001952 259054 1002008
rect 261022 1002516 261078 1002552
rect 261022 1002496 261024 1002516
rect 261024 1002496 261076 1002516
rect 261076 1002496 261078 1002516
rect 260194 1002380 260250 1002416
rect 260194 1002360 260196 1002380
rect 260196 1002360 260248 1002380
rect 260248 1002360 260250 1002380
rect 259826 1002244 259882 1002280
rect 259826 1002224 259828 1002244
rect 259828 1002224 259880 1002244
rect 259880 1002224 259882 1002244
rect 261022 1002108 261078 1002144
rect 261022 1002088 261024 1002108
rect 261024 1002088 261076 1002108
rect 261076 1002088 261078 1002108
rect 260194 1001972 260250 1002008
rect 260194 1001952 260196 1001972
rect 260196 1001952 260248 1001972
rect 260248 1001952 260250 1001972
rect 261850 1001952 261906 1002008
rect 263506 1002108 263562 1002144
rect 263506 1002088 263508 1002108
rect 263508 1002088 263560 1002108
rect 263560 1002088 263562 1002108
rect 263874 1001972 263930 1002008
rect 263874 1001952 263876 1001972
rect 263876 1001952 263928 1001972
rect 263928 1001952 263930 1001972
rect 270406 995016 270462 995072
rect 298098 998824 298154 998880
rect 298098 995968 298154 996024
rect 298650 997736 298706 997792
rect 298466 996376 298522 996432
rect 282734 995696 282790 995752
rect 286782 995696 286838 995752
rect 293590 995696 293646 995752
rect 295338 995696 295394 995752
rect 297270 995696 297326 995752
rect 298282 995696 298338 995752
rect 293222 995560 293278 995616
rect 295522 995560 295578 995616
rect 296902 995560 296958 995616
rect 279422 995288 279478 995344
rect 285954 994472 286010 994528
rect 287794 994744 287850 994800
rect 291474 994744 291530 994800
rect 298466 995560 298522 995616
rect 287150 994200 287206 994256
rect 292118 994200 292174 994256
rect 299386 1002224 299442 1002280
rect 299202 996920 299258 996976
rect 300490 998824 300546 998880
rect 306930 1006324 306986 1006360
rect 306930 1006304 306932 1006324
rect 306932 1006304 306984 1006324
rect 306984 1006304 306986 1006324
rect 314658 1006324 314714 1006360
rect 314658 1006304 314660 1006324
rect 314660 1006304 314712 1006324
rect 314712 1006304 314714 1006324
rect 304906 1006188 304962 1006224
rect 304906 1006168 304908 1006188
rect 304908 1006168 304960 1006188
rect 304960 1006168 304962 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006052 311862 1006088
rect 311806 1006032 311808 1006052
rect 311808 1006032 311860 1006052
rect 311860 1006032 311862 1006052
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 307298 1005236 307354 1005272
rect 307298 1005216 307300 1005236
rect 307300 1005216 307352 1005236
rect 307352 1005216 307354 1005236
rect 301686 997736 301742 997792
rect 303250 1002244 303306 1002280
rect 303250 1002224 303252 1002244
rect 303252 1002224 303304 1002244
rect 303304 1002224 303306 1002244
rect 304078 1002108 304134 1002144
rect 304078 1002088 304080 1002108
rect 304080 1002088 304132 1002108
rect 304132 1002088 304134 1002108
rect 302882 997192 302938 997248
rect 302238 996648 302294 996704
rect 301502 995560 301558 995616
rect 308954 1005100 309010 1005136
rect 308954 1005080 308956 1005100
rect 308956 1005080 309008 1005100
rect 309008 1005080 309010 1005100
rect 305274 1003332 305330 1003368
rect 305274 1003312 305276 1003332
rect 305276 1003312 305328 1003332
rect 305328 1003312 305330 1003332
rect 308126 1004828 308182 1004864
rect 308126 1004808 308128 1004828
rect 308128 1004808 308180 1004828
rect 308180 1004808 308182 1004828
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 306930 1004692 306986 1004728
rect 306930 1004672 306932 1004692
rect 306932 1004672 306984 1004692
rect 306984 1004672 306986 1004692
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 310610 1002496 310666 1002552
rect 306102 1002244 306158 1002280
rect 306102 1002224 306104 1002244
rect 306104 1002224 306156 1002244
rect 306156 1002224 306158 1002244
rect 306102 1001972 306158 1002008
rect 306102 1001952 306104 1001972
rect 306104 1001952 306156 1001972
rect 306156 1001952 306158 1001972
rect 308954 1001972 309010 1002008
rect 308954 1001952 308956 1001972
rect 308956 1001952 309008 1001972
rect 309008 1001952 309010 1001972
rect 308770 995560 308826 995616
rect 308770 995016 308826 995072
rect 309782 1001952 309838 1002008
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 310610 1002244 310666 1002280
rect 310610 1002224 310612 1002244
rect 310612 1002224 310664 1002244
rect 310664 1002224 310666 1002244
rect 309138 994744 309194 994800
rect 304262 994472 304318 994528
rect 300306 994200 300362 994256
rect 357714 1006188 357770 1006224
rect 357714 1006168 357716 1006188
rect 357716 1006168 357768 1006188
rect 357768 1006168 357770 1006188
rect 354862 1006032 354918 1006088
rect 355690 1006052 355746 1006088
rect 355690 1006032 355692 1006052
rect 355692 1006032 355744 1006052
rect 355744 1006032 355746 1006052
rect 356518 1005252 356520 1005272
rect 356520 1005252 356572 1005272
rect 356572 1005252 356574 1005272
rect 356518 1005216 356574 1005252
rect 355690 1004964 355746 1005000
rect 355690 1004944 355692 1004964
rect 355692 1004944 355744 1004964
rect 355744 1004944 355746 1004964
rect 356518 1004828 356574 1004864
rect 356518 1004808 356520 1004828
rect 356520 1004808 356572 1004828
rect 356572 1004808 356574 1004828
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 358542 1002244 358598 1002280
rect 358542 1002224 358544 1002244
rect 358544 1002224 358596 1002244
rect 358596 1002224 358598 1002244
rect 357714 1002108 357770 1002144
rect 357714 1002088 357716 1002108
rect 357716 1002088 357768 1002108
rect 357768 1002088 357770 1002108
rect 356886 1001952 356942 1002008
rect 358542 1001952 358598 1002008
rect 360566 1005388 360568 1005408
rect 360568 1005388 360620 1005408
rect 360620 1005388 360622 1005408
rect 360566 1005352 360622 1005388
rect 360198 1001972 360254 1002008
rect 360198 1001952 360200 1001972
rect 360200 1001952 360252 1001972
rect 360252 1001952 360254 1001972
rect 359462 995832 359518 995888
rect 365074 1006188 365130 1006224
rect 365074 1006168 365076 1006188
rect 365076 1006168 365128 1006188
rect 365128 1006168 365130 1006188
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 363418 1006052 363474 1006088
rect 363418 1006032 363420 1006052
rect 363420 1006032 363472 1006052
rect 363472 1006032 363474 1006052
rect 365074 1005100 365130 1005136
rect 365074 1005080 365076 1005100
rect 365076 1005080 365128 1005100
rect 365128 1005080 365130 1005100
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 428370 1006884 428372 1006904
rect 428372 1006884 428424 1006904
rect 428424 1006884 428426 1006904
rect 428370 1006848 428426 1006884
rect 507858 1006884 507860 1006904
rect 507860 1006884 507912 1006904
rect 507912 1006884 507914 1006904
rect 507858 1006848 507914 1006884
rect 429198 1006748 429200 1006768
rect 429200 1006748 429252 1006768
rect 429252 1006748 429254 1006768
rect 429198 1006712 429254 1006748
rect 372526 996920 372582 996976
rect 372342 996648 372398 996704
rect 373262 995968 373318 996024
rect 431682 1006612 431684 1006632
rect 431684 1006612 431736 1006632
rect 431736 1006612 431738 1006632
rect 431682 1006576 431738 1006612
rect 429198 1006460 429254 1006496
rect 429198 1006440 429200 1006460
rect 429200 1006440 429252 1006460
rect 429252 1006440 429254 1006460
rect 376022 998280 376078 998336
rect 381542 996240 381598 996296
rect 380898 995968 380954 996024
rect 382278 995696 382334 995752
rect 383474 995424 383530 995480
rect 399942 996920 399998 996976
rect 388718 995696 388774 995752
rect 385406 994982 385462 995038
rect 385958 994880 386014 994936
rect 388166 995424 388222 995480
rect 392398 995424 392454 995480
rect 393686 995424 393742 995480
rect 396538 995424 396594 995480
rect 423494 1006324 423550 1006360
rect 423494 1006304 423496 1006324
rect 423496 1006304 423548 1006324
rect 423548 1006304 423550 1006324
rect 421838 1006032 421894 1006088
rect 423494 1006052 423550 1006088
rect 423494 1006032 423496 1006052
rect 423496 1006032 423548 1006052
rect 423548 1006032 423550 1006052
rect 414478 996376 414534 996432
rect 416134 995696 416190 995752
rect 415398 995444 415454 995480
rect 415398 995424 415400 995444
rect 415400 995424 415452 995444
rect 415452 995424 415454 995444
rect 426346 1005660 426348 1005680
rect 426348 1005660 426400 1005680
rect 426400 1005660 426402 1005680
rect 426346 1005624 426402 1005660
rect 425518 1005524 425520 1005544
rect 425520 1005524 425572 1005544
rect 425572 1005524 425574 1005544
rect 425518 1005488 425574 1005524
rect 424322 1005388 424324 1005408
rect 424324 1005388 424376 1005408
rect 424376 1005388 424378 1005408
rect 424322 1005352 424378 1005388
rect 425150 1005252 425152 1005272
rect 425152 1005252 425204 1005272
rect 425204 1005252 425206 1005272
rect 425150 1005216 425206 1005252
rect 431682 1006052 431738 1006088
rect 431682 1006032 431684 1006052
rect 431684 1006032 431736 1006052
rect 431736 1006032 431738 1006052
rect 428002 1004980 428004 1005000
rect 428004 1004980 428056 1005000
rect 428056 1004980 428058 1005000
rect 428002 1004944 428058 1004980
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 426346 1004028 426348 1004048
rect 426348 1004028 426400 1004048
rect 426400 1004028 426402 1004048
rect 426346 1003992 426402 1004028
rect 427174 1002088 427230 1002144
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 424322 1001972 424378 1002008
rect 424322 1001952 424324 1001972
rect 424324 1001952 424376 1001972
rect 424376 1001952 424378 1001972
rect 427542 1001988 427544 1002008
rect 427544 1001988 427596 1002008
rect 427596 1001988 427598 1002008
rect 427542 1001952 427598 1001988
rect 432878 1004692 432934 1004728
rect 432878 1004672 432880 1004692
rect 432880 1004672 432932 1004692
rect 432932 1004672 432934 1004692
rect 428370 998844 428426 998880
rect 428370 998824 428372 998844
rect 428372 998824 428424 998844
rect 428424 998824 428426 998844
rect 430854 998572 430910 998608
rect 430854 998552 430856 998572
rect 430856 998552 430908 998572
rect 430908 998552 430910 998572
rect 430026 998300 430082 998336
rect 430026 998280 430028 998300
rect 430028 998280 430080 998300
rect 430080 998280 430082 998300
rect 431222 998164 431278 998200
rect 431222 998144 431224 998164
rect 431224 998144 431276 998164
rect 431276 998144 431278 998164
rect 432050 998028 432106 998064
rect 432050 998008 432052 998028
rect 432052 998008 432104 998028
rect 432104 998008 432106 998028
rect 430026 997772 430028 997792
rect 430028 997772 430080 997792
rect 430080 997772 430082 997792
rect 430026 997736 430082 997772
rect 435362 997736 435418 997792
rect 505006 1006732 505062 1006768
rect 505006 1006712 505008 1006732
rect 505008 1006712 505060 1006732
rect 505060 1006712 505062 1006732
rect 501326 1006596 501382 1006632
rect 501326 1006576 501328 1006596
rect 501328 1006576 501380 1006596
rect 501380 1006576 501382 1006596
rect 439686 997192 439742 997248
rect 439870 996920 439926 996976
rect 445022 996240 445078 996296
rect 462962 995560 463018 995616
rect 456798 995288 456854 995344
rect 505374 1006324 505430 1006360
rect 505374 1006304 505376 1006324
rect 505376 1006304 505428 1006324
rect 505428 1006304 505430 1006324
rect 507030 1006188 507086 1006224
rect 507030 1006168 507032 1006188
rect 507032 1006168 507084 1006188
rect 507084 1006168 507086 1006188
rect 466366 995968 466422 996024
rect 464342 994744 464398 994800
rect 447782 994472 447838 994528
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 502522 1006052 502578 1006088
rect 502522 1006032 502524 1006052
rect 502524 1006032 502576 1006052
rect 502576 1006032 502578 1006052
rect 506202 1006052 506258 1006088
rect 506202 1006032 506204 1006052
rect 506204 1006032 506256 1006052
rect 506256 1006032 506258 1006052
rect 509054 1006052 509110 1006088
rect 509054 1006032 509056 1006052
rect 509056 1006032 509108 1006052
rect 509108 1006032 509110 1006052
rect 471150 996240 471206 996296
rect 471426 995832 471482 995888
rect 469862 995016 469918 995072
rect 445666 994200 445722 994256
rect 488906 997192 488962 997248
rect 489090 996920 489146 996976
rect 478326 995696 478382 995752
rect 478970 995696 479026 995752
rect 485778 995696 485834 995752
rect 477682 995560 477738 995616
rect 489734 996648 489790 996704
rect 489918 996648 489974 996704
rect 472254 995016 472310 995072
rect 472438 995016 472494 995072
rect 474738 995016 474794 995072
rect 474922 995016 474978 995072
rect 476118 995016 476174 995072
rect 476302 995016 476358 995072
rect 480810 995288 480866 995344
rect 482926 994472 482982 994528
rect 485686 995424 485742 995480
rect 489274 995424 489330 995480
rect 486606 994744 486662 994800
rect 498842 1005252 498844 1005272
rect 498844 1005252 498896 1005272
rect 498896 1005252 498898 1005272
rect 498842 1005216 498898 1005252
rect 500498 1004964 500554 1005000
rect 500498 1004944 500500 1004964
rect 500500 1004944 500552 1004964
rect 500552 1004944 500554 1004964
rect 499670 1004828 499726 1004864
rect 499670 1004808 499672 1004828
rect 499672 1004808 499724 1004828
rect 499724 1004808 499726 1004828
rect 500498 1004692 500554 1004728
rect 500498 1004672 500500 1004692
rect 500500 1004672 500552 1004692
rect 500552 1004672 500554 1004692
rect 504546 1004420 504602 1004456
rect 504546 1004400 504548 1004420
rect 504548 1004400 504600 1004420
rect 504600 1004400 504602 1004420
rect 501694 1003332 501750 1003368
rect 501694 1003312 501696 1003332
rect 501696 1003312 501748 1003332
rect 501748 1003312 501750 1003332
rect 503350 1002380 503406 1002416
rect 503350 1002360 503352 1002380
rect 503352 1002360 503404 1002380
rect 503404 1002360 503406 1002380
rect 503350 1002108 503406 1002144
rect 503350 1002088 503352 1002108
rect 503352 1002088 503404 1002108
rect 503404 1002088 503406 1002108
rect 501694 1001972 501750 1002008
rect 501694 1001952 501696 1001972
rect 501696 1001952 501748 1001972
rect 501748 1001952 501750 1001972
rect 502522 1001952 502578 1002008
rect 504178 1001972 504234 1002008
rect 504178 1001952 504180 1001972
rect 504180 1001952 504232 1001972
rect 504232 1001952 504234 1001972
rect 505374 1001972 505430 1002008
rect 505374 1001952 505376 1001972
rect 505376 1001952 505428 1001972
rect 505428 1001952 505430 1001972
rect 508226 1005100 508282 1005136
rect 508226 1005080 508228 1005100
rect 508228 1005080 508280 1005100
rect 508280 1005080 508282 1005100
rect 508226 1004828 508282 1004864
rect 508226 1004808 508228 1004828
rect 508228 1004808 508280 1004828
rect 508280 1004808 508282 1004828
rect 507398 1004692 507454 1004728
rect 507398 1004672 507400 1004692
rect 507400 1004672 507452 1004692
rect 507452 1004672 507454 1004692
rect 509882 1002108 509938 1002144
rect 509882 1002088 509884 1002108
rect 509884 1002088 509936 1002108
rect 509936 1002088 509938 1002108
rect 510342 1001972 510398 1002008
rect 510342 1001952 510344 1001972
rect 510344 1001952 510396 1001972
rect 510396 1001952 510398 1001972
rect 510986 997192 511042 997248
rect 481914 994200 481970 994256
rect 516874 998552 516930 998608
rect 516690 996376 516746 996432
rect 517058 996920 517114 996976
rect 516874 995696 516930 995752
rect 517518 995288 517574 995344
rect 555974 1006732 556030 1006768
rect 555974 1006712 555976 1006732
rect 555976 1006712 556028 1006732
rect 556028 1006712 556030 1006732
rect 556802 1006596 556858 1006632
rect 556802 1006576 556804 1006596
rect 556804 1006576 556856 1006596
rect 556856 1006576 556858 1006596
rect 553122 1006460 553178 1006496
rect 553122 1006440 553124 1006460
rect 553124 1006440 553176 1006460
rect 553176 1006440 553178 1006460
rect 552294 1006324 552350 1006360
rect 552294 1006304 552296 1006324
rect 552296 1006304 552348 1006324
rect 552348 1006304 552350 1006324
rect 551466 1006188 551522 1006224
rect 551466 1006168 551468 1006188
rect 551468 1006168 551520 1006188
rect 551520 1006168 551522 1006188
rect 551098 1006032 551154 1006088
rect 555974 1006052 556030 1006088
rect 555974 1006032 555976 1006052
rect 555976 1006032 556028 1006052
rect 556028 1006032 556030 1006052
rect 520922 995968 520978 996024
rect 552294 1005388 552296 1005408
rect 552296 1005388 552348 1005408
rect 552348 1005388 552350 1005408
rect 552294 1005352 552350 1005388
rect 551466 1005252 551468 1005272
rect 551468 1005252 551520 1005272
rect 551520 1005252 551522 1005272
rect 551466 1005216 551522 1005252
rect 557170 1003892 557172 1003912
rect 557172 1003892 557224 1003912
rect 557224 1003892 557226 1003912
rect 557170 1003856 557226 1003892
rect 553950 1002380 554006 1002416
rect 553950 1002360 553952 1002380
rect 553952 1002360 554004 1002380
rect 554004 1002360 554006 1002380
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 523498 996648 523554 996704
rect 524050 997192 524106 997248
rect 555146 1002244 555202 1002280
rect 555146 1002224 555148 1002244
rect 555148 1002224 555200 1002244
rect 555200 1002224 555202 1002244
rect 554318 1001972 554374 1002008
rect 554318 1001952 554320 1001972
rect 554320 1001952 554372 1001972
rect 554372 1001952 554374 1001972
rect 555146 999132 555148 999152
rect 555148 999132 555200 999152
rect 555200 999132 555202 999152
rect 555146 999096 555202 999132
rect 553950 997772 553952 997792
rect 553952 997772 554004 997792
rect 554004 997772 554006 997792
rect 553950 997736 554006 997772
rect 540886 996920 540942 996976
rect 524050 996376 524106 996432
rect 549442 996396 549498 996432
rect 549442 996376 549444 996396
rect 549444 996376 549496 996396
rect 549496 996376 549498 996396
rect 529018 995696 529074 995752
rect 529662 995696 529718 995752
rect 532238 995696 532294 995752
rect 532790 995696 532846 995752
rect 534630 995696 534686 995752
rect 536562 995696 536618 995752
rect 527914 995016 527970 995072
rect 529846 995560 529902 995616
rect 535642 995288 535698 995344
rect 529662 995016 529718 995072
rect 538586 994508 538588 994528
rect 538588 994508 538640 994528
rect 538640 994508 538642 994528
rect 538586 994472 538642 994508
rect 557998 998300 558054 998336
rect 557998 998280 558000 998300
rect 558000 998280 558052 998300
rect 558052 998280 558054 998300
rect 557998 998028 558054 998064
rect 557998 998008 558000 998028
rect 558000 998008 558052 998028
rect 558052 998008 558054 998028
rect 557630 997892 557686 997928
rect 557630 997872 557632 997892
rect 557632 997872 557684 997892
rect 557684 997872 557686 997892
rect 560850 1004692 560906 1004728
rect 560850 1004672 560852 1004692
rect 560852 1004672 560904 1004692
rect 560904 1004672 560906 1004692
rect 560850 1002516 560906 1002552
rect 560850 1002496 560852 1002516
rect 560852 1002496 560904 1002516
rect 560904 1002496 560906 1002516
rect 560482 1002380 560538 1002416
rect 560482 1002360 560484 1002380
rect 560484 1002360 560536 1002380
rect 560536 1002360 560538 1002380
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 558826 998436 558882 998472
rect 558826 998416 558828 998436
rect 558828 998416 558880 998436
rect 558880 998416 558882 998436
rect 558826 998164 558882 998200
rect 558826 998144 558828 998164
rect 558828 998144 558880 998164
rect 558880 998144 558882 998164
rect 560022 997892 560078 997928
rect 560022 997872 560024 997892
rect 560024 997872 560076 997892
rect 560076 997872 560078 997892
rect 570418 994744 570474 994800
rect 590566 996920 590622 996976
rect 623686 997192 623742 997248
rect 590566 996648 590622 996704
rect 590566 996412 590568 996432
rect 590568 996412 590620 996432
rect 590620 996412 590622 996432
rect 590566 996376 590622 996412
rect 590750 995288 590806 995344
rect 590566 995016 590622 995072
rect 625434 995968 625490 996024
rect 625618 995696 625674 995752
rect 627182 995696 627238 995752
rect 627918 995696 627974 995752
rect 629574 995696 629630 995752
rect 630310 995696 630366 995752
rect 633990 995696 634046 995752
rect 635278 995696 635334 995752
rect 637026 995696 637082 995752
rect 630862 994744 630918 994800
rect 634726 995288 634782 995344
rect 640982 995016 641038 995072
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 937216 660358 937272
rect 664442 947280 664498 947336
rect 663062 941704 663118 941760
rect 665822 939800 665878 939856
rect 674378 966048 674434 966104
rect 673366 962784 673422 962840
rect 673182 962512 673238 962568
rect 672998 958704 673054 958760
rect 668582 938440 668638 938496
rect 672170 938032 672226 938088
rect 667202 937760 667258 937816
rect 672814 937760 672870 937816
rect 672630 937488 672686 937544
rect 672170 937216 672226 937272
rect 671802 936672 671858 936728
rect 658922 935992 658978 936048
rect 671618 935720 671674 935776
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 55862 892744 55918 892800
rect 54482 892472 54538 892528
rect 53286 892200 53342 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62762 858608 62818 858664
rect 62118 845552 62174 845608
rect 53102 799040 53158 799096
rect 62118 832496 62174 832552
rect 54482 774288 54538 774344
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 652390 856296 652446 856352
rect 652022 842968 652078 843024
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 62946 793600 63002 793656
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 55862 772792 55918 772848
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 50342 730496 50398 730552
rect 48962 669296 49018 669352
rect 47398 638152 47454 638208
rect 47398 618840 47454 618896
rect 45374 598032 45430 598088
rect 62762 743008 62818 743064
rect 651470 789928 651526 789984
rect 651470 776600 651526 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62946 741648 63002 741704
rect 62118 741240 62174 741296
rect 51722 691328 51778 691384
rect 51722 646584 51778 646640
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 50342 626592 50398 626648
rect 51722 601704 51778 601760
rect 48962 601296 49018 601352
rect 651470 723424 651526 723480
rect 652574 736752 652630 736808
rect 652022 718256 652078 718312
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652574 710232 652630 710288
rect 62762 697856 62818 697912
rect 652390 696940 652392 696960
rect 652392 696940 652444 696960
rect 652444 696940 652446 696960
rect 652390 696904 652446 696940
rect 62118 689152 62174 689208
rect 652022 683576 652078 683632
rect 62118 676096 62174 676152
rect 651470 670384 651526 670440
rect 62118 663040 62174 663096
rect 651470 657056 651526 657112
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 651470 630536 651526 630592
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 54482 600888 54538 600944
rect 47582 582392 47638 582448
rect 48962 557776 49018 557832
rect 51722 557504 51778 557560
rect 45558 556824 45614 556880
rect 45098 555600 45154 555656
rect 44822 555192 44878 555248
rect 44638 428848 44694 428904
rect 45006 551520 45062 551576
rect 45374 550840 45430 550896
rect 45190 548664 45246 548720
rect 45190 536968 45246 537024
rect 45374 532752 45430 532808
rect 45006 529624 45062 529680
rect 45558 429664 45614 429720
rect 45006 429256 45062 429312
rect 44822 428032 44878 428088
rect 44362 427216 44418 427272
rect 44454 426808 44510 426864
rect 44178 385600 44234 385656
rect 44638 421504 44694 421560
rect 44822 420688 44878 420744
rect 44638 406952 44694 407008
rect 44638 385192 44694 385248
rect 44454 383968 44510 384024
rect 45190 427624 45246 427680
rect 45006 386688 45062 386744
rect 45374 422320 45430 422376
rect 45374 405592 45430 405648
rect 45374 386008 45430 386064
rect 45190 384784 45246 384840
rect 45006 384376 45062 384432
rect 44454 377848 44510 377904
rect 44270 377440 44326 377496
rect 44454 364928 44510 364984
rect 44270 356632 44326 356688
rect 45190 383560 45246 383616
rect 43902 354184 43958 354240
rect 44730 353776 44786 353832
rect 28538 351192 28594 351248
rect 38290 346296 38346 346352
rect 28906 344256 28962 344312
rect 28538 343848 28594 343904
rect 45006 341672 45062 341728
rect 45558 383152 45614 383208
rect 45742 379072 45798 379128
rect 47582 430072 47638 430128
rect 46938 426400 46994 426456
rect 47122 423544 47178 423600
rect 47122 400152 47178 400208
rect 46938 399744 46994 399800
rect 46938 380704 46994 380760
rect 46202 366968 46258 367024
rect 45742 364248 45798 364304
rect 45558 356904 45614 356960
rect 45650 356632 45706 356688
rect 45926 355816 45982 355872
rect 45374 343304 45430 343360
rect 45190 340856 45246 340912
rect 35806 339768 35862 339824
rect 35806 338952 35862 339008
rect 31022 338544 31078 338600
rect 31022 329024 31078 329080
rect 45650 338408 45706 338464
rect 45466 337184 45522 337240
rect 37922 335280 37978 335336
rect 42798 334600 42854 334656
rect 43166 334600 43222 334656
rect 44270 334600 44326 334656
rect 36542 328344 36598 328400
rect 41786 326712 41842 326768
rect 41786 325352 41842 325408
rect 41786 324672 41842 324728
rect 42246 323584 42302 323640
rect 42062 322768 42118 322824
rect 42430 321408 42486 321464
rect 41786 321136 41842 321192
rect 42430 320048 42486 320104
rect 42430 318824 42486 318880
rect 42982 334328 43038 334384
rect 42982 323584 43038 323640
rect 43442 322904 43498 322960
rect 43166 322768 43222 322824
rect 42430 316376 42486 316432
rect 42154 315968 42210 316024
rect 41878 315560 41934 315616
rect 42154 313656 42210 313712
rect 42430 312704 42486 312760
rect 42062 312568 42118 312624
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 42890 299648 42946 299704
rect 41786 296792 41842 296848
rect 41326 295976 41382 296032
rect 32402 294752 32458 294808
rect 41786 292440 41842 292496
rect 41786 290400 41842 290456
rect 41326 290264 41382 290320
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42430 278704 42486 278760
rect 42338 278432 42394 278488
rect 41786 277888 41842 277944
rect 42154 277888 42210 277944
rect 42062 277072 42118 277128
rect 42062 276528 42118 276584
rect 41786 274216 41842 274272
rect 42062 273400 42118 273456
rect 42062 272992 42118 273048
rect 41786 270408 41842 270464
rect 42430 270408 42486 270464
rect 41786 269048 41842 269104
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 43258 298832 43314 298888
rect 43074 295160 43130 295216
rect 43074 276528 43130 276584
rect 42890 256808 42946 256864
rect 44270 320048 44326 320104
rect 45650 318824 45706 318880
rect 45466 315968 45522 316024
rect 44730 311480 44786 311536
rect 44362 311208 44418 311264
rect 44546 311072 44602 311128
rect 47122 379888 47178 379944
rect 47122 357312 47178 357368
rect 46938 356088 46994 356144
rect 46938 340040 46994 340096
rect 47582 333104 47638 333160
rect 46938 313656 46994 313712
rect 46386 303048 46442 303104
rect 44730 300056 44786 300112
rect 44546 299240 44602 299296
rect 44362 298424 44418 298480
rect 44178 298016 44234 298072
rect 43626 293936 43682 293992
rect 43810 293120 43866 293176
rect 43994 291896 44050 291952
rect 43810 279792 43866 279848
rect 43994 277072 44050 277128
rect 43626 272992 43682 273048
rect 43442 257624 43498 257680
rect 43626 256400 43682 256456
rect 43258 255992 43314 256048
rect 42982 255584 43038 255640
rect 42798 254768 42854 254824
rect 35438 253408 35494 253464
rect 35622 253000 35678 253056
rect 35806 252592 35862 252648
rect 35806 252184 35862 252240
rect 41326 252184 41382 252240
rect 42614 252184 42670 252240
rect 41694 242836 41696 242856
rect 41696 242836 41748 242856
rect 41748 242836 41750 242856
rect 41694 242800 41750 242836
rect 42338 242800 42394 242856
rect 40682 242528 40738 242584
rect 41786 240080 41842 240136
rect 42062 238448 42118 238504
rect 41786 235864 41842 235920
rect 42154 235320 42210 235376
rect 42522 238040 42578 238096
rect 42246 234096 42302 234152
rect 42430 233824 42486 233880
rect 42338 233144 42394 233200
rect 42430 231784 42486 231840
rect 42154 230152 42210 230208
rect 42430 229336 42486 229392
rect 41970 227296 42026 227352
rect 42154 226616 42210 226672
rect 42430 225664 42486 225720
rect 40682 222808 40738 222864
rect 35530 217912 35586 217968
rect 35530 214240 35586 214296
rect 35806 214240 35862 214296
rect 43442 251096 43498 251152
rect 43258 242528 43314 242584
rect 44638 297200 44694 297256
rect 44362 294344 44418 294400
rect 44362 270408 44418 270464
rect 44178 255176 44234 255232
rect 44638 254360 44694 254416
rect 44178 253952 44234 254008
rect 43350 226616 43406 226672
rect 43166 225664 43222 225720
rect 43718 249056 43774 249112
rect 43718 231784 43774 231840
rect 43534 213696 43590 213752
rect 42982 212880 43038 212936
rect 42798 212064 42854 212120
rect 35806 211384 35862 211440
rect 44546 251912 44602 251968
rect 44362 248648 44418 248704
rect 44362 234096 44418 234152
rect 44546 233144 44602 233200
rect 45006 293528 45062 293584
rect 45190 291624 45246 291680
rect 46202 290672 46258 290728
rect 45190 277888 45246 277944
rect 45006 273400 45062 273456
rect 45558 250688 45614 250744
rect 45006 248240 45062 248296
rect 45006 235320 45062 235376
rect 45834 250280 45890 250336
rect 46018 249464 46074 249520
rect 46018 233824 46074 233880
rect 45834 230152 45890 230208
rect 45558 229336 45614 229392
rect 44822 214920 44878 214976
rect 45006 213288 45062 213344
rect 44178 211248 44234 211304
rect 43258 210840 43314 210896
rect 42798 209344 42854 209400
rect 35806 208936 35862 208992
rect 41694 208936 41750 208992
rect 40038 207712 40094 207768
rect 35622 204040 35678 204096
rect 35806 203632 35862 203688
rect 35622 202136 35678 202192
rect 37922 197784 37978 197840
rect 41786 197104 41842 197160
rect 41878 195744 41934 195800
rect 42614 195472 42670 195528
rect 41786 195200 41842 195256
rect 42430 193160 42486 193216
rect 42614 192888 42670 192944
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41786 187176 41842 187232
rect 42338 186088 42394 186144
rect 41970 185816 42026 185872
rect 42430 184864 42486 184920
rect 42430 183096 42486 183152
rect 42982 206352 43038 206408
rect 44178 210432 44234 210488
rect 43442 207984 43498 208040
rect 43258 206216 43314 206272
rect 43994 206760 44050 206816
rect 42982 191120 43038 191176
rect 43810 205536 43866 205592
rect 43626 205128 43682 205184
rect 43442 202136 43498 202192
rect 43258 183096 43314 183152
rect 43626 191664 43682 191720
rect 43994 193160 44050 193216
rect 43810 190440 43866 190496
rect 44362 208528 44418 208584
rect 44546 205944 44602 206000
rect 44362 189896 44418 189952
rect 44822 204720 44878 204776
rect 44546 187584 44602 187640
rect 44178 184864 44234 184920
rect 46938 247016 46994 247072
rect 46938 238448 46994 238504
rect 50342 430888 50398 430944
rect 48962 386960 49018 387016
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 49146 346296 49202 346352
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 212472 48006 212528
rect 47950 192344 48006 192400
rect 48778 190440 48834 190496
rect 49146 289856 49202 289912
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 62118 597896 62174 597952
rect 651470 590708 651526 590744
rect 651470 590688 651472 590708
rect 651472 590688 651524 590708
rect 651524 590688 651526 590708
rect 62118 584840 62174 584896
rect 669226 879144 669282 879200
rect 664442 868672 664498 868728
rect 668214 868128 668270 868184
rect 663062 760824 663118 760880
rect 661682 760416 661738 760472
rect 660302 625232 660358 625288
rect 660302 599528 660358 599584
rect 652022 582936 652078 582992
rect 666282 777008 666338 777064
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661866 643728 661922 643784
rect 661682 581032 661738 581088
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 658922 553968 658978 554024
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 652574 497664 652630 497720
rect 62118 493584 62174 493640
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 55862 408448 55918 408504
rect 651470 404640 651526 404696
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51722 301280 51778 301336
rect 51722 289856 51778 289912
rect 50342 257760 50398 257816
rect 50526 247696 50582 247752
rect 50342 246472 50398 246528
rect 49330 208936 49386 208992
rect 49514 206216 49570 206272
rect 49330 196424 49386 196480
rect 49514 194384 49570 194440
rect 50710 203224 50766 203280
rect 652574 391448 652630 391504
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 652022 378120 652078 378176
rect 62118 376216 62174 376272
rect 651654 364792 651710 364848
rect 62118 363296 62174 363352
rect 651470 351600 651526 351656
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 55862 278704 55918 278760
rect 651470 338272 651526 338328
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 651470 285232 651526 285288
rect 62946 285096 63002 285152
rect 62762 267008 62818 267064
rect 54482 217912 54538 217968
rect 136546 269728 136602 269784
rect 139950 269764 139952 269784
rect 139952 269764 140004 269784
rect 140004 269764 140006 269784
rect 139950 269728 140006 269764
rect 485732 267436 485788 267472
rect 485732 267416 485734 267436
rect 485734 267416 485786 267436
rect 485786 267416 485788 267436
rect 485686 266872 485742 266928
rect 486054 266872 486110 266928
rect 487250 267436 487306 267472
rect 487250 267416 487252 267436
rect 487252 267416 487304 267436
rect 487304 267416 487306 267436
rect 492310 267824 492366 267880
rect 494150 270000 494206 270056
rect 498198 267824 498254 267880
rect 499578 267164 499634 267200
rect 499578 267144 499580 267164
rect 499580 267144 499632 267164
rect 499632 267144 499634 267164
rect 501050 267144 501106 267200
rect 504178 270544 504234 270600
rect 503074 269592 503130 269648
rect 504546 269628 504548 269648
rect 504548 269628 504600 269648
rect 504600 269628 504602 269648
rect 504546 269592 504602 269628
rect 507858 270544 507914 270600
rect 511722 271396 511724 271416
rect 511724 271396 511776 271416
rect 511776 271396 511778 271416
rect 511722 271360 511778 271396
rect 509882 269728 509938 269784
rect 513194 272312 513250 272368
rect 515310 271396 515312 271416
rect 515312 271396 515364 271416
rect 515364 271396 515366 271416
rect 515310 271360 515366 271396
rect 516598 274100 516654 274136
rect 516598 274080 516600 274100
rect 516600 274080 516652 274100
rect 516652 274080 516654 274100
rect 517058 274080 517114 274136
rect 518438 272312 518494 272368
rect 518438 268504 518494 268560
rect 518990 268504 519046 268560
rect 516966 267688 517022 267744
rect 519174 268368 519230 268424
rect 518990 267708 519046 267744
rect 518990 267688 518992 267708
rect 518992 267688 519044 267708
rect 519044 267688 519046 267708
rect 519174 267144 519230 267200
rect 521106 273672 521162 273728
rect 520462 268388 520518 268424
rect 520462 268368 520464 268388
rect 520464 268368 520516 268388
rect 520516 268368 520518 268388
rect 521474 272584 521530 272640
rect 522026 270852 522028 270872
rect 522028 270852 522080 270872
rect 522080 270852 522082 270872
rect 522026 270816 522082 270852
rect 524234 273672 524290 273728
rect 523958 271632 524014 271688
rect 523314 269728 523370 269784
rect 521658 269456 521714 269512
rect 524878 272620 524880 272640
rect 524880 272620 524932 272640
rect 524932 272620 524934 272640
rect 524878 272584 524934 272620
rect 524510 272312 524566 272368
rect 525798 275712 525854 275768
rect 524694 271632 524750 271688
rect 524786 270852 524788 270872
rect 524788 270852 524840 270872
rect 524840 270852 524842 270872
rect 524786 270816 524842 270852
rect 526258 270952 526314 271008
rect 525522 268640 525578 268696
rect 527362 275732 527418 275768
rect 527362 275712 527364 275732
rect 527364 275712 527416 275732
rect 527416 275712 527418 275732
rect 528006 273808 528062 273864
rect 527178 267144 527234 267200
rect 528650 270716 528652 270736
rect 528652 270716 528704 270736
rect 528704 270716 528706 270736
rect 528650 270680 528706 270716
rect 529202 271224 529258 271280
rect 529570 270952 529626 271008
rect 531594 272312 531650 272368
rect 531410 270000 531466 270056
rect 530950 269456 531006 269512
rect 530950 269048 531006 269104
rect 533894 274216 533950 274272
rect 533894 273808 533950 273864
rect 534906 275712 534962 275768
rect 535090 275032 535146 275088
rect 534078 272720 534134 272776
rect 533710 272448 533766 272504
rect 534170 272484 534172 272504
rect 534172 272484 534224 272504
rect 534224 272484 534226 272504
rect 534170 272448 534226 272484
rect 533158 270680 533214 270736
rect 533526 269728 533582 269784
rect 532238 267008 532294 267064
rect 534354 269728 534410 269784
rect 533894 269048 533950 269104
rect 533894 268640 533950 268696
rect 533894 267980 533950 268016
rect 533894 267960 533896 267980
rect 533896 267960 533948 267980
rect 533948 267960 533950 267980
rect 533986 267708 534042 267744
rect 533986 267688 533988 267708
rect 533988 267688 534040 267708
rect 534040 267688 534042 267708
rect 533894 267300 533950 267336
rect 533894 267280 533896 267300
rect 533896 267280 533948 267300
rect 533948 267280 533950 267300
rect 534170 267280 534226 267336
rect 538034 275712 538090 275768
rect 538218 275460 538274 275496
rect 538218 275440 538220 275460
rect 538220 275440 538272 275460
rect 538272 275440 538274 275460
rect 536746 273808 536802 273864
rect 535918 269456 535974 269512
rect 535458 267960 535514 268016
rect 538402 275032 538458 275088
rect 538678 275032 538734 275088
rect 538218 274760 538274 274816
rect 539046 275440 539102 275496
rect 539046 274216 539102 274272
rect 537022 269220 537024 269240
rect 537024 269220 537076 269240
rect 537076 269220 537078 269240
rect 537022 269184 537078 269220
rect 538310 270544 538366 270600
rect 538034 269728 538090 269784
rect 541162 275032 541218 275088
rect 538678 269184 538734 269240
rect 539230 268096 539286 268152
rect 538310 267688 538366 267744
rect 538678 266620 538734 266656
rect 538678 266600 538680 266620
rect 538680 266600 538732 266620
rect 538732 266600 538734 266620
rect 543186 274760 543242 274816
rect 544474 272720 544530 272776
rect 543002 272448 543058 272504
rect 541990 269456 542046 269512
rect 542174 267280 542230 267336
rect 543554 271496 543610 271552
rect 546222 271496 546278 271552
rect 543554 270544 543610 270600
rect 543554 267708 543610 267744
rect 547510 268388 547566 268424
rect 547510 268368 547512 268388
rect 547512 268368 547564 268388
rect 547564 268368 547566 268388
rect 547694 268096 547750 268152
rect 543554 267688 543556 267708
rect 543556 267688 543608 267708
rect 543608 267688 543610 267708
rect 546590 267708 546646 267744
rect 546590 267688 546592 267708
rect 546592 267688 546644 267708
rect 546644 267688 546646 267708
rect 543554 266600 543610 266656
rect 552202 270680 552258 270736
rect 549258 268368 549314 268424
rect 553398 270680 553454 270736
rect 574926 270272 574982 270328
rect 607862 267280 607918 267336
rect 625066 271088 625122 271144
rect 627918 270000 627974 270056
rect 635646 273808 635702 273864
rect 637578 269728 637634 269784
rect 645122 272448 645178 272504
rect 629298 267008 629354 267064
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553674 255584 553730 255640
rect 553490 251252 553546 251288
rect 553490 251232 553492 251252
rect 553492 251232 553544 251252
rect 553544 251232 553546 251252
rect 554502 253428 554558 253464
rect 554502 253408 554504 253428
rect 554504 253408 554556 253428
rect 554556 253408 554558 253428
rect 553858 249056 553914 249112
rect 554410 246880 554466 246936
rect 554502 244704 554558 244760
rect 553950 242528 554006 242584
rect 553858 240352 553914 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 62946 222808 63002 222864
rect 73066 226888 73122 226944
rect 68926 224168 68982 224224
rect 69754 220088 69810 220144
rect 72882 220360 72938 220416
rect 79966 228248 80022 228304
rect 103610 229744 103666 229800
rect 101862 221448 101918 221504
rect 123390 222808 123446 222864
rect 133786 227840 133842 227896
rect 139306 226480 139362 226536
rect 136546 225256 136602 225312
rect 138294 221720 138350 221776
rect 137834 219136 137890 219192
rect 138110 219156 138166 219192
rect 138110 219136 138112 219156
rect 138112 219136 138164 219156
rect 138164 219136 138166 219156
rect 141330 227860 141386 227896
rect 141330 227840 141332 227860
rect 141332 227840 141384 227860
rect 141384 227840 141386 227860
rect 142158 227160 142214 227216
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 142250 225292 142252 225312
rect 142252 225292 142304 225312
rect 142304 225292 142306 225312
rect 142250 225256 142306 225292
rect 143078 227160 143134 227216
rect 143170 225528 143226 225584
rect 140962 223932 140964 223952
rect 140964 223932 141016 223952
rect 141016 223932 141018 223952
rect 140962 223896 141018 223932
rect 140778 220108 140834 220144
rect 140778 220088 140780 220108
rect 140780 220088 140832 220108
rect 140832 220088 140834 220108
rect 142434 221176 142490 221232
rect 142250 219020 142306 219056
rect 142250 219000 142252 219020
rect 142252 219000 142304 219020
rect 142304 219000 142306 219020
rect 145654 229744 145710 229800
rect 146298 229356 146354 229392
rect 146298 229336 146300 229356
rect 146300 229336 146352 229356
rect 146352 229336 146354 229356
rect 145930 225256 145986 225312
rect 145654 224032 145710 224088
rect 145378 223896 145434 223952
rect 144182 221196 144238 221232
rect 144182 221176 144184 221196
rect 144184 221176 144236 221196
rect 144236 221176 144238 221196
rect 145654 219000 145710 219056
rect 147034 225936 147090 225992
rect 147954 229336 148010 229392
rect 147678 228520 147734 228576
rect 147402 225564 147404 225584
rect 147404 225564 147456 225584
rect 147456 225564 147458 225584
rect 147402 225528 147458 225564
rect 147770 224032 147826 224088
rect 147310 222128 147366 222184
rect 146574 221720 146630 221776
rect 147494 221856 147550 221912
rect 147494 220244 147550 220280
rect 147494 220224 147496 220244
rect 147496 220224 147548 220244
rect 147548 220224 147550 220244
rect 146390 220088 146446 220144
rect 147034 219408 147090 219464
rect 147494 218748 147550 218784
rect 147494 218728 147496 218748
rect 147496 218728 147548 218748
rect 147548 218728 147550 218748
rect 148230 220224 148286 220280
rect 148046 219408 148102 219464
rect 149794 228520 149850 228576
rect 150162 227180 150218 227216
rect 150162 227160 150164 227180
rect 150164 227160 150216 227180
rect 150216 227160 150218 227180
rect 149058 221856 149114 221912
rect 150070 220768 150126 220824
rect 148598 218728 148654 218784
rect 151910 227432 151966 227488
rect 151726 223760 151782 223816
rect 151082 219816 151138 219872
rect 152922 227432 152978 227488
rect 153106 226072 153162 226128
rect 152830 225936 152886 225992
rect 152462 224304 152518 224360
rect 152094 222128 152150 222184
rect 153290 225256 153346 225312
rect 153658 220496 153714 220552
rect 152094 218884 152150 218920
rect 152094 218864 152096 218884
rect 152096 218864 152148 218884
rect 152148 218864 152150 218884
rect 154578 227160 154634 227216
rect 155866 227976 155922 228032
rect 155314 226888 155370 226944
rect 155038 223080 155094 223136
rect 153842 218864 153898 218920
rect 156142 220768 156198 220824
rect 157430 228520 157486 228576
rect 157982 229336 158038 229392
rect 157798 227976 157854 228032
rect 157614 226108 157616 226128
rect 157616 226108 157668 226128
rect 157668 226108 157670 226128
rect 157614 226072 157670 226108
rect 156694 224032 156750 224088
rect 157062 224304 157118 224360
rect 157430 224032 157486 224088
rect 157246 223760 157302 223816
rect 157246 223388 157248 223408
rect 157248 223388 157300 223408
rect 157300 223388 157302 223408
rect 157246 223352 157302 223388
rect 157430 223388 157432 223408
rect 157432 223388 157484 223408
rect 157484 223388 157486 223408
rect 157430 223352 157486 223388
rect 157062 223116 157064 223136
rect 157064 223116 157116 223136
rect 157116 223116 157118 223136
rect 157062 223080 157118 223116
rect 157338 220380 157394 220416
rect 157338 220360 157340 220380
rect 157340 220360 157392 220380
rect 157392 220360 157394 220380
rect 157246 218592 157302 218648
rect 157706 218592 157762 218648
rect 158810 228520 158866 228576
rect 159638 227452 159694 227488
rect 159638 227432 159640 227452
rect 159640 227432 159692 227452
rect 159692 227432 159694 227452
rect 160466 228248 160522 228304
rect 158350 223080 158406 223136
rect 160834 222536 160890 222592
rect 161570 225528 161626 225584
rect 162306 222536 162362 222592
rect 161478 220360 161534 220416
rect 163870 229356 163926 229392
rect 163870 229336 163872 229356
rect 163872 229336 163924 229356
rect 163924 229336 163926 229356
rect 162950 224304 163006 224360
rect 163962 223896 164018 223952
rect 166630 228384 166686 228440
rect 166446 227432 166502 227488
rect 166814 225836 166816 225856
rect 166816 225836 166868 225856
rect 166868 225836 166870 225856
rect 166814 225800 166870 225836
rect 166722 225528 166778 225584
rect 166538 225020 166540 225040
rect 166540 225020 166592 225040
rect 166592 225020 166594 225040
rect 166538 224984 166594 225020
rect 165802 223116 165804 223136
rect 165804 223116 165856 223136
rect 165856 223116 165858 223136
rect 165802 223080 165858 223116
rect 165618 222808 165674 222864
rect 166814 223252 166816 223272
rect 166816 223252 166868 223272
rect 166868 223252 166870 223272
rect 166814 223216 166870 223252
rect 166262 219136 166318 219192
rect 166446 218884 166502 218920
rect 166446 218864 166448 218884
rect 166448 218864 166500 218884
rect 166500 218864 166502 218884
rect 166538 218612 166594 218648
rect 166538 218592 166540 218612
rect 166540 218592 166592 218612
rect 166592 218592 166594 218612
rect 167182 219136 167238 219192
rect 166998 218864 167054 218920
rect 167182 218592 167238 218648
rect 166262 218320 166318 218376
rect 167366 218320 167422 218376
rect 169850 225800 169906 225856
rect 171138 228656 171194 228712
rect 171230 228384 171286 228440
rect 170862 225936 170918 225992
rect 171230 225972 171232 225992
rect 171232 225972 171284 225992
rect 171284 225972 171286 225992
rect 171230 225936 171286 225972
rect 171046 225700 171048 225720
rect 171048 225700 171100 225720
rect 171100 225700 171102 225720
rect 171046 225664 171102 225700
rect 171046 225020 171048 225040
rect 171048 225020 171100 225040
rect 171100 225020 171102 225040
rect 171046 224984 171102 225020
rect 170954 224204 170956 224224
rect 170956 224204 171008 224224
rect 171008 224204 171010 224224
rect 170954 224168 171010 224204
rect 172426 228792 172482 228848
rect 172242 228676 172298 228712
rect 172242 228656 172244 228676
rect 172244 228656 172296 228676
rect 172296 228656 172298 228676
rect 171414 224168 171470 224224
rect 170954 223896 171010 223952
rect 170402 223216 170458 223272
rect 171230 222264 171286 222320
rect 171046 221856 171102 221912
rect 171506 221876 171562 221912
rect 171506 221856 171508 221876
rect 171508 221856 171560 221876
rect 171560 221856 171562 221876
rect 174174 228812 174230 228848
rect 174174 228792 174176 228812
rect 174176 228792 174228 228812
rect 174228 228792 174230 228812
rect 174818 228792 174874 228848
rect 175738 228812 175794 228848
rect 175738 228792 175740 228812
rect 175740 228792 175792 228812
rect 175792 228792 175794 228812
rect 176658 226072 176714 226128
rect 176934 225664 176990 225720
rect 176474 225256 176530 225312
rect 176750 225256 176806 225312
rect 176106 222028 176108 222048
rect 176108 222028 176160 222048
rect 176160 222028 176162 222048
rect 176106 221992 176162 222028
rect 176658 222264 176714 222320
rect 176842 221992 176898 222048
rect 177394 221720 177450 221776
rect 178038 221448 178094 221504
rect 180798 226072 180854 226128
rect 181074 226072 181130 226128
rect 181258 221448 181314 221504
rect 184846 225664 184902 225720
rect 186042 226072 186098 226128
rect 186272 226024 186328 226026
rect 186272 225972 186274 226024
rect 186274 225972 186326 226024
rect 186326 225972 186328 226024
rect 186272 225970 186328 225972
rect 185674 225428 185676 225448
rect 185676 225428 185728 225448
rect 185728 225428 185730 225448
rect 185674 225392 185730 225428
rect 186410 225664 186466 225720
rect 186594 225392 186650 225448
rect 186870 225392 186926 225448
rect 186318 225120 186374 225176
rect 187238 225936 187294 225992
rect 185030 221720 185086 221776
rect 185858 221448 185914 221504
rect 188342 228812 188398 228848
rect 188342 228792 188344 228812
rect 188344 228792 188396 228812
rect 188396 228792 188398 228812
rect 190366 228792 190422 228848
rect 194874 225392 194930 225448
rect 195518 225120 195574 225176
rect 195058 219272 195114 219328
rect 196070 219292 196126 219328
rect 196070 219272 196072 219292
rect 196072 219272 196124 219292
rect 196124 219272 196126 219292
rect 202694 225120 202750 225176
rect 205086 225156 205088 225176
rect 205088 225156 205140 225176
rect 205140 225156 205142 225176
rect 205086 225120 205142 225156
rect 484582 219408 484638 219464
rect 486606 220904 486662 220960
rect 487802 218048 487858 218104
rect 490562 219136 490618 219192
rect 491114 219136 491170 219192
rect 490286 218864 490342 218920
rect 491114 218592 491170 218648
rect 492126 217096 492182 217152
rect 492954 219136 493010 219192
rect 493598 219136 493654 219192
rect 494794 219680 494850 219736
rect 493598 217232 493654 217288
rect 497738 219136 497794 219192
rect 496910 218320 496966 218376
rect 497554 217232 497610 217288
rect 498658 217776 498714 217832
rect 500038 218340 500094 218376
rect 500038 218320 500040 218340
rect 500040 218320 500092 218340
rect 500092 218320 500094 218340
rect 500222 218320 500278 218376
rect 502522 219136 502578 219192
rect 502706 219136 502762 219192
rect 503534 217504 503590 217560
rect 505098 219136 505154 219192
rect 505282 219136 505338 219192
rect 504822 218592 504878 218648
rect 505006 218628 505008 218648
rect 505008 218628 505060 218648
rect 505060 218628 505062 218648
rect 505006 218592 505062 218628
rect 504638 218320 504694 218376
rect 505282 218320 505338 218376
rect 504822 217776 504878 217832
rect 505834 217776 505890 217832
rect 506018 217776 506074 217832
rect 508502 217776 508558 217832
rect 510158 218592 510214 218648
rect 510986 219952 511042 220008
rect 509698 218320 509754 218376
rect 513378 221604 513434 221640
rect 513378 221584 513380 221604
rect 513380 221584 513432 221604
rect 513432 221584 513434 221604
rect 512642 219952 512698 220008
rect 515770 221176 515826 221232
rect 514758 219136 514814 219192
rect 514942 219156 514998 219192
rect 514942 219136 514944 219156
rect 514944 219136 514996 219156
rect 514996 219136 514998 219156
rect 517702 221720 517758 221776
rect 519542 220224 519598 220280
rect 519542 219680 519598 219736
rect 519818 219680 519874 219736
rect 522578 219716 522580 219736
rect 522580 219716 522632 219736
rect 522632 219716 522634 219736
rect 522578 219680 522634 219716
rect 526442 219952 526498 220008
rect 530030 219952 530086 220008
rect 533710 220496 533766 220552
rect 533710 219952 533766 220008
rect 533618 217776 533674 217832
rect 534446 217504 534502 217560
rect 541898 220496 541954 220552
rect 544658 220496 544714 220552
rect 544198 220224 544254 220280
rect 547418 220496 547474 220552
rect 547602 219136 547658 219192
rect 548154 219136 548210 219192
rect 548154 218592 548210 218648
rect 549074 220496 549130 220552
rect 549258 218320 549314 218376
rect 553490 220516 553546 220552
rect 553490 220496 553492 220516
rect 553492 220496 553544 220516
rect 553544 220496 553546 220516
rect 553674 218320 553730 218376
rect 554042 218320 554098 218376
rect 555422 221992 555478 222048
rect 554962 220496 555018 220552
rect 555238 220224 555294 220280
rect 555606 220632 555662 220688
rect 558550 220652 558606 220688
rect 558550 220632 558552 220652
rect 558552 220632 558604 220652
rect 558604 220632 558606 220652
rect 558550 219680 558606 219736
rect 559746 220496 559802 220552
rect 559102 219680 559158 219736
rect 559378 219680 559434 219736
rect 562230 222264 562286 222320
rect 562046 220496 562102 220552
rect 562598 221992 562654 222048
rect 563150 221992 563206 222048
rect 563426 220496 563482 220552
rect 562874 219680 562930 219736
rect 562874 218048 562930 218104
rect 563242 217640 563298 217696
rect 565726 222536 565782 222592
rect 567382 222536 567438 222592
rect 565680 217368 565736 217424
rect 566002 217402 566058 217458
rect 568026 219680 568082 219736
rect 571246 218150 571302 218206
rect 571890 222264 571946 222320
rect 572626 222536 572682 222592
rect 572166 222152 572222 222208
rect 572350 220496 572406 220552
rect 572166 219680 572222 219736
rect 572994 220088 573050 220144
rect 575938 222128 575994 222184
rect 572626 218592 572682 218648
rect 572810 218456 572866 218512
rect 574742 218286 574798 218342
rect 572166 217912 572222 217968
rect 572442 217504 572498 217560
rect 574466 218048 574522 218104
rect 574282 217504 574338 217560
rect 574926 217504 574982 217560
rect 575478 215056 575534 215112
rect 577594 220632 577650 220688
rect 576858 215056 576914 215112
rect 576306 214920 576362 214976
rect 582102 220088 582158 220144
rect 582102 219136 582158 219192
rect 582286 219172 582288 219192
rect 582288 219172 582340 219192
rect 582340 219172 582342 219192
rect 582286 219136 582342 219172
rect 586150 219136 586206 219192
rect 586334 219136 586390 219192
rect 582332 218592 582388 218648
rect 582194 218456 582250 218512
rect 586518 218320 586574 218376
rect 586334 218204 586390 218240
rect 586334 218184 586336 218204
rect 586336 218184 586388 218204
rect 586388 218184 586390 218204
rect 586518 218048 586574 218104
rect 591486 217776 591542 217832
rect 591670 217776 591726 217832
rect 591026 217504 591082 217560
rect 590842 217232 590898 217288
rect 591486 217232 591542 217288
rect 592038 216960 592094 217016
rect 590842 216724 590844 216744
rect 590844 216724 590896 216744
rect 590896 216724 590898 216744
rect 590842 216688 590898 216724
rect 591026 216688 591082 216744
rect 582102 215892 582158 215928
rect 582102 215872 582104 215892
rect 582104 215872 582156 215892
rect 582156 215872 582158 215892
rect 586702 215328 586758 215384
rect 578606 213968 578662 214024
rect 579434 211656 579490 211712
rect 578790 209908 578846 209944
rect 578790 209888 578792 209908
rect 578792 209888 578844 209908
rect 578844 209888 578846 209908
rect 597466 222012 597522 222048
rect 597466 221992 597468 222012
rect 597468 221992 597520 222012
rect 597520 221992 597522 222012
rect 599490 221448 599546 221504
rect 599030 220224 599086 220280
rect 597926 217504 597982 217560
rect 595166 216960 595222 217016
rect 595626 216724 595628 216744
rect 595628 216724 595680 216744
rect 595680 216724 595682 216744
rect 595626 216688 595682 216724
rect 595810 216688 595866 216744
rect 595994 216436 596050 216472
rect 595994 216416 595996 216436
rect 595996 216416 596048 216436
rect 596048 216416 596050 216436
rect 595810 215328 595866 215384
rect 595994 215328 596050 215384
rect 595718 215056 595774 215112
rect 597558 216552 597614 216608
rect 598478 217232 598534 217288
rect 599030 216144 599086 216200
rect 602250 221992 602306 222048
rect 600778 221176 600834 221232
rect 599766 219136 599822 219192
rect 601790 220224 601846 220280
rect 600962 218864 601018 218920
rect 600962 218320 601018 218376
rect 601146 218320 601202 218376
rect 601146 217776 601202 217832
rect 600962 216144 601018 216200
rect 600962 215328 601018 215384
rect 604090 219136 604146 219192
rect 606758 220224 606814 220280
rect 606758 219680 606814 219736
rect 616878 221720 616934 221776
rect 611634 220904 611690 220960
rect 611358 215872 611414 215928
rect 614486 218592 614542 218648
rect 617062 219952 617118 220008
rect 620558 215872 620614 215928
rect 618902 215600 618958 215656
rect 626446 218048 626502 218104
rect 630954 219680 631010 219736
rect 630770 219408 630826 219464
rect 629942 218320 629998 218376
rect 631138 218592 631194 218648
rect 652206 298424 652262 298480
rect 640246 231376 640302 231432
rect 639602 230016 639658 230072
rect 638866 219136 638922 219192
rect 640062 218864 640118 218920
rect 650642 223080 650698 223136
rect 643190 220360 643246 220416
rect 641442 220088 641498 220144
rect 642086 217232 642142 217288
rect 643006 215872 643062 215928
rect 642178 213152 642234 213208
rect 644938 217504 644994 217560
rect 646594 215600 646650 215656
rect 649906 218592 649962 218648
rect 647146 214512 647202 214568
rect 651838 222808 651894 222864
rect 651194 221448 651250 221504
rect 651010 214784 651066 214840
rect 579434 207304 579490 207360
rect 578238 205828 578294 205864
rect 578238 205808 578240 205828
rect 578240 205808 578292 205828
rect 578292 205808 578294 205828
rect 660302 405592 660358 405648
rect 659106 360032 659162 360088
rect 666466 742736 666522 742792
rect 666282 705472 666338 705528
rect 667754 786664 667810 786720
rect 667570 743144 667626 743200
rect 667202 671064 667258 671120
rect 668398 783808 668454 783864
rect 668214 752256 668270 752312
rect 668214 733624 668270 733680
rect 667754 710776 667810 710832
rect 667754 688880 667810 688936
rect 667570 665896 667626 665952
rect 666466 665352 666522 665408
rect 665822 626048 665878 626104
rect 664442 579672 664498 579728
rect 666466 603064 666522 603120
rect 668398 708736 668454 708792
rect 668398 692824 668454 692880
rect 668214 662496 668270 662552
rect 668214 654200 668270 654256
rect 667754 621152 667810 621208
rect 668950 773744 669006 773800
rect 668766 734304 668822 734360
rect 668766 731448 668822 731504
rect 668582 670520 668638 670576
rect 671158 872208 671214 872264
rect 670606 867856 670662 867912
rect 669778 864184 669834 864240
rect 669594 789384 669650 789440
rect 669226 755112 669282 755168
rect 669410 741104 669466 741160
rect 668950 709960 669006 710016
rect 669226 705064 669282 705120
rect 668766 664536 668822 664592
rect 669042 648624 669098 648680
rect 668398 620200 668454 620256
rect 668398 601704 668454 601760
rect 668214 574096 668270 574152
rect 668214 564440 668270 564496
rect 667202 534112 667258 534168
rect 666466 529896 666522 529952
rect 664626 493992 664682 494048
rect 662050 491952 662106 492008
rect 661866 406272 661922 406328
rect 663062 315424 663118 315480
rect 661682 268096 661738 268152
rect 666006 494672 666062 494728
rect 668858 593680 668914 593736
rect 668582 535880 668638 535936
rect 669042 573144 669098 573200
rect 669042 559000 669098 559056
rect 668858 528536 668914 528592
rect 668398 526496 668454 526552
rect 668214 485152 668270 485208
rect 665822 358672 665878 358728
rect 664442 271088 664498 271144
rect 663246 234096 663302 234152
rect 658922 233824 658978 233880
rect 661682 229472 661738 229528
rect 660946 229200 661002 229256
rect 652758 226344 652814 226400
rect 654782 225528 654838 225584
rect 653034 220632 653090 220688
rect 655886 225256 655942 225312
rect 655426 216416 655482 216472
rect 660210 224984 660266 225040
rect 658186 224440 658242 224496
rect 656622 223624 656678 223680
rect 658002 221720 658058 221776
rect 659566 223896 659622 223952
rect 658922 223352 658978 223408
rect 661498 213424 661554 213480
rect 663062 231784 663118 231840
rect 663246 231104 663302 231160
rect 664442 230560 664498 230616
rect 664626 215056 664682 215112
rect 664810 213696 664866 213752
rect 665546 230832 665602 230888
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 579526 198872 579582 198928
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 579526 192208 579582 192264
rect 589462 191664 589518 191720
rect 579526 190712 579582 190768
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 579526 187992 579582 188048
rect 589462 186768 589518 186824
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 589462 185136 589518 185192
rect 579526 184320 579582 184376
rect 589462 183504 589518 183560
rect 579526 181872 579582 181928
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 578790 180104 578846 180160
rect 589462 178608 589518 178664
rect 579526 177656 579582 177712
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 579526 171012 579582 171048
rect 579526 170992 579528 171012
rect 579528 170992 579580 171012
rect 579580 170992 579582 171012
rect 578330 169224 578386 169280
rect 578974 166912 579030 166968
rect 578882 164464 578938 164520
rect 579434 162424 579490 162480
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589462 170448 589518 170504
rect 579250 159840 579306 159896
rect 579158 158208 579214 158264
rect 579526 155916 579582 155952
rect 579526 155896 579528 155916
rect 579528 155896 579580 155916
rect 579580 155896 579582 155916
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 578238 153992 578294 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147192 579582 147248
rect 578606 142976 578662 143032
rect 578698 138760 578754 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589462 157412 589518 157448
rect 589462 157392 589464 157412
rect 589464 157392 589516 157412
rect 589516 157392 589518 157412
rect 579526 140564 579528 140584
rect 579528 140564 579580 140584
rect 579580 140564 579582 140584
rect 579526 140528 579582 140564
rect 578882 136584 578938 136640
rect 578330 134408 578386 134464
rect 578238 132232 578294 132288
rect 578330 127744 578386 127800
rect 579526 129684 579528 129704
rect 579528 129684 579580 129704
rect 579580 129684 579582 129704
rect 579526 129648 579582 129684
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 589462 150864 589518 150920
rect 589186 149232 589242 149288
rect 579250 125296 579306 125352
rect 579250 123528 579306 123584
rect 579066 121116 579068 121136
rect 579068 121116 579120 121136
rect 579120 121116 579122 121136
rect 579066 121080 579122 121116
rect 578514 118360 578570 118416
rect 578330 108332 578332 108352
rect 578332 108332 578384 108352
rect 578384 108332 578386 108352
rect 578330 108296 578386 108332
rect 578330 105848 578386 105904
rect 578514 93064 578570 93120
rect 578514 86400 578570 86456
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579526 114436 579582 114472
rect 579526 114416 579528 114436
rect 579528 114416 579580 114436
rect 579580 114416 579582 114436
rect 579526 112648 579582 112704
rect 579434 110236 579436 110256
rect 579436 110236 579488 110256
rect 579488 110236 579490 110256
rect 579434 110200 579490 110236
rect 579526 103300 579528 103320
rect 579528 103300 579580 103320
rect 579580 103300 579582 103320
rect 579526 103264 579582 103300
rect 579250 101768 579306 101824
rect 579526 99204 579582 99240
rect 579526 99184 579528 99204
rect 579528 99184 579580 99204
rect 579580 99184 579582 99204
rect 579526 97452 579528 97472
rect 579528 97452 579580 97472
rect 579580 97452 579582 97472
rect 579526 97416 579582 97452
rect 579526 95004 579528 95024
rect 579528 95004 579580 95024
rect 579580 95004 579582 95024
rect 579526 94968 579582 95004
rect 579066 90888 579122 90944
rect 578882 80008 578938 80064
rect 579526 88032 579582 88088
rect 579342 83988 579344 84008
rect 579344 83988 579396 84008
rect 579396 83988 579398 84008
rect 579342 83952 579398 83988
rect 579250 82184 579306 82240
rect 579066 77832 579122 77888
rect 578606 73108 578608 73128
rect 578608 73108 578660 73128
rect 578660 73108 578662 73128
rect 578606 73072 578662 73108
rect 578514 61784 578570 61840
rect 579250 75556 579252 75576
rect 579252 75556 579304 75576
rect 579304 75556 579306 75576
rect 579250 75520 579306 75556
rect 589370 147600 589426 147656
rect 589462 145968 589518 146024
rect 589922 144336 589978 144392
rect 589462 142704 589518 142760
rect 589094 141072 589150 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589278 136176 589334 136232
rect 589462 134544 589518 134600
rect 588542 132912 588598 132968
rect 579066 71304 579122 71360
rect 579526 68040 579582 68096
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579526 64504 579582 64560
rect 579526 60288 579582 60344
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 579526 56072 579582 56128
rect 581642 54984 581698 55040
rect 590106 131280 590162 131336
rect 589462 129648 589518 129704
rect 589462 128016 589518 128072
rect 589462 124752 589518 124808
rect 589462 123120 589518 123176
rect 589462 121508 589518 121544
rect 589462 121488 589464 121508
rect 589464 121488 589516 121508
rect 589516 121488 589518 121508
rect 590290 126384 590346 126440
rect 589922 119856 589978 119912
rect 588726 118224 588782 118280
rect 589462 116592 589518 116648
rect 589646 114960 589702 115016
rect 589554 113328 589610 113384
rect 589462 111696 589518 111752
rect 589278 110064 589334 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589462 105168 589518 105224
rect 667202 313656 667258 313712
rect 667018 223352 667074 223408
rect 666834 223080 666890 223136
rect 667018 222128 667074 222184
rect 666834 219408 666890 219464
rect 666466 215328 666522 215384
rect 666466 200912 666522 200968
rect 666190 186904 666246 186960
rect 667018 214512 667074 214568
rect 666834 174800 666890 174856
rect 667386 181328 667442 181384
rect 669042 483112 669098 483168
rect 669778 750896 669834 750952
rect 669778 738520 669834 738576
rect 669594 709552 669650 709608
rect 669594 695136 669650 695192
rect 669410 663584 669466 663640
rect 670330 782992 670386 783048
rect 670146 780544 670202 780600
rect 670146 710368 670202 710424
rect 670974 781088 671030 781144
rect 670606 751712 670662 751768
rect 670790 750080 670846 750136
rect 671342 763000 671398 763056
rect 673182 934632 673238 934688
rect 674194 957072 674250 957128
rect 673366 932592 673422 932648
rect 672998 930552 673054 930608
rect 675206 966048 675262 966104
rect 675758 965096 675814 965152
rect 675206 963600 675262 963656
rect 675390 963328 675446 963384
rect 674930 962512 674986 962568
rect 674654 962104 674710 962160
rect 674378 933000 674434 933056
rect 675482 962784 675538 962840
rect 675390 962104 675446 962160
rect 675206 959248 675262 959304
rect 675114 958704 675170 958760
rect 675298 957752 675354 957808
rect 675758 957752 675814 957808
rect 675482 957072 675538 957128
rect 675758 956392 675814 956448
rect 675022 954488 675078 954544
rect 674838 953400 674894 953456
rect 674654 932184 674710 932240
rect 674194 930144 674250 930200
rect 671986 928240 672042 928296
rect 671802 758648 671858 758704
rect 671526 758240 671582 758296
rect 671158 752528 671214 752584
rect 671158 737024 671214 737080
rect 671066 730496 671122 730552
rect 670790 727912 670846 727968
rect 670790 712408 670846 712464
rect 670330 707512 670386 707568
rect 670606 699760 670662 699816
rect 670330 687384 670386 687440
rect 669962 673104 670018 673160
rect 669778 666168 669834 666224
rect 669778 645360 669834 645416
rect 669594 620608 669650 620664
rect 669962 644816 670018 644872
rect 669778 574912 669834 574968
rect 669962 571512 670018 571568
rect 669410 570288 669466 570344
rect 669778 556144 669834 556200
rect 669594 553424 669650 553480
rect 669410 500928 669466 500984
rect 670974 706696 671030 706752
rect 670974 685480 671030 685536
rect 670790 667664 670846 667720
rect 671158 662360 671214 662416
rect 670790 623872 670846 623928
rect 670422 619384 670478 619440
rect 670422 618160 670478 618216
rect 670606 607280 670662 607336
rect 670330 598848 670386 598904
rect 670146 537784 670202 537840
rect 669778 483520 669834 483576
rect 669594 482296 669650 482352
rect 669226 456184 669282 456240
rect 671158 640464 671214 640520
rect 670974 619792 671030 619848
rect 671710 757832 671766 757888
rect 671710 757424 671766 757480
rect 671526 713632 671582 713688
rect 671526 713224 671582 713280
rect 672538 873568 672594 873624
rect 672354 784352 672410 784408
rect 672170 770616 672226 770672
rect 672170 733896 672226 733952
rect 671986 732808 672042 732864
rect 671710 712816 671766 712872
rect 671986 688608 672042 688664
rect 671618 668480 671674 668536
rect 671802 668072 671858 668128
rect 671526 667256 671582 667312
rect 671342 627816 671398 627872
rect 671618 624416 671674 624472
rect 671802 623464 671858 623520
rect 671710 623056 671766 623112
rect 671434 622648 671490 622704
rect 670790 578992 670846 579048
rect 670790 578584 670846 578640
rect 671250 594768 671306 594824
rect 671066 577768 671122 577824
rect 670790 569472 670846 569528
rect 670974 535064 671030 535120
rect 670606 529624 670662 529680
rect 670330 528128 670386 528184
rect 671066 533432 671122 533488
rect 671066 532888 671122 532944
rect 671434 579808 671490 579864
rect 671526 579400 671582 579456
rect 673366 929464 673422 929520
rect 672998 870032 673054 870088
rect 672722 760280 672778 760336
rect 672722 759872 672778 759928
rect 672538 754160 672594 754216
rect 672538 738248 672594 738304
rect 673182 759056 673238 759112
rect 672998 755384 673054 755440
rect 672906 751304 672962 751360
rect 672354 709144 672410 709200
rect 672446 670112 672502 670168
rect 672446 669840 672502 669896
rect 672170 661544 672226 661600
rect 672170 638696 672226 638752
rect 672078 616664 672134 616720
rect 672078 614896 672134 614952
rect 671710 578176 671766 578232
rect 671710 576136 671766 576192
rect 671710 555192 671766 555248
rect 671434 534656 671490 534712
rect 671526 534384 671582 534440
rect 671250 525680 671306 525736
rect 671526 490864 671582 490920
rect 671066 489232 671122 489288
rect 671710 485968 671766 486024
rect 672814 715264 672870 715320
rect 672814 714856 672870 714912
rect 675390 953400 675446 953456
rect 675206 951360 675262 951416
rect 675850 951360 675906 951416
rect 675206 951088 675262 951144
rect 675022 934224 675078 934280
rect 677506 951496 677562 951552
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 676494 938032 676550 938088
rect 676034 937760 676090 937816
rect 675206 933816 675262 933872
rect 678242 950680 678298 950736
rect 678242 935584 678298 935640
rect 683118 947280 683174 947336
rect 683118 939664 683174 939720
rect 682382 935176 682438 935232
rect 681002 933544 681058 933600
rect 677506 931096 677562 931152
rect 683118 929056 683174 929112
rect 675298 879144 675354 879200
rect 675758 875880 675814 875936
rect 675390 873976 675446 874032
rect 675390 873568 675446 873624
rect 675114 873160 675170 873216
rect 675390 872208 675446 872264
rect 674930 870848 674986 870904
rect 675114 870032 675170 870088
rect 673918 864864 673974 864920
rect 673734 779184 673790 779240
rect 673550 777416 673606 777472
rect 673366 732808 673422 732864
rect 673918 771976 673974 772032
rect 674470 788024 674526 788080
rect 674286 779864 674342 779920
rect 673918 752120 673974 752176
rect 673366 730088 673422 730144
rect 673366 728476 673422 728512
rect 673366 728456 673368 728476
rect 673368 728456 673420 728476
rect 673420 728456 673422 728476
rect 673182 714448 673238 714504
rect 672998 714040 673054 714096
rect 673182 698264 673238 698320
rect 672998 685752 673054 685808
rect 672814 669432 672870 669488
rect 672814 668888 672870 668944
rect 672630 662360 672686 662416
rect 672630 661136 672686 661192
rect 672446 625096 672502 625152
rect 672446 604288 672502 604344
rect 672170 574504 672226 574560
rect 672262 532616 672318 532672
rect 672814 635432 672870 635488
rect 672814 622240 672870 622296
rect 673826 728184 673882 728240
rect 673826 727640 673882 727696
rect 674148 727912 674204 727968
rect 675298 868400 675354 868456
rect 674838 868128 674894 868184
rect 674838 867448 674894 867504
rect 675482 867856 675538 867912
rect 675482 867448 675538 867504
rect 675390 864864 675446 864920
rect 675482 864184 675538 864240
rect 674930 789384 674986 789440
rect 675298 863096 675354 863152
rect 674930 787480 674986 787536
rect 674838 787208 674894 787264
rect 675482 788024 675538 788080
rect 675482 787480 675538 787536
rect 675390 787208 675446 787264
rect 675482 786664 675538 786720
rect 675482 784352 675538 784408
rect 675482 783808 675538 783864
rect 675482 782992 675538 783048
rect 675298 781088 675354 781144
rect 675482 780544 675538 780600
rect 675482 779864 675538 779920
rect 675482 779184 675538 779240
rect 675482 778776 675538 778832
rect 675482 777416 675538 777472
rect 675574 775648 675630 775704
rect 675758 775512 675814 775568
rect 675022 774560 675078 774616
rect 675114 774288 675170 774344
rect 674838 768168 674894 768224
rect 675390 773744 675446 773800
rect 682382 772656 682438 772712
rect 675114 766536 675170 766592
rect 674654 757152 674710 757208
rect 676034 763000 676090 763056
rect 677046 761912 677102 761968
rect 676770 761776 676826 761832
rect 676034 760688 676090 760744
rect 676034 757172 676090 757208
rect 676034 757152 676036 757172
rect 676036 757152 676088 757172
rect 676088 757152 676090 757172
rect 675850 755792 675906 755848
rect 683210 771976 683266 772032
rect 683394 770888 683450 770944
rect 682382 757016 682438 757072
rect 677046 754976 677102 755032
rect 676770 754568 676826 754624
rect 683578 770616 683634 770672
rect 683578 759464 683634 759520
rect 683302 756608 683358 756664
rect 683486 753752 683542 753808
rect 683118 752936 683174 752992
rect 675114 743144 675170 743200
rect 674930 742736 674986 742792
rect 675390 742464 675446 742520
rect 675114 741512 675170 741568
rect 674930 741104 674986 741160
rect 675114 739608 675170 739664
rect 675022 738520 675078 738576
rect 675206 738316 675262 738372
rect 675114 737024 675170 737080
rect 674286 726824 674342 726880
rect 674930 734304 674986 734360
rect 675114 733896 675170 733952
rect 675114 733624 675170 733680
rect 675114 731448 675170 731504
rect 675482 730496 675538 730552
rect 675298 730088 675354 730144
rect 674746 727640 674802 727696
rect 683486 726824 683542 726880
rect 674010 726552 674066 726608
rect 674562 726552 674618 726608
rect 682382 725736 682438 725792
rect 673550 724104 673606 724160
rect 673550 689560 673606 689616
rect 673366 666440 673422 666496
rect 673366 660728 673422 660784
rect 673366 659912 673422 659968
rect 673182 620880 673238 620936
rect 672998 615712 673054 615768
rect 673090 604560 673146 604616
rect 672814 577360 672870 577416
rect 672814 576952 672870 577008
rect 672906 559408 672962 559464
rect 672814 548392 672870 548448
rect 672630 546216 672686 546272
rect 672630 533840 672686 533896
rect 672446 528944 672502 529000
rect 673182 530576 673238 530632
rect 672722 490048 672778 490104
rect 672446 489640 672502 489696
rect 671986 455368 672042 455424
rect 670882 455096 670938 455152
rect 671986 455116 672042 455152
rect 671986 455096 671988 455116
rect 671988 455096 672040 455116
rect 672040 455096 672042 455116
rect 672262 453736 672318 453792
rect 669962 403688 670018 403744
rect 670606 393488 670662 393544
rect 668766 360848 668822 360904
rect 669962 347248 670018 347304
rect 668582 312840 668638 312896
rect 668306 302232 668362 302288
rect 668582 234504 668638 234560
rect 668122 230852 668178 230888
rect 668122 230832 668124 230852
rect 668124 230832 668176 230852
rect 668176 230832 668178 230852
rect 667938 229744 667994 229800
rect 668398 224984 668454 225040
rect 668398 223624 668454 223680
rect 668398 220360 668454 220416
rect 668398 219816 668454 219872
rect 667938 192480 667994 192536
rect 667938 189252 667940 189272
rect 667940 189252 667992 189272
rect 667992 189252 667994 189272
rect 667938 189216 667994 189252
rect 668122 182688 668178 182744
rect 667754 178744 667810 178800
rect 667938 174564 667940 174584
rect 667940 174564 667992 174584
rect 667992 174564 667994 174584
rect 667938 174528 667994 174564
rect 668030 169668 668032 169688
rect 668032 169668 668084 169688
rect 668084 169668 668086 169688
rect 668030 169632 668086 169668
rect 667938 164772 667940 164792
rect 667940 164772 667992 164792
rect 667992 164772 667994 164792
rect 667938 164736 667994 164772
rect 668306 163104 668362 163160
rect 668950 236680 669006 236736
rect 669410 230852 669466 230888
rect 669410 230832 669412 230852
rect 669412 230832 669464 230852
rect 669464 230832 669466 230852
rect 669410 226344 669466 226400
rect 669410 225664 669466 225720
rect 669410 216416 669466 216472
rect 669410 214104 669466 214160
rect 669318 199044 669320 199064
rect 669320 199044 669372 199064
rect 669372 199044 669374 199064
rect 669318 199008 669374 199044
rect 669134 197376 669190 197432
rect 669410 197104 669466 197160
rect 669226 196016 669282 196072
rect 669410 194148 669412 194168
rect 669412 194148 669464 194168
rect 669464 194148 669466 194168
rect 669410 194112 669466 194148
rect 669226 187584 669282 187640
rect 669226 184320 669282 184376
rect 669778 168136 669834 168192
rect 669134 164192 669190 164248
rect 668950 159840 669006 159896
rect 668766 153312 668822 153368
rect 668766 149096 668822 149152
rect 668490 148416 668546 148472
rect 668490 145152 668546 145208
rect 667570 135904 667626 135960
rect 668030 135360 668086 135416
rect 667202 134544 667258 134600
rect 667018 133048 667074 133104
rect 669134 138624 669190 138680
rect 668950 128288 669006 128344
rect 668766 125568 668822 125624
rect 670422 257624 670478 257680
rect 670422 235864 670478 235920
rect 670146 232872 670202 232928
rect 672630 488008 672686 488064
rect 672446 401648 672502 401704
rect 672446 400424 672502 400480
rect 672906 485560 672962 485616
rect 676034 718256 676090 718312
rect 676034 715672 676090 715728
rect 683302 724104 683358 724160
rect 682382 711592 682438 711648
rect 683302 707920 683358 707976
rect 683670 726416 683726 726472
rect 683854 725464 683910 725520
rect 683670 711184 683726 711240
rect 683854 708328 683910 708384
rect 683486 707104 683542 707160
rect 674378 706288 674434 706344
rect 674010 693504 674066 693560
rect 673734 680992 673790 681048
rect 673734 647808 673790 647864
rect 673550 636792 673606 636848
rect 673550 603472 673606 603528
rect 674194 690104 674250 690160
rect 674930 699760 674986 699816
rect 675114 698264 675170 698320
rect 675390 696768 675446 696824
rect 675114 695136 675170 695192
rect 675666 694320 675722 694376
rect 675114 693504 675170 693560
rect 675114 692824 675170 692880
rect 675390 690104 675446 690160
rect 675298 689560 675354 689616
rect 674930 688880 674986 688936
rect 675298 688880 675354 688936
rect 675114 688608 675170 688664
rect 674838 686432 674894 686488
rect 675482 687384 675538 687440
rect 675482 685752 675538 685808
rect 675206 685480 675262 685536
rect 674838 670112 674894 670168
rect 674838 669432 674894 669488
rect 683210 682624 683266 682680
rect 676494 673104 676550 673160
rect 676494 671064 676550 671120
rect 676494 666168 676550 666224
rect 676494 665352 676550 665408
rect 683670 682352 683726 682408
rect 683486 680992 683542 681048
rect 683210 664536 683266 664592
rect 683670 666984 683726 667040
rect 683486 662904 683542 662960
rect 675390 654200 675446 654256
rect 675574 652840 675630 652896
rect 675390 651480 675446 651536
rect 675206 649712 675262 649768
rect 675390 648896 675446 648952
rect 674470 647536 674526 647592
rect 674378 645088 674434 645144
rect 674194 641688 674250 641744
rect 673918 618568 673974 618624
rect 674010 599120 674066 599176
rect 673826 598440 673882 598496
rect 674838 647536 674894 647592
rect 675022 647264 675078 647320
rect 675482 648624 675538 648680
rect 675482 647808 675538 647864
rect 675482 645360 675538 645416
rect 675390 644816 675446 644872
rect 675758 644272 675814 644328
rect 675206 644000 675262 644056
rect 675206 643728 675262 643784
rect 675482 643456 675538 643512
rect 675298 641688 675354 641744
rect 674838 640736 674894 640792
rect 674378 624824 674434 624880
rect 674378 606464 674434 606520
rect 674194 592864 674250 592920
rect 673734 591096 673790 591152
rect 674194 552064 674250 552120
rect 674010 545672 674066 545728
rect 674010 535336 674066 535392
rect 674010 534112 674066 534168
rect 673826 532208 673882 532264
rect 673826 531800 673882 531856
rect 673642 528400 673698 528456
rect 673366 488416 673422 488472
rect 673090 484744 673146 484800
rect 675390 640464 675446 640520
rect 674930 631352 674986 631408
rect 674746 617344 674802 617400
rect 674838 603200 674894 603256
rect 675022 601704 675078 601760
rect 674838 601024 674894 601080
rect 675022 600480 675078 600536
rect 675022 599664 675078 599720
rect 674838 598848 674894 598904
rect 674838 598032 674894 598088
rect 675022 596808 675078 596864
rect 675482 638696 675538 638752
rect 675390 638016 675446 638072
rect 677506 637880 677562 637936
rect 675758 637608 675814 637664
rect 674930 595448 674986 595504
rect 674562 592592 674618 592648
rect 675758 631352 675814 631408
rect 675850 627816 675906 627872
rect 676494 625640 676550 625696
rect 683302 636792 683358 636848
rect 683118 624824 683174 624880
rect 677506 621968 677562 622024
rect 683670 635432 683726 635488
rect 683670 624416 683726 624472
rect 683302 617888 683358 617944
rect 683118 617072 683174 617128
rect 675482 607688 675538 607744
rect 675482 607280 675538 607336
rect 675482 606464 675538 606520
rect 675482 604560 675538 604616
rect 675482 604288 675538 604344
rect 675482 603472 675538 603528
rect 675482 602928 675538 602984
rect 675482 601024 675538 601080
rect 675482 600480 675538 600536
rect 675482 599120 675538 599176
rect 675482 598440 675538 598496
rect 675482 598032 675538 598088
rect 675482 596808 675538 596864
rect 675390 595448 675446 595504
rect 675482 594768 675538 594824
rect 675390 593680 675446 593736
rect 683302 592864 683358 592920
rect 675758 592320 675814 592376
rect 675574 592048 675630 592104
rect 674654 558320 674710 558376
rect 674378 547032 674434 547088
rect 674470 535064 674526 535120
rect 674470 534112 674526 534168
rect 674838 556144 674894 556200
rect 674838 554784 674894 554840
rect 675574 586200 675630 586256
rect 683118 592592 683174 592648
rect 676034 582936 676090 582992
rect 676034 580216 676090 580272
rect 675758 576544 675814 576600
rect 682382 575592 682438 575648
rect 683118 573960 683174 574016
rect 683486 591096 683542 591152
rect 683302 573144 683358 573200
rect 683486 572328 683542 572384
rect 683118 570696 683174 570752
rect 675206 564440 675262 564496
rect 675390 563080 675446 563136
rect 675482 561176 675538 561232
rect 675298 559408 675354 559464
rect 675298 559000 675354 559056
rect 675390 558320 675446 558376
rect 675298 557504 675354 557560
rect 675390 555192 675446 555248
rect 675298 554784 675354 554840
rect 675298 553968 675354 554024
rect 675390 553424 675446 553480
rect 675390 552064 675446 552120
rect 675758 550704 675814 550760
rect 675114 549616 675170 549672
rect 674838 547576 674894 547632
rect 674838 545944 674894 546000
rect 675482 549616 675538 549672
rect 675482 548392 675538 548448
rect 675850 547596 675906 547632
rect 675850 547576 675852 547596
rect 675852 547576 675904 547596
rect 675904 547576 675906 547596
rect 675298 546488 675354 546544
rect 674930 503784 674986 503840
rect 676402 546216 676458 546272
rect 676034 537784 676090 537840
rect 676034 535676 676090 535732
rect 675758 529624 675814 529680
rect 675758 529148 675814 529204
rect 675022 503512 675078 503568
rect 675022 503240 675078 503296
rect 675850 503784 675906 503840
rect 676034 503532 676090 503568
rect 676034 503512 676036 503532
rect 676036 503512 676088 503532
rect 676088 503512 676090 503532
rect 676034 503240 676090 503296
rect 674930 500928 674986 500984
rect 674654 484336 674710 484392
rect 674194 483928 674250 483984
rect 674746 464752 674802 464808
rect 673826 456864 673882 456920
rect 674746 456864 674802 456920
rect 673946 456204 674002 456240
rect 673946 456184 673948 456204
rect 673948 456184 674000 456204
rect 674000 456184 674002 456204
rect 673596 455660 673652 455696
rect 673596 455640 673598 455660
rect 673598 455640 673650 455660
rect 673650 455640 673652 455660
rect 673504 455388 673560 455424
rect 673504 455368 673506 455388
rect 673506 455368 673558 455388
rect 673558 455368 673560 455388
rect 673386 455132 673388 455152
rect 673388 455132 673440 455152
rect 673440 455132 673442 455152
rect 673386 455096 673442 455132
rect 675298 486376 675354 486432
rect 673162 454844 673218 454880
rect 673162 454824 673164 454844
rect 673164 454824 673216 454844
rect 673216 454824 673218 454844
rect 674930 454824 674986 454880
rect 683210 547032 683266 547088
rect 679622 546488 679678 546544
rect 678242 531392 678298 531448
rect 683394 545672 683450 545728
rect 683210 531800 683266 531856
rect 679622 530984 679678 531040
rect 683578 532208 683634 532264
rect 683394 527720 683450 527776
rect 683578 526496 683634 526552
rect 676862 525680 676918 525736
rect 677874 524456 677930 524512
rect 683210 503648 683266 503704
rect 676034 493992 676090 494048
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 675482 454552 675538 454608
rect 675850 481888 675906 481944
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 675666 454280 675722 454336
rect 672814 454044 672816 454064
rect 672816 454044 672868 454064
rect 672868 454044 672870 454064
rect 672814 454008 672870 454044
rect 676034 480664 676090 480720
rect 677322 492360 677378 492416
rect 677322 487192 677378 487248
rect 681002 487600 681058 487656
rect 679622 486784 679678 486840
rect 683578 494672 683634 494728
rect 683394 491680 683450 491736
rect 683578 491272 683634 491328
rect 683210 482704 683266 482760
rect 682382 481480 682438 481536
rect 676770 455640 676826 455696
rect 676034 454008 676090 454064
rect 675850 453736 675906 453792
rect 683118 406272 683174 406328
rect 676034 405592 676090 405648
rect 676034 403416 676090 403472
rect 683118 403280 683174 403336
rect 674654 402192 674710 402248
rect 674194 401376 674250 401432
rect 672630 400016 672686 400072
rect 673182 398792 673238 398848
rect 672998 397160 673054 397216
rect 672630 393896 672686 393952
rect 672814 392536 672870 392592
rect 672630 376216 672686 376272
rect 672446 355816 672502 355872
rect 672446 355408 672502 355464
rect 672262 351328 672318 351384
rect 671986 348880 672042 348936
rect 672262 335280 672318 335336
rect 671986 332288 672042 332344
rect 672630 348472 672686 348528
rect 672446 310800 672502 310856
rect 671986 301960 672042 302016
rect 671342 269728 671398 269784
rect 671526 264016 671582 264072
rect 671342 262112 671398 262168
rect 671342 244704 671398 244760
rect 671802 258848 671858 258904
rect 671802 241440 671858 241496
rect 671526 238176 671582 238232
rect 671066 227160 671122 227216
rect 671066 226616 671122 226672
rect 671066 225664 671122 225720
rect 671066 225392 671122 225448
rect 670928 224440 670984 224496
rect 670882 224032 670938 224088
rect 670698 223932 670700 223952
rect 670700 223932 670752 223952
rect 670752 223932 670754 223952
rect 670698 223896 670754 223932
rect 670698 220360 670754 220416
rect 670698 219816 670754 219872
rect 670606 211112 670662 211168
rect 670606 210840 670662 210896
rect 671802 229472 671858 229528
rect 672630 256944 672686 257000
rect 672170 234504 672226 234560
rect 672170 231376 672226 231432
rect 672262 227024 672318 227080
rect 672262 226480 672318 226536
rect 671986 226344 672042 226400
rect 671802 225936 671858 225992
rect 670606 190304 670662 190360
rect 670606 170312 670662 170368
rect 670330 165552 670386 165608
rect 669594 122712 669650 122768
rect 669226 121352 669282 121408
rect 668950 120672 669006 120728
rect 668214 119040 668270 119096
rect 668030 117408 668086 117464
rect 671986 224984 672042 225040
rect 672262 224984 672318 225040
rect 671802 221720 671858 221776
rect 671802 220904 671858 220960
rect 672262 224712 672318 224768
rect 672262 224032 672318 224088
rect 671986 219816 672042 219872
rect 672170 214784 672226 214840
rect 672078 213696 672134 213752
rect 672078 200640 672134 200696
rect 672262 196016 672318 196072
rect 672078 183504 672134 183560
rect 671894 176432 671950 176488
rect 671894 166912 671950 166968
rect 671710 158208 671766 158264
rect 671526 150048 671582 150104
rect 670606 147600 670662 147656
rect 671342 131688 671398 131744
rect 669226 114144 669282 114200
rect 671526 130872 671582 130928
rect 668214 112512 668270 112568
rect 668306 111832 668362 111888
rect 668030 109248 668086 109304
rect 666650 105984 666706 106040
rect 667202 105984 667258 106040
rect 590106 103536 590162 103592
rect 589462 101904 589518 101960
rect 585782 77832 585838 77888
rect 584402 54712 584458 54768
rect 635738 96600 635794 96656
rect 637026 96600 637082 96656
rect 626446 95376 626502 95432
rect 643190 95104 643246 95160
rect 626262 94424 626318 94480
rect 626446 93472 626502 93528
rect 625618 92520 625674 92576
rect 625434 91568 625490 91624
rect 626446 90616 626502 90672
rect 625250 89664 625306 89720
rect 643374 89664 643430 89720
rect 626446 88848 626502 88904
rect 626446 87896 626502 87952
rect 643558 87080 643614 87136
rect 625618 86944 625674 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 625618 84124 625620 84144
rect 625620 84124 625672 84144
rect 625672 84124 625674 84144
rect 625618 84088 625674 84124
rect 624422 82864 624478 82920
rect 644938 92112 644994 92168
rect 644754 84632 644810 84688
rect 643742 82728 643798 82784
rect 628654 81640 628710 81696
rect 629206 80824 629262 80880
rect 633898 80416 633954 80472
rect 639602 77832 639658 77888
rect 655242 94152 655298 94208
rect 655058 93336 655114 93392
rect 654874 92520 654930 92576
rect 654138 90616 654194 90672
rect 655426 91432 655482 91488
rect 663246 93064 663302 93120
rect 655794 89800 655850 89856
rect 663706 91976 663762 92032
rect 664166 88984 664222 89040
rect 647054 74432 647110 74488
rect 646870 72936 646926 72992
rect 647330 69944 647386 70000
rect 646226 68856 646282 68912
rect 648986 71440 649042 71496
rect 649170 66952 649226 67008
rect 647514 65456 647570 65512
rect 646134 64368 646190 64424
rect 604458 54440 604514 54496
rect 580262 54168 580318 54224
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 308034 50224 308090 50280
rect 461904 52808 461960 52864
rect 465722 52808 465778 52864
rect 309690 49680 309746 49736
rect 458178 46960 458234 47016
rect 458362 46688 458418 46744
rect 431222 44784 431278 44840
rect 142618 44240 142674 44296
rect 310426 44104 310482 44160
rect 364890 44104 364946 44160
rect 308954 42744 309010 42800
rect 194322 42064 194378 42120
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 419906 41792 419962 41848
rect 443550 42200 443606 42256
rect 443550 41520 443606 41576
rect 460110 44784 460166 44840
rect 460846 43424 460902 43480
rect 461950 44376 462006 44432
rect 462502 44376 462558 44432
rect 463698 44104 463754 44160
rect 462962 43832 463018 43888
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463698 42880 463754 42936
rect 544014 47504 544070 47560
rect 549994 48864 550050 48920
rect 553674 50224 553730 50280
rect 552018 48048 552074 48104
rect 547878 47776 547934 47832
rect 665178 93336 665234 93392
rect 665362 90616 665418 90672
rect 664626 89800 664682 89856
rect 672602 230288 672658 230344
rect 672998 377984 673054 378040
rect 673366 396344 673422 396400
rect 673826 396072 673882 396128
rect 673366 382200 673422 382256
rect 674010 395664 674066 395720
rect 673826 381384 673882 381440
rect 674010 375400 674066 375456
rect 674470 394440 674526 394496
rect 674470 377712 674526 377768
rect 676034 399336 676090 399392
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675114 377712 675170 377768
rect 675206 377440 675262 377496
rect 675758 377168 675814 377224
rect 675390 376216 675446 376272
rect 675390 375400 675446 375456
rect 675758 372952 675814 373008
rect 675114 372544 675170 372600
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 357448 674710 357504
rect 674654 357040 674710 357096
rect 674194 356632 674250 356688
rect 674102 356224 674158 356280
rect 673182 355000 673238 355056
rect 672998 354592 673054 354648
rect 673182 353368 673238 353424
rect 673918 352552 673974 352608
rect 673550 352144 673606 352200
rect 673366 349696 673422 349752
rect 673182 340720 673238 340776
rect 673366 335824 673422 335880
rect 673734 350512 673790 350568
rect 673918 336640 673974 336696
rect 673734 331064 673790 331120
rect 673550 325624 673606 325680
rect 673918 312024 673974 312080
rect 673182 311208 673238 311264
rect 672998 309984 673054 310040
rect 672998 304272 673054 304328
rect 672998 287816 673054 287872
rect 673734 305496 673790 305552
rect 673366 304680 673422 304736
rect 673366 289992 673422 290048
rect 673734 285504 673790 285560
rect 674470 349424 674526 349480
rect 674286 347656 674342 347712
rect 676034 353776 676090 353832
rect 675942 349152 675998 349208
rect 675114 340720 675170 340776
rect 675758 340312 675814 340368
rect 675390 338952 675446 339008
rect 674470 332832 674526 332888
rect 674286 327528 674342 327584
rect 675574 337728 675630 337784
rect 675114 336640 675170 336696
rect 675758 336640 675814 336696
rect 675482 335824 675538 335880
rect 675298 335280 675354 335336
rect 675390 332832 675446 332888
rect 675114 332288 675170 332344
rect 675758 332152 675814 332208
rect 675114 331064 675170 331120
rect 675758 328344 675814 328400
rect 675114 327528 675170 327584
rect 675114 325624 675170 325680
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 312432 674710 312488
rect 674102 311616 674158 311672
rect 674470 310392 674526 310448
rect 674194 309576 674250 309632
rect 673918 267416 673974 267472
rect 673182 266464 673238 266520
rect 674010 266192 674066 266248
rect 673182 263744 673238 263800
rect 672998 260072 673054 260128
rect 672998 244976 673054 245032
rect 674838 309168 674894 309224
rect 674654 303864 674710 303920
rect 676034 308352 676090 308408
rect 675022 307944 675078 308000
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 676402 305904 676458 305960
rect 676034 303456 676090 303512
rect 674838 298016 674894 298072
rect 675298 298016 675354 298072
rect 674838 296792 674894 296848
rect 675022 296520 675078 296576
rect 676034 301960 676090 302016
rect 676678 305088 676734 305144
rect 676402 301552 676458 301608
rect 676678 301416 676734 301472
rect 678978 306312 679034 306368
rect 678242 297336 678298 297392
rect 676126 296792 676182 296848
rect 675942 296520 675998 296576
rect 675758 296248 675814 296304
rect 675758 295840 675814 295896
rect 675758 295160 675814 295216
rect 675758 291488 675814 291544
rect 675114 289992 675170 290048
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 683118 271088 683174 271144
rect 676034 269728 676090 269784
rect 676034 268232 676090 268288
rect 683118 268096 683174 268152
rect 674654 267008 674710 267064
rect 674470 265784 674526 265840
rect 674378 265376 674434 265432
rect 674194 264968 674250 265024
rect 673734 259664 673790 259720
rect 673366 259256 673422 259312
rect 673918 258440 673974 258496
rect 673734 245520 673790 245576
rect 673366 242800 673422 242856
rect 673526 236700 673582 236736
rect 673526 236680 673528 236700
rect 673528 236680 673580 236700
rect 673580 236680 673582 236700
rect 673182 233144 673238 233200
rect 673182 232872 673238 232928
rect 672998 231376 673054 231432
rect 673366 230288 673422 230344
rect 673090 229744 673146 229800
rect 673090 229472 673146 229528
rect 673458 230016 673514 230072
rect 673458 229084 673514 229120
rect 673458 229064 673460 229084
rect 673460 229064 673512 229084
rect 673512 229064 673514 229084
rect 673504 228828 673506 228848
rect 673506 228828 673558 228848
rect 673558 228828 673560 228848
rect 673504 228792 673560 228828
rect 672906 228656 672962 228712
rect 673386 228540 673442 228576
rect 673386 228520 673388 228540
rect 673388 228520 673440 228540
rect 673440 228520 673442 228540
rect 673182 226752 673238 226808
rect 673182 225120 673238 225176
rect 672906 224576 672962 224632
rect 672722 224304 672778 224360
rect 672814 220360 672870 220416
rect 673504 225392 673560 225448
rect 674286 260888 674342 260944
rect 674286 246880 674342 246936
rect 674102 235184 674158 235240
rect 674470 234912 674526 234968
rect 674838 264424 674894 264480
rect 676494 264016 676550 264072
rect 674838 263744 674894 263800
rect 676494 263608 676550 263664
rect 678242 263200 678298 263256
rect 676218 262792 676274 262848
rect 674930 251504 674986 251560
rect 674930 249328 674986 249384
rect 678426 261160 678482 261216
rect 675850 251540 675852 251560
rect 675852 251540 675904 251560
rect 675904 251540 675906 251560
rect 675850 251504 675906 251540
rect 675758 250280 675814 250336
rect 675390 249600 675446 249656
rect 675114 246880 675170 246936
rect 675114 245520 675170 245576
rect 674838 245248 674894 245304
rect 675114 242800 675170 242856
rect 675114 241440 675170 241496
rect 675206 240216 675262 240272
rect 675114 238176 675170 238232
rect 675390 236816 675446 236872
rect 675114 235864 675170 235920
rect 675666 235184 675722 235240
rect 674654 234368 674710 234424
rect 675850 234912 675906 234968
rect 675850 234388 675906 234424
rect 675850 234368 675852 234388
rect 675852 234368 675904 234388
rect 675904 234368 675906 234388
rect 675178 231804 675234 231840
rect 675178 231784 675180 231804
rect 675180 231784 675232 231804
rect 675232 231784 675234 231804
rect 674954 231276 674956 231296
rect 674956 231276 675008 231296
rect 675008 231276 675010 231296
rect 674954 231240 675010 231276
rect 674838 231140 674840 231160
rect 674840 231140 674892 231160
rect 674892 231140 674894 231160
rect 675850 231260 675906 231296
rect 675850 231240 675852 231260
rect 675852 231240 675904 231260
rect 675904 231240 675906 231260
rect 674838 231104 674894 231140
rect 674730 230868 674732 230888
rect 674732 230868 674784 230888
rect 674784 230868 674786 230888
rect 674730 230832 674786 230868
rect 674516 230288 674572 230344
rect 675022 230560 675078 230616
rect 676770 230288 676826 230344
rect 674056 230016 674112 230072
rect 675114 230016 675170 230072
rect 673826 223624 673882 223680
rect 673918 222808 673974 222864
rect 673734 220632 673790 220688
rect 673366 216144 673422 216200
rect 672722 214648 672778 214704
rect 672906 209888 672962 209944
rect 672446 177792 672502 177848
rect 672538 175208 672594 175264
rect 672354 169088 672410 169144
rect 672354 153040 672410 153096
rect 672078 140256 672134 140312
rect 672722 149096 672778 149152
rect 672538 130464 672594 130520
rect 672354 124344 672410 124400
rect 671894 115776 671950 115832
rect 673550 212880 673606 212936
rect 673550 206896 673606 206952
rect 673366 201864 673422 201920
rect 673550 201592 673606 201648
rect 673366 174392 673422 174448
rect 673090 172896 673146 172952
rect 673182 169904 673238 169960
rect 673182 151680 673238 151736
rect 673918 209616 673974 209672
rect 673918 203224 673974 203280
rect 675114 229472 675170 229528
rect 675114 229064 675170 229120
rect 675114 228792 675170 228848
rect 675022 227024 675078 227080
rect 674286 225664 674342 225720
rect 674562 221856 674618 221912
rect 674378 220224 674434 220280
rect 674102 179424 674158 179480
rect 674194 176840 674250 176896
rect 674010 168680 674066 168736
rect 673734 168408 673790 168464
rect 674010 151000 674066 151056
rect 675206 226072 675262 226128
rect 675022 221448 675078 221504
rect 674930 220496 674986 220552
rect 674746 218592 674802 218648
rect 675390 224848 675446 224904
rect 675850 224576 675906 224632
rect 675390 222128 675446 222184
rect 675850 220496 675906 220552
rect 676034 219988 676036 220008
rect 676036 219988 676088 220008
rect 676088 219988 676090 220008
rect 676034 219952 676090 219988
rect 676034 219716 676036 219736
rect 676036 219716 676088 219736
rect 676088 219716 676090 219736
rect 676034 219680 676090 219716
rect 674930 217504 674986 217560
rect 674930 216824 674986 216880
rect 674746 216552 674802 216608
rect 674930 215872 674986 215928
rect 675298 219136 675354 219192
rect 675666 219000 675722 219056
rect 675298 215736 675354 215792
rect 675114 215600 675170 215656
rect 675022 212880 675078 212936
rect 674746 204992 674802 205048
rect 676034 217776 676090 217832
rect 675850 215092 675852 215112
rect 675852 215092 675904 215112
rect 675904 215092 675906 215112
rect 675850 215056 675906 215092
rect 675850 213424 675906 213480
rect 675850 213188 675852 213208
rect 675852 213188 675904 213208
rect 675904 213188 675906 213208
rect 675850 213152 675906 213188
rect 675666 212880 675722 212936
rect 676862 209616 676918 209672
rect 676126 207168 676182 207224
rect 679254 223760 679310 223816
rect 683854 234096 683910 234152
rect 683302 233824 683358 233880
rect 683302 223080 683358 223136
rect 679990 222264 680046 222320
rect 679806 221448 679862 221504
rect 679622 220632 679678 220688
rect 683854 222672 683910 222728
rect 683486 219816 683542 219872
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 677782 206896 677838 206952
rect 675758 205536 675814 205592
rect 675482 204992 675538 205048
rect 674838 202680 674894 202736
rect 675390 202680 675446 202736
rect 675482 201864 675538 201920
rect 675022 200912 675078 200968
rect 675206 200640 675262 200696
rect 675758 200640 675814 200696
rect 675574 198192 675630 198248
rect 675390 197104 675446 197160
rect 675758 197104 675814 197160
rect 675666 193160 675722 193216
rect 675758 191528 675814 191584
rect 675298 190304 675354 190360
rect 683118 186904 683174 186960
rect 676494 181328 676550 181384
rect 676034 178064 676090 178120
rect 683118 178744 683174 178800
rect 674562 177248 674618 177304
rect 674654 176024 674710 176080
rect 674378 175616 674434 175672
rect 674378 169496 674434 169552
rect 674378 155352 674434 155408
rect 674194 132096 674250 132152
rect 678242 173168 678298 173224
rect 674838 172760 674894 172816
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 676586 166368 676642 166424
rect 676034 165552 676090 165608
rect 681002 171536 681058 171592
rect 679622 171128 679678 171184
rect 675942 161880 675998 161936
rect 676126 161336 676182 161392
rect 675758 160656 675814 160712
rect 675758 159296 675814 159352
rect 674838 157528 674894 157584
rect 675482 157528 675538 157584
rect 675390 156984 675446 157040
rect 675758 156304 675814 156360
rect 675114 155352 675170 155408
rect 675114 153040 675170 153096
rect 675758 153040 675814 153096
rect 675114 151680 675170 151736
rect 675114 151000 675170 151056
rect 675666 148416 675722 148472
rect 675114 147600 675170 147656
rect 675666 147600 675722 147656
rect 675758 145968 675814 146024
rect 683118 135904 683174 135960
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 683118 132640 683174 132696
rect 674654 131280 674710 131336
rect 675942 130056 675998 130112
rect 673366 129648 673422 129704
rect 674102 129240 674158 129296
rect 673274 125976 673330 126032
rect 672906 123936 672962 123992
rect 673090 123936 673146 123992
rect 672814 123120 672870 123176
rect 672814 121352 672870 121408
rect 672538 121080 672594 121136
rect 673366 123528 673422 123584
rect 672538 110880 672594 110936
rect 672354 110200 672410 110256
rect 671526 107616 671582 107672
rect 673090 111424 673146 111480
rect 672814 106392 672870 106448
rect 674286 128288 674342 128344
rect 675942 128288 675998 128344
rect 674102 111832 674158 111888
rect 673366 105576 673422 105632
rect 668306 104352 668362 104408
rect 682382 127744 682438 127800
rect 674838 127608 674894 127664
rect 674654 125568 674710 125624
rect 674470 125160 674526 125216
rect 675022 126384 675078 126440
rect 675298 113056 675354 113112
rect 675114 111424 675170 111480
rect 674654 110200 674710 110256
rect 675666 108024 675722 108080
rect 675114 106392 675170 106448
rect 675758 106120 675814 106176
rect 675114 105576 675170 105632
rect 675758 103128 675814 103184
rect 675666 102584 675722 102640
rect 668490 102176 668546 102232
rect 674286 102176 674342 102232
rect 675758 101360 675814 101416
rect 663982 48456 664038 48512
rect 663798 47776 663854 47832
rect 662418 47368 662474 47424
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40432 141754 40488
<< metal3 >>
rect 106825 1007314 106891 1007317
rect 106628 1007312 106891 1007314
rect 106628 1007256 106830 1007312
rect 106886 1007256 106891 1007312
rect 106628 1007254 106891 1007256
rect 106825 1007251 106891 1007254
rect 425513 1007178 425579 1007181
rect 425513 1007176 425776 1007178
rect 425513 1007120 425518 1007176
rect 425574 1007120 425776 1007176
rect 425513 1007118 425776 1007120
rect 425513 1007115 425579 1007118
rect 359733 1007042 359799 1007045
rect 359628 1007040 359799 1007042
rect 359628 1006984 359738 1007040
rect 359794 1006984 359799 1007040
rect 359628 1006982 359799 1006984
rect 359733 1006979 359799 1006982
rect 359365 1006906 359431 1006909
rect 428365 1006906 428431 1006909
rect 507853 1006906 507919 1006909
rect 359168 1006904 359431 1006906
rect 359168 1006848 359370 1006904
rect 359426 1006848 359431 1006904
rect 359168 1006846 359431 1006848
rect 428260 1006904 428431 1006906
rect 428260 1006848 428370 1006904
rect 428426 1006848 428431 1006904
rect 428260 1006846 428431 1006848
rect 507656 1006904 507919 1006906
rect 507656 1006848 507858 1006904
rect 507914 1006848 507919 1006904
rect 507656 1006846 507919 1006848
rect 359365 1006843 359431 1006846
rect 428365 1006843 428431 1006846
rect 507853 1006843 507919 1006846
rect 361389 1006770 361455 1006773
rect 429193 1006770 429259 1006773
rect 505001 1006770 505067 1006773
rect 555969 1006770 556035 1006773
rect 361192 1006768 361455 1006770
rect 361192 1006712 361394 1006768
rect 361450 1006712 361455 1006768
rect 361192 1006710 361455 1006712
rect 428996 1006768 429259 1006770
rect 428996 1006712 429198 1006768
rect 429254 1006712 429259 1006768
rect 428996 1006710 429259 1006712
rect 504804 1006768 505067 1006770
rect 504804 1006712 505006 1006768
rect 505062 1006712 505067 1006768
rect 504804 1006710 505067 1006712
rect 555772 1006768 556035 1006770
rect 555772 1006712 555974 1006768
rect 556030 1006712 556035 1006768
rect 555772 1006710 556035 1006712
rect 361389 1006707 361455 1006710
rect 429193 1006707 429259 1006710
rect 505001 1006707 505067 1006710
rect 555969 1006707 556035 1006710
rect 101949 1006634 102015 1006637
rect 153745 1006634 153811 1006637
rect 157425 1006634 157491 1006637
rect 101949 1006632 102212 1006634
rect 101949 1006576 101954 1006632
rect 102010 1006576 102212 1006632
rect 101949 1006574 102212 1006576
rect 153548 1006632 153811 1006634
rect 153548 1006576 153750 1006632
rect 153806 1006576 153811 1006632
rect 153548 1006574 153811 1006576
rect 157228 1006632 157491 1006634
rect 157228 1006576 157430 1006632
rect 157486 1006576 157491 1006632
rect 157228 1006574 157491 1006576
rect 101949 1006571 102015 1006574
rect 153745 1006571 153811 1006574
rect 157425 1006571 157491 1006574
rect 431677 1006634 431743 1006637
rect 501321 1006634 501387 1006637
rect 556797 1006634 556863 1006637
rect 431677 1006632 431940 1006634
rect 431677 1006576 431682 1006632
rect 431738 1006576 431940 1006632
rect 431677 1006574 431940 1006576
rect 501124 1006632 501387 1006634
rect 501124 1006576 501326 1006632
rect 501382 1006576 501387 1006632
rect 501124 1006574 501387 1006576
rect 556600 1006632 556863 1006634
rect 556600 1006576 556802 1006632
rect 556858 1006576 556863 1006632
rect 556600 1006574 556863 1006576
rect 431677 1006571 431743 1006574
rect 501321 1006571 501387 1006574
rect 556797 1006571 556863 1006574
rect 104801 1006498 104867 1006501
rect 152917 1006498 152983 1006501
rect 158253 1006498 158319 1006501
rect 256141 1006498 256207 1006501
rect 104604 1006496 104867 1006498
rect 104604 1006440 104806 1006496
rect 104862 1006440 104867 1006496
rect 104604 1006438 104867 1006440
rect 152720 1006496 152983 1006498
rect 152720 1006440 152922 1006496
rect 152978 1006440 152983 1006496
rect 152720 1006438 152983 1006440
rect 158056 1006496 158319 1006498
rect 158056 1006440 158258 1006496
rect 158314 1006440 158319 1006496
rect 158056 1006438 158319 1006440
rect 255944 1006496 256207 1006498
rect 255944 1006440 256146 1006496
rect 256202 1006440 256207 1006496
rect 255944 1006438 256207 1006440
rect 104801 1006435 104867 1006438
rect 152917 1006435 152983 1006438
rect 158253 1006435 158319 1006438
rect 256141 1006435 256207 1006438
rect 307753 1006498 307819 1006501
rect 360561 1006498 360627 1006501
rect 429193 1006498 429259 1006501
rect 553117 1006498 553183 1006501
rect 307753 1006496 307924 1006498
rect 307753 1006440 307758 1006496
rect 307814 1006440 307924 1006496
rect 307753 1006438 307924 1006440
rect 360561 1006496 360824 1006498
rect 360561 1006440 360566 1006496
rect 360622 1006440 360824 1006496
rect 360561 1006438 360824 1006440
rect 429193 1006496 429456 1006498
rect 429193 1006440 429198 1006496
rect 429254 1006440 429456 1006496
rect 429193 1006438 429456 1006440
rect 552920 1006496 553183 1006498
rect 552920 1006440 553122 1006496
rect 553178 1006440 553183 1006496
rect 552920 1006438 553183 1006440
rect 307753 1006435 307819 1006438
rect 360561 1006435 360627 1006438
rect 429193 1006435 429259 1006438
rect 553117 1006435 553183 1006438
rect 100293 1006362 100359 1006365
rect 158621 1006362 158687 1006365
rect 258993 1006362 259059 1006365
rect 100293 1006360 100556 1006362
rect 100293 1006304 100298 1006360
rect 100354 1006304 100556 1006360
rect 100293 1006302 100556 1006304
rect 158621 1006360 158884 1006362
rect 158621 1006304 158626 1006360
rect 158682 1006304 158884 1006360
rect 158621 1006302 158884 1006304
rect 258796 1006360 259059 1006362
rect 258796 1006304 258998 1006360
rect 259054 1006304 259059 1006360
rect 258796 1006302 259059 1006304
rect 100293 1006299 100359 1006302
rect 158621 1006299 158687 1006302
rect 258993 1006299 259059 1006302
rect 306925 1006362 306991 1006365
rect 314653 1006362 314719 1006365
rect 423489 1006362 423555 1006365
rect 505369 1006362 505435 1006365
rect 552289 1006362 552355 1006365
rect 306925 1006360 307188 1006362
rect 306925 1006304 306930 1006360
rect 306986 1006304 307188 1006360
rect 306925 1006302 307188 1006304
rect 314548 1006360 314719 1006362
rect 314548 1006304 314658 1006360
rect 314714 1006304 314719 1006360
rect 314548 1006302 314719 1006304
rect 423292 1006360 423555 1006362
rect 423292 1006304 423494 1006360
rect 423550 1006304 423555 1006360
rect 423292 1006302 423555 1006304
rect 505172 1006360 505435 1006362
rect 505172 1006304 505374 1006360
rect 505430 1006304 505435 1006360
rect 505172 1006302 505435 1006304
rect 552092 1006360 552355 1006362
rect 552092 1006304 552294 1006360
rect 552350 1006304 552355 1006360
rect 552092 1006302 552355 1006304
rect 306925 1006299 306991 1006302
rect 314653 1006299 314719 1006302
rect 423489 1006299 423555 1006302
rect 505369 1006299 505435 1006302
rect 552289 1006299 552355 1006302
rect 103973 1006226 104039 1006229
rect 105997 1006226 106063 1006229
rect 103973 1006224 104236 1006226
rect 103973 1006168 103978 1006224
rect 104034 1006168 104236 1006224
rect 103973 1006166 104236 1006168
rect 105892 1006224 106063 1006226
rect 105892 1006168 106002 1006224
rect 106058 1006168 106063 1006224
rect 105892 1006166 106063 1006168
rect 103973 1006163 104039 1006166
rect 105997 1006163 106063 1006166
rect 151261 1006226 151327 1006229
rect 152089 1006226 152155 1006229
rect 160277 1006226 160343 1006229
rect 210417 1006226 210483 1006229
rect 262673 1006226 262739 1006229
rect 151261 1006224 151524 1006226
rect 151261 1006168 151266 1006224
rect 151322 1006168 151524 1006224
rect 151261 1006166 151524 1006168
rect 152089 1006224 152352 1006226
rect 152089 1006168 152094 1006224
rect 152150 1006168 152352 1006224
rect 152089 1006166 152352 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 210220 1006224 210483 1006226
rect 210220 1006168 210422 1006224
rect 210478 1006168 210483 1006224
rect 210220 1006166 210483 1006168
rect 262476 1006224 262739 1006226
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 151261 1006163 151327 1006166
rect 152089 1006163 152155 1006166
rect 160277 1006163 160343 1006166
rect 210417 1006163 210483 1006166
rect 262673 1006163 262739 1006166
rect 304901 1006226 304967 1006229
rect 357709 1006226 357775 1006229
rect 365069 1006226 365135 1006229
rect 507025 1006226 507091 1006229
rect 304901 1006224 305164 1006226
rect 304901 1006168 304906 1006224
rect 304962 1006168 305164 1006224
rect 304901 1006166 305164 1006168
rect 357604 1006224 357775 1006226
rect 357604 1006168 357714 1006224
rect 357770 1006168 357775 1006224
rect 357604 1006166 357775 1006168
rect 364872 1006224 365135 1006226
rect 364872 1006168 365074 1006224
rect 365130 1006168 365135 1006224
rect 364872 1006166 365135 1006168
rect 506828 1006224 507091 1006226
rect 506828 1006168 507030 1006224
rect 507086 1006168 507091 1006224
rect 506828 1006166 507091 1006168
rect 304901 1006163 304967 1006166
rect 357709 1006163 357775 1006166
rect 365069 1006163 365135 1006166
rect 507025 1006163 507091 1006166
rect 551461 1006226 551527 1006229
rect 551461 1006224 551724 1006226
rect 551461 1006168 551466 1006224
rect 551522 1006168 551724 1006224
rect 551461 1006166 551724 1006168
rect 551461 1006163 551527 1006166
rect 98269 1006090 98335 1006093
rect 102317 1006090 102383 1006093
rect 108481 1006090 108547 1006093
rect 98269 1006088 98900 1006090
rect 98269 1006032 98274 1006088
rect 98330 1006032 98900 1006088
rect 98269 1006030 98900 1006032
rect 102317 1006088 102580 1006090
rect 102317 1006032 102322 1006088
rect 102378 1006032 102580 1006088
rect 102317 1006030 102580 1006032
rect 108284 1006088 108547 1006090
rect 108284 1006032 108486 1006088
rect 108542 1006032 108547 1006088
rect 108284 1006030 108547 1006032
rect 98269 1006027 98335 1006030
rect 102317 1006027 102383 1006030
rect 108481 1006027 108547 1006030
rect 147121 1006090 147187 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 158253 1006090 158319 1006093
rect 159449 1006090 159515 1006093
rect 201033 1006090 201099 1006093
rect 208393 1006090 208459 1006093
rect 252461 1006090 252527 1006093
rect 257337 1006090 257403 1006093
rect 261845 1006090 261911 1006093
rect 147121 1006088 148935 1006090
rect 147121 1006032 147126 1006088
rect 147182 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 147121 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 158253 1006088 158516 1006090
rect 158253 1006032 158258 1006088
rect 158314 1006032 158516 1006088
rect 158253 1006030 158516 1006032
rect 159449 1006088 159712 1006090
rect 159449 1006032 159454 1006088
rect 159510 1006032 159712 1006088
rect 159449 1006030 159712 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 208393 1006088 208656 1006090
rect 208393 1006032 208398 1006088
rect 208454 1006032 208656 1006088
rect 208393 1006030 208656 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 257337 1006088 257600 1006090
rect 257337 1006032 257342 1006088
rect 257398 1006032 257600 1006088
rect 257337 1006030 257600 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 147121 1006027 147187 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 158253 1006027 158319 1006030
rect 159449 1006027 159515 1006030
rect 201033 1006027 201099 1006030
rect 208393 1006027 208459 1006030
rect 252461 1006027 252527 1006030
rect 257337 1006027 257403 1006030
rect 261845 1006027 261911 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 354857 1006090 354923 1006093
rect 355685 1006090 355751 1006093
rect 363413 1006090 363479 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314653 1006088 314916 1006090
rect 314653 1006032 314658 1006088
rect 314714 1006032 314916 1006088
rect 314653 1006030 314916 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 355685 1006088 355948 1006090
rect 355685 1006032 355690 1006088
rect 355746 1006032 355948 1006088
rect 355685 1006030 355948 1006032
rect 363308 1006088 363479 1006090
rect 363308 1006032 363418 1006088
rect 363474 1006032 363479 1006088
rect 363308 1006030 363479 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 354857 1006027 354923 1006030
rect 355685 1006027 355751 1006030
rect 363413 1006027 363479 1006030
rect 421833 1006090 421899 1006093
rect 423489 1006090 423555 1006093
rect 431677 1006090 431743 1006093
rect 421833 1006088 422556 1006090
rect 421833 1006032 421838 1006088
rect 421894 1006032 422556 1006088
rect 421833 1006030 422556 1006032
rect 423489 1006088 423752 1006090
rect 423489 1006032 423494 1006088
rect 423550 1006032 423752 1006088
rect 423489 1006030 423752 1006032
rect 431480 1006088 431743 1006090
rect 431480 1006032 431682 1006088
rect 431738 1006032 431743 1006088
rect 431480 1006030 431743 1006032
rect 421833 1006027 421899 1006030
rect 423489 1006027 423555 1006030
rect 431677 1006027 431743 1006030
rect 498837 1006090 498903 1006093
rect 502517 1006090 502583 1006093
rect 506197 1006090 506263 1006093
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 502517 1006088 502780 1006090
rect 502517 1006032 502522 1006088
rect 502578 1006032 502780 1006088
rect 502517 1006030 502780 1006032
rect 506000 1006088 506263 1006090
rect 506000 1006032 506202 1006088
rect 506258 1006032 506263 1006088
rect 506000 1006030 506263 1006032
rect 498837 1006027 498903 1006030
rect 502517 1006027 502583 1006030
rect 506197 1006027 506263 1006030
rect 509049 1006090 509115 1006093
rect 551093 1006090 551159 1006093
rect 509049 1006088 509312 1006090
rect 509049 1006032 509054 1006088
rect 509110 1006032 509312 1006088
rect 509049 1006030 509312 1006032
rect 550436 1006088 551159 1006090
rect 550436 1006032 551098 1006088
rect 551154 1006032 551159 1006088
rect 550436 1006030 551159 1006032
rect 509049 1006027 509115 1006030
rect 551093 1006027 551159 1006030
rect 555969 1006090 556035 1006093
rect 555969 1006088 556232 1006090
rect 555969 1006032 555974 1006088
rect 556030 1006032 556232 1006088
rect 555969 1006030 556232 1006032
rect 555969 1006027 556035 1006030
rect 426341 1005682 426407 1005685
rect 426144 1005680 426407 1005682
rect 426144 1005624 426346 1005680
rect 426402 1005624 426407 1005680
rect 426144 1005622 426407 1005624
rect 426341 1005619 426407 1005622
rect 425513 1005546 425579 1005549
rect 425316 1005544 425579 1005546
rect 425316 1005488 425518 1005544
rect 425574 1005488 425579 1005544
rect 425316 1005486 425579 1005488
rect 425513 1005483 425579 1005486
rect 360561 1005410 360627 1005413
rect 424317 1005410 424383 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 424120 1005408 424383 1005410
rect 424120 1005352 424322 1005408
rect 424378 1005352 424383 1005408
rect 424120 1005350 424383 1005352
rect 360561 1005347 360627 1005350
rect 424317 1005347 424383 1005350
rect 552289 1005410 552355 1005413
rect 552289 1005408 552552 1005410
rect 552289 1005352 552294 1005408
rect 552350 1005352 552552 1005408
rect 552289 1005350 552552 1005352
rect 552289 1005347 552355 1005350
rect 108849 1005274 108915 1005277
rect 212073 1005274 212139 1005277
rect 108849 1005272 109112 1005274
rect 108849 1005216 108854 1005272
rect 108910 1005216 109112 1005272
rect 108849 1005214 109112 1005216
rect 211876 1005272 212139 1005274
rect 211876 1005216 212078 1005272
rect 212134 1005216 212139 1005272
rect 211876 1005214 212139 1005216
rect 108849 1005211 108915 1005214
rect 212073 1005211 212139 1005214
rect 307293 1005274 307359 1005277
rect 356513 1005274 356579 1005277
rect 425145 1005274 425211 1005277
rect 498837 1005274 498903 1005277
rect 551461 1005274 551527 1005277
rect 307293 1005272 307556 1005274
rect 307293 1005216 307298 1005272
rect 307354 1005216 307556 1005272
rect 307293 1005214 307556 1005216
rect 356316 1005272 356579 1005274
rect 356316 1005216 356518 1005272
rect 356574 1005216 356579 1005272
rect 356316 1005214 356579 1005216
rect 424948 1005272 425211 1005274
rect 424948 1005216 425150 1005272
rect 425206 1005216 425211 1005272
rect 424948 1005214 425211 1005216
rect 498732 1005272 498903 1005274
rect 498732 1005216 498842 1005272
rect 498898 1005216 498903 1005272
rect 498732 1005214 498903 1005216
rect 551356 1005272 551527 1005274
rect 551356 1005216 551466 1005272
rect 551522 1005216 551527 1005272
rect 551356 1005214 551527 1005216
rect 307293 1005211 307359 1005214
rect 356513 1005211 356579 1005214
rect 425145 1005211 425211 1005214
rect 498837 1005211 498903 1005214
rect 551461 1005211 551527 1005214
rect 152917 1005138 152983 1005141
rect 258165 1005138 258231 1005141
rect 308949 1005138 309015 1005141
rect 152917 1005136 153180 1005138
rect 152917 1005080 152922 1005136
rect 152978 1005080 153180 1005136
rect 152917 1005078 153180 1005080
rect 258165 1005136 258428 1005138
rect 258165 1005080 258170 1005136
rect 258226 1005080 258428 1005136
rect 258165 1005078 258428 1005080
rect 308752 1005136 309015 1005138
rect 308752 1005080 308954 1005136
rect 309010 1005080 309015 1005136
rect 308752 1005078 309015 1005080
rect 152917 1005075 152983 1005078
rect 258165 1005075 258231 1005078
rect 308949 1005075 309015 1005078
rect 365069 1005138 365135 1005141
rect 508221 1005138 508287 1005141
rect 365069 1005136 365332 1005138
rect 365069 1005080 365074 1005136
rect 365130 1005080 365332 1005136
rect 365069 1005078 365332 1005080
rect 508221 1005136 508484 1005138
rect 508221 1005080 508226 1005136
rect 508282 1005080 508484 1005136
rect 508221 1005078 508484 1005080
rect 365069 1005075 365135 1005078
rect 508221 1005075 508287 1005078
rect 153745 1005002 153811 1005005
rect 209221 1005002 209287 1005005
rect 263041 1005002 263107 1005005
rect 355685 1005002 355751 1005005
rect 153745 1005000 153916 1005002
rect 153745 1004944 153750 1005000
rect 153806 1004944 153916 1005000
rect 153745 1004942 153916 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 262844 1005000 263107 1005002
rect 262844 1004944 263046 1005000
rect 263102 1004944 263107 1005000
rect 262844 1004942 263107 1004944
rect 355488 1005000 355751 1005002
rect 355488 1004944 355690 1005000
rect 355746 1004944 355751 1005000
rect 355488 1004942 355751 1004944
rect 153745 1004939 153811 1004942
rect 209221 1004939 209287 1004942
rect 263041 1004939 263107 1004942
rect 355685 1004939 355751 1004942
rect 361389 1005002 361455 1005005
rect 427997 1005002 428063 1005005
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 427800 1005000 428063 1005002
rect 427800 1004944 428002 1005000
rect 428058 1004944 428063 1005000
rect 427800 1004942 428063 1004944
rect 361389 1004939 361455 1004942
rect 427997 1004939 428063 1004942
rect 500493 1005002 500559 1005005
rect 500493 1005000 500756 1005002
rect 500493 1004944 500498 1005000
rect 500554 1004944 500756 1005000
rect 500493 1004942 500756 1004944
rect 500493 1004939 500559 1004942
rect 151721 1004866 151787 1004869
rect 160645 1004866 160711 1004869
rect 151721 1004864 151892 1004866
rect 151721 1004808 151726 1004864
rect 151782 1004808 151892 1004864
rect 151721 1004806 151892 1004808
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 151721 1004803 151787 1004806
rect 160645 1004803 160711 1004806
rect 211245 1004866 211311 1004869
rect 258165 1004866 258231 1004869
rect 211245 1004864 211508 1004866
rect 211245 1004808 211250 1004864
rect 211306 1004808 211508 1004864
rect 211245 1004806 211508 1004808
rect 257968 1004864 258231 1004866
rect 257968 1004808 258170 1004864
rect 258226 1004808 258231 1004864
rect 257968 1004806 258231 1004808
rect 211245 1004803 211311 1004806
rect 258165 1004803 258231 1004806
rect 308121 1004866 308187 1004869
rect 313825 1004866 313891 1004869
rect 308121 1004864 308384 1004866
rect 308121 1004808 308126 1004864
rect 308182 1004808 308384 1004864
rect 308121 1004806 308384 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 308121 1004803 308187 1004806
rect 313825 1004803 313891 1004806
rect 356513 1004866 356579 1004869
rect 362585 1004866 362651 1004869
rect 356513 1004864 356684 1004866
rect 356513 1004808 356518 1004864
rect 356574 1004808 356684 1004864
rect 356513 1004806 356684 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 356513 1004803 356579 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 499665 1004866 499731 1004869
rect 508221 1004866 508287 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 499665 1004864 499928 1004866
rect 499665 1004808 499670 1004864
rect 499726 1004808 499928 1004864
rect 499665 1004806 499928 1004808
rect 508116 1004864 508287 1004866
rect 508116 1004808 508226 1004864
rect 508282 1004808 508287 1004864
rect 508116 1004806 508287 1004808
rect 422661 1004803 422727 1004806
rect 499665 1004803 499731 1004806
rect 508221 1004803 508287 1004806
rect 108481 1004730 108547 1004733
rect 154113 1004730 154179 1004733
rect 161105 1004730 161171 1004733
rect 209221 1004730 209287 1004733
rect 306925 1004730 306991 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 432873 1004730 432939 1004733
rect 500493 1004730 500559 1004733
rect 507393 1004730 507459 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 154113 1004728 154376 1004730
rect 154113 1004672 154118 1004728
rect 154174 1004672 154376 1004728
rect 154113 1004670 154376 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 306728 1004728 306991 1004730
rect 306728 1004672 306930 1004728
rect 306986 1004672 306991 1004728
rect 306728 1004670 306991 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 432676 1004728 432939 1004730
rect 432676 1004672 432878 1004728
rect 432934 1004672 432939 1004728
rect 432676 1004670 432939 1004672
rect 500296 1004728 500559 1004730
rect 500296 1004672 500498 1004728
rect 500554 1004672 500559 1004728
rect 500296 1004670 500559 1004672
rect 507196 1004728 507459 1004730
rect 507196 1004672 507398 1004728
rect 507454 1004672 507459 1004728
rect 507196 1004670 507459 1004672
rect 108481 1004667 108547 1004670
rect 154113 1004667 154179 1004670
rect 161105 1004667 161171 1004670
rect 209221 1004667 209287 1004670
rect 306925 1004667 306991 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 432873 1004667 432939 1004670
rect 500493 1004667 500559 1004670
rect 507393 1004667 507459 1004670
rect 560845 1004730 560911 1004733
rect 560845 1004728 561108 1004730
rect 560845 1004672 560850 1004728
rect 560906 1004672 561108 1004728
rect 560845 1004670 561108 1004672
rect 560845 1004667 560911 1004670
rect 504541 1004458 504607 1004461
rect 504436 1004456 504607 1004458
rect 504436 1004400 504546 1004456
rect 504602 1004400 504607 1004456
rect 504436 1004398 504607 1004400
rect 504541 1004395 504607 1004398
rect 426341 1004050 426407 1004053
rect 426341 1004048 426604 1004050
rect 426341 1003992 426346 1004048
rect 426402 1003992 426604 1004048
rect 426341 1003990 426604 1003992
rect 426341 1003987 426407 1003990
rect 103145 1003914 103211 1003917
rect 255313 1003914 255379 1003917
rect 557165 1003914 557231 1003917
rect 103145 1003912 103408 1003914
rect 103145 1003856 103150 1003912
rect 103206 1003856 103408 1003912
rect 103145 1003854 103408 1003856
rect 255116 1003912 255379 1003914
rect 255116 1003856 255318 1003912
rect 255374 1003856 255379 1003912
rect 255116 1003854 255379 1003856
rect 557060 1003912 557231 1003914
rect 557060 1003856 557170 1003912
rect 557226 1003856 557231 1003912
rect 557060 1003854 557231 1003856
rect 103145 1003851 103211 1003854
rect 255313 1003851 255379 1003854
rect 557165 1003851 557231 1003854
rect 305269 1003370 305335 1003373
rect 501689 1003370 501755 1003373
rect 305269 1003368 305532 1003370
rect 305269 1003312 305274 1003368
rect 305330 1003312 305532 1003368
rect 305269 1003310 305532 1003312
rect 501492 1003368 501755 1003370
rect 501492 1003312 501694 1003368
rect 501750 1003312 501755 1003368
rect 501492 1003310 501755 1003312
rect 305269 1003307 305335 1003310
rect 501689 1003307 501755 1003310
rect 101949 1002690 102015 1002693
rect 101752 1002688 102015 1002690
rect 101752 1002632 101954 1002688
rect 102010 1002632 102015 1002688
rect 101752 1002630 102015 1002632
rect 101949 1002627 102015 1002630
rect 256141 1002690 256207 1002693
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 256141 1002627 256207 1002630
rect 100293 1002554 100359 1002557
rect 100096 1002552 100359 1002554
rect 100096 1002496 100298 1002552
rect 100354 1002496 100359 1002552
rect 100096 1002494 100359 1002496
rect 100293 1002491 100359 1002494
rect 254117 1002554 254183 1002557
rect 261017 1002554 261083 1002557
rect 310605 1002554 310671 1002557
rect 560845 1002554 560911 1002557
rect 254117 1002552 254380 1002554
rect 254117 1002496 254122 1002552
rect 254178 1002496 254380 1002552
rect 254117 1002494 254380 1002496
rect 260820 1002552 261083 1002554
rect 260820 1002496 261022 1002552
rect 261078 1002496 261083 1002552
rect 260820 1002494 261083 1002496
rect 310408 1002552 310671 1002554
rect 310408 1002496 310610 1002552
rect 310666 1002496 310671 1002552
rect 310408 1002494 310671 1002496
rect 560740 1002552 560911 1002554
rect 560740 1002496 560850 1002552
rect 560906 1002496 560911 1002552
rect 560740 1002494 560911 1002496
rect 254117 1002491 254183 1002494
rect 261017 1002491 261083 1002494
rect 310605 1002491 310671 1002494
rect 560845 1002491 560911 1002494
rect 99097 1002418 99163 1002421
rect 107653 1002418 107719 1002421
rect 99097 1002416 99268 1002418
rect 99097 1002360 99102 1002416
rect 99158 1002360 99268 1002416
rect 99097 1002358 99268 1002360
rect 107456 1002416 107719 1002418
rect 107456 1002360 107658 1002416
rect 107714 1002360 107719 1002416
rect 107456 1002358 107719 1002360
rect 99097 1002355 99163 1002358
rect 107653 1002355 107719 1002358
rect 150893 1002418 150959 1002421
rect 254485 1002418 254551 1002421
rect 260189 1002418 260255 1002421
rect 503345 1002418 503411 1002421
rect 150893 1002416 151156 1002418
rect 150893 1002360 150898 1002416
rect 150954 1002360 151156 1002416
rect 150893 1002358 151156 1002360
rect 254485 1002416 254748 1002418
rect 254485 1002360 254490 1002416
rect 254546 1002360 254748 1002416
rect 254485 1002358 254748 1002360
rect 260084 1002416 260255 1002418
rect 260084 1002360 260194 1002416
rect 260250 1002360 260255 1002416
rect 260084 1002358 260255 1002360
rect 503148 1002416 503411 1002418
rect 503148 1002360 503350 1002416
rect 503406 1002360 503411 1002416
rect 503148 1002358 503411 1002360
rect 150893 1002355 150959 1002358
rect 254485 1002355 254551 1002358
rect 260189 1002355 260255 1002358
rect 503345 1002355 503411 1002358
rect 553945 1002418 554011 1002421
rect 560477 1002418 560543 1002421
rect 553945 1002416 554116 1002418
rect 553945 1002360 553950 1002416
rect 554006 1002360 554116 1002416
rect 553945 1002358 554116 1002360
rect 560280 1002416 560543 1002418
rect 560280 1002360 560482 1002416
rect 560538 1002360 560543 1002416
rect 560280 1002358 560543 1002360
rect 553945 1002355 554011 1002358
rect 560477 1002355 560543 1002358
rect 101121 1002282 101187 1002285
rect 105629 1002282 105695 1002285
rect 108021 1002282 108087 1002285
rect 155769 1002282 155835 1002285
rect 206369 1002282 206435 1002285
rect 206737 1002282 206803 1002285
rect 100924 1002280 101187 1002282
rect 100924 1002224 101126 1002280
rect 101182 1002224 101187 1002280
rect 100924 1002222 101187 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 107916 1002280 108087 1002282
rect 107916 1002224 108026 1002280
rect 108082 1002224 108087 1002280
rect 107916 1002222 108087 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 206172 1002280 206435 1002282
rect 206172 1002224 206374 1002280
rect 206430 1002224 206435 1002280
rect 206172 1002222 206435 1002224
rect 206540 1002280 206803 1002282
rect 206540 1002224 206742 1002280
rect 206798 1002224 206803 1002280
rect 206540 1002222 206803 1002224
rect 101121 1002219 101187 1002222
rect 105629 1002219 105695 1002222
rect 108021 1002219 108087 1002222
rect 155769 1002219 155835 1002222
rect 206369 1002219 206435 1002222
rect 206737 1002219 206803 1002222
rect 256509 1002282 256575 1002285
rect 259821 1002282 259887 1002285
rect 256509 1002280 256772 1002282
rect 256509 1002224 256514 1002280
rect 256570 1002224 256772 1002280
rect 256509 1002222 256772 1002224
rect 259624 1002280 259887 1002282
rect 259624 1002224 259826 1002280
rect 259882 1002224 259887 1002280
rect 259624 1002222 259887 1002224
rect 256509 1002219 256575 1002222
rect 259821 1002219 259887 1002222
rect 299381 1002282 299447 1002285
rect 303245 1002282 303311 1002285
rect 306097 1002282 306163 1002285
rect 299381 1002280 303311 1002282
rect 299381 1002224 299386 1002280
rect 299442 1002224 303250 1002280
rect 303306 1002224 303311 1002280
rect 299381 1002222 303311 1002224
rect 305900 1002280 306163 1002282
rect 305900 1002224 306102 1002280
rect 306158 1002224 306163 1002280
rect 305900 1002222 306163 1002224
rect 299381 1002219 299447 1002222
rect 303245 1002219 303311 1002222
rect 306097 1002219 306163 1002222
rect 310605 1002282 310671 1002285
rect 358537 1002282 358603 1002285
rect 310605 1002280 310868 1002282
rect 310605 1002224 310610 1002280
rect 310666 1002224 310868 1002280
rect 310605 1002222 310868 1002224
rect 358340 1002280 358603 1002282
rect 358340 1002224 358542 1002280
rect 358598 1002224 358603 1002280
rect 358340 1002222 358603 1002224
rect 310605 1002219 310671 1002222
rect 358537 1002219 358603 1002222
rect 555141 1002282 555207 1002285
rect 555141 1002280 555404 1002282
rect 555141 1002224 555146 1002280
rect 555202 1002224 555404 1002280
rect 555141 1002222 555404 1002224
rect 555141 1002219 555207 1002222
rect 99465 1002146 99531 1002149
rect 103145 1002146 103211 1002149
rect 99465 1002144 99728 1002146
rect 99465 1002088 99470 1002144
rect 99526 1002088 99728 1002144
rect 99465 1002086 99728 1002088
rect 102948 1002144 103211 1002146
rect 102948 1002088 103150 1002144
rect 103206 1002088 103211 1002144
rect 102948 1002086 103211 1002088
rect 99465 1002083 99531 1002086
rect 103145 1002083 103211 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 154573 1002146 154639 1002149
rect 157793 1002146 157859 1002149
rect 154573 1002144 154836 1002146
rect 154573 1002088 154578 1002144
rect 154634 1002088 154836 1002144
rect 154573 1002086 154836 1002088
rect 157596 1002144 157859 1002146
rect 157596 1002088 157798 1002144
rect 157854 1002088 157859 1002144
rect 157596 1002086 157859 1002088
rect 154573 1002083 154639 1002086
rect 157793 1002083 157859 1002086
rect 207197 1002146 207263 1002149
rect 210877 1002146 210943 1002149
rect 255313 1002146 255379 1002149
rect 261017 1002146 261083 1002149
rect 263501 1002146 263567 1002149
rect 304073 1002146 304139 1002149
rect 207197 1002144 207460 1002146
rect 207197 1002088 207202 1002144
rect 207258 1002088 207460 1002144
rect 207197 1002086 207460 1002088
rect 210877 1002144 211140 1002146
rect 210877 1002088 210882 1002144
rect 210938 1002088 211140 1002144
rect 210877 1002086 211140 1002088
rect 255313 1002144 255576 1002146
rect 255313 1002088 255318 1002144
rect 255374 1002088 255576 1002144
rect 255313 1002086 255576 1002088
rect 261017 1002144 261280 1002146
rect 261017 1002088 261022 1002144
rect 261078 1002088 261280 1002144
rect 261017 1002086 261280 1002088
rect 263304 1002144 263567 1002146
rect 263304 1002088 263506 1002144
rect 263562 1002088 263567 1002144
rect 263304 1002086 263567 1002088
rect 303876 1002144 304139 1002146
rect 303876 1002088 304078 1002144
rect 304134 1002088 304139 1002144
rect 303876 1002086 304139 1002088
rect 207197 1002083 207263 1002086
rect 210877 1002083 210943 1002086
rect 255313 1002083 255379 1002086
rect 261017 1002083 261083 1002086
rect 263501 1002083 263567 1002086
rect 304073 1002083 304139 1002086
rect 357709 1002146 357775 1002149
rect 427169 1002146 427235 1002149
rect 357709 1002144 357972 1002146
rect 357709 1002088 357714 1002144
rect 357770 1002088 357972 1002144
rect 357709 1002086 357972 1002088
rect 426972 1002144 427235 1002146
rect 426972 1002088 427174 1002144
rect 427230 1002088 427235 1002144
rect 426972 1002086 427235 1002088
rect 357709 1002083 357775 1002086
rect 427169 1002083 427235 1002086
rect 503345 1002146 503411 1002149
rect 509877 1002146 509943 1002149
rect 503345 1002144 503608 1002146
rect 503345 1002088 503350 1002144
rect 503406 1002088 503608 1002144
rect 503345 1002086 503608 1002088
rect 509680 1002144 509943 1002146
rect 509680 1002088 509882 1002144
rect 509938 1002088 509943 1002144
rect 509680 1002086 509943 1002088
rect 503345 1002083 503411 1002086
rect 509877 1002083 509943 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101121 1002010 101187 1002013
rect 104801 1002010 104867 1002013
rect 105997 1002010 106063 1002013
rect 149237 1002010 149303 1002013
rect 154941 1002010 155007 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 202689 1002010 202755 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 104801 1002008 104972 1002010
rect 104801 1001952 104806 1002008
rect 104862 1001952 104972 1002008
rect 104801 1001950 104972 1001952
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 155769 1002008 156032 1002010
rect 155769 1001952 155774 1002008
rect 155830 1001952 156032 1002008
rect 155769 1001950 156032 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 202492 1002008 202755 1002010
rect 202492 1001952 202694 1002008
rect 202750 1001952 202755 1002008
rect 202492 1001950 202755 1001952
rect 101121 1001947 101187 1001950
rect 104801 1001947 104867 1001950
rect 105997 1001947 106063 1001950
rect 149237 1001947 149303 1001950
rect 154941 1001947 155007 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 202689 1001947 202755 1001950
rect 205541 1002010 205607 1002013
rect 206737 1002010 206803 1002013
rect 207565 1002010 207631 1002013
rect 212533 1002010 212599 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 206737 1002008 207000 1002010
rect 206737 1001952 206742 1002008
rect 206798 1001952 207000 1002008
rect 206737 1001950 207000 1001952
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 212336 1002008 212599 1002010
rect 212336 1001952 212538 1002008
rect 212594 1001952 212599 1002008
rect 212336 1001950 212599 1001952
rect 205541 1001947 205607 1001950
rect 206737 1001947 206803 1001950
rect 207565 1001947 207631 1001950
rect 212533 1001947 212599 1001950
rect 256969 1002010 257035 1002013
rect 258993 1002010 259059 1002013
rect 260189 1002010 260255 1002013
rect 261845 1002010 261911 1002013
rect 263869 1002010 263935 1002013
rect 256969 1002008 257140 1002010
rect 256969 1001952 256974 1002008
rect 257030 1001952 257140 1002008
rect 256969 1001950 257140 1001952
rect 258993 1002008 259164 1002010
rect 258993 1001952 258998 1002008
rect 259054 1001952 259164 1002008
rect 258993 1001950 259164 1001952
rect 260189 1002008 260452 1002010
rect 260189 1001952 260194 1002008
rect 260250 1001952 260452 1002008
rect 260189 1001950 260452 1001952
rect 261845 1002008 262108 1002010
rect 261845 1001952 261850 1002008
rect 261906 1001952 262108 1002008
rect 261845 1001950 262108 1001952
rect 263764 1002008 263935 1002010
rect 263764 1001952 263874 1002008
rect 263930 1001952 263935 1002008
rect 263764 1001950 263935 1001952
rect 256969 1001947 257035 1001950
rect 258993 1001947 259059 1001950
rect 260189 1001947 260255 1001950
rect 261845 1001947 261911 1001950
rect 263869 1001947 263935 1001950
rect 306097 1002010 306163 1002013
rect 308949 1002010 309015 1002013
rect 309777 1002010 309843 1002013
rect 310145 1002010 310211 1002013
rect 306097 1002008 306360 1002010
rect 306097 1001952 306102 1002008
rect 306158 1001952 306360 1002008
rect 306097 1001950 306360 1001952
rect 308949 1002008 309212 1002010
rect 308949 1001952 308954 1002008
rect 309010 1001952 309212 1002008
rect 308949 1001950 309212 1001952
rect 309580 1002008 309843 1002010
rect 309580 1001952 309782 1002008
rect 309838 1001952 309843 1002008
rect 309580 1001950 309843 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 306097 1001947 306163 1001950
rect 308949 1001947 309015 1001950
rect 309777 1001947 309843 1001950
rect 310145 1001947 310211 1001950
rect 354029 1002010 354095 1002013
rect 356881 1002010 356947 1002013
rect 358537 1002010 358603 1002013
rect 360193 1002010 360259 1002013
rect 365897 1002010 365963 1002013
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 356881 1002008 357144 1002010
rect 356881 1001952 356886 1002008
rect 356942 1001952 357144 1002008
rect 356881 1001950 357144 1001952
rect 358537 1002008 358800 1002010
rect 358537 1001952 358542 1002008
rect 358598 1001952 358800 1002008
rect 358537 1001950 358800 1001952
rect 359996 1002008 360259 1002010
rect 359996 1001952 360198 1002008
rect 360254 1001952 360259 1002008
rect 359996 1001950 360259 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 354029 1001947 354095 1001950
rect 356881 1001947 356947 1001950
rect 358537 1001947 358603 1001950
rect 360193 1001947 360259 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 424317 1002010 424383 1002013
rect 427537 1002010 427603 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 424317 1002008 424580 1002010
rect 424317 1001952 424322 1002008
rect 424378 1001952 424580 1002008
rect 424317 1001950 424580 1001952
rect 427340 1002008 427603 1002010
rect 427340 1001952 427542 1002008
rect 427598 1001952 427603 1002008
rect 427340 1001950 427603 1001952
rect 421465 1001947 421531 1001950
rect 424317 1001947 424383 1001950
rect 427537 1001947 427603 1001950
rect 501689 1002010 501755 1002013
rect 502517 1002010 502583 1002013
rect 504173 1002010 504239 1002013
rect 501689 1002008 501952 1002010
rect 501689 1001952 501694 1002008
rect 501750 1001952 501952 1002008
rect 501689 1001950 501952 1001952
rect 502412 1002008 502583 1002010
rect 502412 1001952 502522 1002008
rect 502578 1001952 502583 1002008
rect 502412 1001950 502583 1001952
rect 503976 1002008 504239 1002010
rect 503976 1001952 504178 1002008
rect 504234 1001952 504239 1002008
rect 503976 1001950 504239 1001952
rect 501689 1001947 501755 1001950
rect 502517 1001947 502583 1001950
rect 504173 1001947 504239 1001950
rect 505369 1002010 505435 1002013
rect 510337 1002010 510403 1002013
rect 505369 1002008 505632 1002010
rect 505369 1001952 505374 1002008
rect 505430 1001952 505632 1002008
rect 505369 1001950 505632 1001952
rect 510140 1002008 510403 1002010
rect 510140 1001952 510342 1002008
rect 510398 1001952 510403 1002008
rect 510140 1001950 510403 1001952
rect 505369 1001947 505435 1001950
rect 510337 1001947 510403 1001950
rect 554313 1002010 554379 1002013
rect 561673 1002010 561739 1002013
rect 554313 1002008 554576 1002010
rect 554313 1001952 554318 1002008
rect 554374 1001952 554576 1002008
rect 554313 1001950 554576 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 554313 1001947 554379 1001950
rect 561673 1001947 561739 1001950
rect 203885 1001194 203951 1001197
rect 550265 1001194 550331 1001197
rect 203885 1001192 204148 1001194
rect 203885 1001136 203890 1001192
rect 203946 1001136 204148 1001192
rect 203885 1001134 204148 1001136
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 203885 1001131 203951 1001134
rect 550265 1001131 550331 1001134
rect 555141 999154 555207 999157
rect 555036 999152 555207 999154
rect 555036 999096 555146 999152
rect 555202 999096 555207 999152
rect 555036 999094 555207 999096
rect 555141 999091 555207 999094
rect 298093 998882 298159 998885
rect 300485 998882 300551 998885
rect 298093 998880 300551 998882
rect 298093 998824 298098 998880
rect 298154 998824 300490 998880
rect 300546 998824 300551 998880
rect 298093 998822 300551 998824
rect 298093 998819 298159 998822
rect 300485 998819 300551 998822
rect 428365 998882 428431 998885
rect 428365 998880 428628 998882
rect 428365 998824 428370 998880
rect 428426 998824 428628 998880
rect 428365 998822 428628 998824
rect 428365 998819 428431 998822
rect 204345 998746 204411 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 204345 998683 204411 998686
rect 203517 998610 203583 998613
rect 430849 998610 430915 998613
rect 203320 998608 203583 998610
rect 203320 998552 203522 998608
rect 203578 998552 203583 998608
rect 203320 998550 203583 998552
rect 430652 998608 430915 998610
rect 430652 998552 430854 998608
rect 430910 998552 430915 998608
rect 430652 998550 430915 998552
rect 203517 998547 203583 998550
rect 430849 998547 430915 998550
rect 516869 998610 516935 998613
rect 516869 998608 524154 998610
rect 516869 998552 516874 998608
rect 516930 998552 524154 998608
rect 516869 998550 524154 998552
rect 516869 998547 516935 998550
rect 203517 998338 203583 998341
rect 376017 998338 376083 998341
rect 430021 998338 430087 998341
rect 203517 998336 203780 998338
rect 203517 998280 203522 998336
rect 203578 998280 203780 998336
rect 203517 998278 203780 998280
rect 376017 998336 383762 998338
rect 376017 998280 376022 998336
rect 376078 998280 383762 998336
rect 376017 998278 383762 998280
rect 429824 998336 430087 998338
rect 429824 998280 430026 998336
rect 430082 998280 430087 998336
rect 429824 998278 430087 998280
rect 203517 998275 203583 998278
rect 376017 998275 376083 998278
rect 202689 998202 202755 998205
rect 253657 998202 253723 998205
rect 202689 998200 202952 998202
rect 202689 998144 202694 998200
rect 202750 998144 202952 998200
rect 202689 998142 202952 998144
rect 253657 998200 253920 998202
rect 253657 998144 253662 998200
rect 253718 998144 253920 998200
rect 253657 998142 253920 998144
rect 202689 998139 202755 998142
rect 253657 998139 253723 998142
rect 201861 998066 201927 998069
rect 205541 998066 205607 998069
rect 201861 998064 202124 998066
rect 201861 998008 201866 998064
rect 201922 998008 202124 998064
rect 201861 998006 202124 998008
rect 205344 998064 205607 998066
rect 205344 998008 205546 998064
rect 205602 998008 205607 998064
rect 205344 998006 205607 998008
rect 201861 998003 201927 998006
rect 205541 998003 205607 998006
rect 200665 997930 200731 997933
rect 204713 997930 204779 997933
rect 253657 997930 253723 997933
rect 200665 997928 200836 997930
rect 200665 997872 200670 997928
rect 200726 997872 200836 997928
rect 200665 997870 200836 997872
rect 204713 997928 204976 997930
rect 204713 997872 204718 997928
rect 204774 997872 204976 997928
rect 204713 997870 204976 997872
rect 253460 997928 253723 997930
rect 253460 997872 253662 997928
rect 253718 997872 253723 997928
rect 253460 997870 253723 997872
rect 200665 997867 200731 997870
rect 204713 997867 204779 997870
rect 253657 997867 253723 997870
rect 198733 997794 198799 997797
rect 200021 997794 200087 997797
rect 252461 997794 252527 997797
rect 198733 997792 200087 997794
rect 198733 997736 198738 997792
rect 198794 997736 200026 997792
rect 200082 997736 200087 997792
rect 198733 997734 200087 997736
rect 252264 997792 252527 997794
rect 252264 997736 252466 997792
rect 252522 997736 252527 997792
rect 252264 997734 252527 997736
rect 198733 997731 198799 997734
rect 200021 997731 200087 997734
rect 252461 997731 252527 997734
rect 298645 997794 298711 997797
rect 301681 997794 301747 997797
rect 298645 997792 301747 997794
rect 298645 997736 298650 997792
rect 298706 997736 301686 997792
rect 301742 997736 301747 997792
rect 298645 997734 301747 997736
rect 298645 997731 298711 997734
rect 301681 997731 301747 997734
rect 89478 997188 89484 997252
rect 89548 997250 89554 997252
rect 92565 997250 92631 997253
rect 97441 997250 97507 997253
rect 89548 997248 92631 997250
rect 89548 997192 92570 997248
rect 92626 997192 92631 997248
rect 89548 997190 92631 997192
rect 89548 997188 89554 997190
rect 92565 997187 92631 997190
rect 93810 997248 97507 997250
rect 93810 997192 97446 997248
rect 97502 997192 97507 997248
rect 93810 997190 97507 997192
rect 92933 996978 92999 996981
rect 85254 996976 92999 996978
rect 85254 996920 92938 996976
rect 92994 996920 92999 996976
rect 85254 996918 92999 996920
rect 85254 996706 85314 996918
rect 92933 996915 92999 996918
rect 93810 996706 93870 997190
rect 97441 997187 97507 997190
rect 117129 997250 117195 997253
rect 143809 997250 143875 997253
rect 117129 997248 143875 997250
rect 117129 997192 117134 997248
rect 117190 997192 143814 997248
rect 143870 997192 143875 997248
rect 117129 997190 143875 997192
rect 117129 997187 117195 997190
rect 143809 997187 143875 997190
rect 195278 997188 195284 997252
rect 195348 997250 195354 997252
rect 195348 997190 195990 997250
rect 195348 997188 195354 997190
rect 189758 997052 189764 997116
rect 189828 997114 189834 997116
rect 195145 997114 195211 997117
rect 189828 997112 195211 997114
rect 189828 997056 195150 997112
rect 195206 997056 195211 997112
rect 189828 997054 195211 997056
rect 195930 997114 195990 997190
rect 243486 997188 243492 997252
rect 243556 997250 243562 997252
rect 247493 997250 247559 997253
rect 249057 997250 249123 997253
rect 243556 997248 247559 997250
rect 243556 997192 247498 997248
rect 247554 997192 247559 997248
rect 243556 997190 247559 997192
rect 243556 997188 243562 997190
rect 247493 997187 247559 997190
rect 248370 997248 249123 997250
rect 248370 997192 249062 997248
rect 249118 997192 249123 997248
rect 248370 997190 249123 997192
rect 198733 997114 198799 997117
rect 195930 997112 198799 997114
rect 195930 997056 198738 997112
rect 198794 997056 198799 997112
rect 195930 997054 198799 997056
rect 189828 997052 189834 997054
rect 195145 997051 195211 997054
rect 198733 997051 198799 997054
rect 116117 996978 116183 996981
rect 144821 996978 144887 996981
rect 116117 996976 144887 996978
rect 116117 996920 116122 996976
rect 116178 996920 144826 996976
rect 144882 996920 144887 996976
rect 116117 996918 144887 996920
rect 116117 996915 116183 996918
rect 144821 996915 144887 996918
rect 243854 996916 243860 996980
rect 243924 996978 243930 996980
rect 246941 996978 247007 996981
rect 243924 996976 247007 996978
rect 243924 996920 246946 996976
rect 247002 996920 247007 996976
rect 243924 996918 247007 996920
rect 243924 996916 243930 996918
rect 246941 996915 247007 996918
rect 195053 996842 195119 996845
rect 200205 996842 200271 996845
rect 195053 996840 200271 996842
rect 195053 996784 195058 996840
rect 195114 996784 200210 996840
rect 200266 996784 200271 996840
rect 195053 996782 200271 996784
rect 195053 996779 195119 996782
rect 200205 996779 200271 996782
rect 144637 996706 144703 996709
rect 194910 996706 194916 996708
rect 85070 996646 85314 996706
rect 89670 996646 93870 996706
rect 140270 996704 144703 996706
rect 140270 996648 144642 996704
rect 144698 996648 144703 996704
rect 140270 996646 144703 996648
rect 85070 995890 85130 996646
rect 89670 996434 89730 996646
rect 84886 995830 85130 995890
rect 85254 996374 89730 996434
rect 84653 995754 84719 995757
rect 84886 995754 84946 995830
rect 85254 995757 85314 996374
rect 89846 996236 89852 996300
rect 89916 996298 89922 996300
rect 92749 996298 92815 996301
rect 89916 996296 92815 996298
rect 89916 996240 92754 996296
rect 92810 996240 92815 996296
rect 89916 996238 92815 996240
rect 89916 996236 89922 996238
rect 92749 996235 92815 996238
rect 126237 996298 126303 996301
rect 140078 996298 140084 996300
rect 126237 996296 140084 996298
rect 126237 996240 126242 996296
rect 126298 996240 140084 996296
rect 126237 996238 140084 996240
rect 126237 996235 126303 996238
rect 140078 996236 140084 996238
rect 140148 996236 140154 996300
rect 89670 995966 93870 996026
rect 89670 995890 89730 995966
rect 87646 995830 89730 995890
rect 93810 995890 93870 995966
rect 98821 995890 98887 995893
rect 93810 995888 98887 995890
rect 93810 995832 98826 995888
rect 98882 995832 98887 995888
rect 93810 995830 98887 995832
rect 84653 995752 84946 995754
rect 84653 995696 84658 995752
rect 84714 995696 84946 995752
rect 84653 995694 84946 995696
rect 85205 995752 85314 995757
rect 85205 995696 85210 995752
rect 85266 995696 85314 995752
rect 85205 995694 85314 995696
rect 86033 995754 86099 995757
rect 87646 995754 87706 995830
rect 98821 995827 98887 995830
rect 86033 995752 87706 995754
rect 86033 995696 86038 995752
rect 86094 995696 87706 995752
rect 86033 995694 87706 995696
rect 90265 995754 90331 995757
rect 93485 995754 93551 995757
rect 90265 995752 93551 995754
rect 90265 995696 90270 995752
rect 90326 995696 93490 995752
rect 93546 995696 93551 995752
rect 90265 995694 93551 995696
rect 84653 995691 84719 995694
rect 85205 995691 85271 995694
rect 86033 995691 86099 995694
rect 90265 995691 90331 995694
rect 93485 995691 93551 995694
rect 88977 995618 89043 995621
rect 89529 995620 89595 995621
rect 89294 995618 89300 995620
rect 88977 995616 89300 995618
rect 88977 995560 88982 995616
rect 89038 995560 89300 995616
rect 88977 995558 89300 995560
rect 88977 995555 89043 995558
rect 89294 995556 89300 995558
rect 89364 995556 89370 995620
rect 89478 995556 89484 995620
rect 89548 995618 89595 995620
rect 89548 995616 89640 995618
rect 89590 995560 89640 995616
rect 89548 995558 89640 995560
rect 89548 995556 89595 995558
rect 89529 995555 89595 995556
rect 77201 995346 77267 995349
rect 101397 995346 101463 995349
rect 77201 995344 101463 995346
rect 77201 995288 77206 995344
rect 77262 995288 101402 995344
rect 101458 995288 101463 995344
rect 77201 995286 101463 995288
rect 77201 995283 77267 995286
rect 101397 995283 101463 995286
rect 80145 995074 80211 995077
rect 103746 995074 103806 996132
rect 132350 995964 132356 996028
rect 132420 996026 132426 996028
rect 132420 995966 132970 996026
rect 132420 995964 132426 995966
rect 132910 995757 132970 995966
rect 140270 995890 140330 996646
rect 144637 996643 144703 996646
rect 191974 996646 194916 996706
rect 136958 995830 140330 995890
rect 140454 996374 144562 996434
rect 131849 995754 131915 995757
rect 132534 995754 132540 995756
rect 131849 995752 132540 995754
rect 131849 995696 131854 995752
rect 131910 995696 132540 995752
rect 131849 995694 132540 995696
rect 131849 995691 131915 995694
rect 132534 995692 132540 995694
rect 132604 995692 132610 995756
rect 132910 995752 133019 995757
rect 132910 995696 132958 995752
rect 133014 995696 133019 995752
rect 132910 995694 133019 995696
rect 132953 995691 133019 995694
rect 136725 995754 136791 995757
rect 136958 995754 137018 995830
rect 140454 995757 140514 996374
rect 144502 996301 144562 996374
rect 188102 996372 188108 996436
rect 188172 996434 188178 996436
rect 191974 996434 192034 996646
rect 194910 996644 194916 996646
rect 194980 996644 194986 996708
rect 248045 996706 248111 996709
rect 234478 996704 248111 996706
rect 234478 996648 248050 996704
rect 248106 996648 248111 996704
rect 234478 996646 248111 996648
rect 188172 996374 192034 996434
rect 188172 996372 188178 996374
rect 192334 996372 192340 996436
rect 192404 996434 192410 996436
rect 198181 996434 198247 996437
rect 192404 996432 198247 996434
rect 192404 996376 198186 996432
rect 198242 996376 198247 996432
rect 192404 996374 198247 996376
rect 192404 996372 192410 996374
rect 198181 996371 198247 996374
rect 144502 996296 144611 996301
rect 144502 996240 144550 996296
rect 144606 996240 144611 996296
rect 144502 996238 144611 996240
rect 144545 996235 144611 996238
rect 195697 996162 195763 996165
rect 192342 996160 195763 996162
rect 144269 995890 144335 995893
rect 136725 995752 137018 995754
rect 136725 995696 136730 995752
rect 136786 995696 137018 995752
rect 136725 995694 137018 995696
rect 140405 995752 140514 995757
rect 140405 995696 140410 995752
rect 140466 995696 140514 995752
rect 140405 995694 140514 995696
rect 140638 995888 144335 995890
rect 140638 995832 144274 995888
rect 144330 995832 144335 995888
rect 140638 995830 144335 995832
rect 136725 995691 136791 995694
rect 140405 995691 140471 995694
rect 137369 995482 137435 995485
rect 140638 995482 140698 995830
rect 144269 995827 144335 995830
rect 154297 995754 154363 995757
rect 156830 995754 156890 996132
rect 154297 995752 156890 995754
rect 154297 995696 154302 995752
rect 154358 995696 156890 995752
rect 154297 995694 156890 995696
rect 154297 995691 154363 995694
rect 141785 995618 141851 995621
rect 147121 995618 147187 995621
rect 141785 995616 147187 995618
rect 141785 995560 141790 995616
rect 141846 995560 147126 995616
rect 147182 995560 147187 995616
rect 141785 995558 147187 995560
rect 141785 995555 141851 995558
rect 147121 995555 147187 995558
rect 159222 995482 159282 996132
rect 192342 996104 195702 996160
rect 195758 996104 195763 996160
rect 192342 996102 195763 996104
rect 175917 996026 175983 996029
rect 191598 996026 191604 996028
rect 175917 996024 191604 996026
rect 175917 995968 175922 996024
rect 175978 995968 191604 996024
rect 175917 995966 191604 995968
rect 175917 995963 175983 995966
rect 191598 995964 191604 995966
rect 191668 995964 191674 996028
rect 192342 995890 192402 996102
rect 195697 996099 195763 996102
rect 202965 995890 203031 995893
rect 191790 995830 192402 995890
rect 193998 995888 203031 995890
rect 193998 995832 202970 995888
rect 203026 995832 203031 995888
rect 193998 995830 203031 995832
rect 191790 995757 191850 995830
rect 188061 995756 188127 995757
rect 188061 995754 188108 995756
rect 188016 995752 188108 995754
rect 188016 995696 188066 995752
rect 188016 995694 188108 995696
rect 188061 995692 188108 995694
rect 188172 995692 188178 995756
rect 189441 995754 189507 995757
rect 189758 995754 189764 995756
rect 189441 995752 189764 995754
rect 189441 995696 189446 995752
rect 189502 995696 189764 995752
rect 189441 995694 189764 995696
rect 188061 995691 188127 995692
rect 189441 995691 189507 995694
rect 189758 995692 189764 995694
rect 189828 995692 189834 995756
rect 191741 995752 191850 995757
rect 191741 995696 191746 995752
rect 191802 995696 191850 995752
rect 191741 995694 191850 995696
rect 192477 995754 192543 995757
rect 193998 995754 194058 995830
rect 202965 995827 203031 995830
rect 203149 995890 203215 995893
rect 208166 995890 208226 996132
rect 203149 995888 208226 995890
rect 203149 995832 203154 995888
rect 203210 995832 208226 995888
rect 203149 995830 208226 995832
rect 208393 995890 208459 995893
rect 209822 995890 209882 996132
rect 208393 995888 209882 995890
rect 208393 995832 208398 995888
rect 208454 995832 209882 995888
rect 208393 995830 209882 995832
rect 203149 995827 203215 995830
rect 208393 995827 208459 995830
rect 192477 995752 194058 995754
rect 192477 995696 192482 995752
rect 192538 995696 194058 995752
rect 192477 995694 194058 995696
rect 191741 995691 191807 995694
rect 192477 995691 192543 995694
rect 192293 995620 192359 995621
rect 192293 995618 192340 995620
rect 192248 995616 192340 995618
rect 192248 995560 192298 995616
rect 192248 995558 192340 995560
rect 192293 995556 192340 995558
rect 192404 995556 192410 995620
rect 194317 995618 194383 995621
rect 195053 995618 195119 995621
rect 210650 995618 210710 996132
rect 234478 995757 234538 996646
rect 248045 996643 248111 996646
rect 248370 996434 248430 997190
rect 249057 997187 249123 997190
rect 287830 997188 287836 997252
rect 287900 997250 287906 997252
rect 302877 997250 302943 997253
rect 287900 997248 302943 997250
rect 287900 997192 302882 997248
rect 302938 997192 302943 997248
rect 287900 997190 302943 997192
rect 383702 997250 383762 998278
rect 430021 998275 430087 998278
rect 431217 998202 431283 998205
rect 431020 998200 431283 998202
rect 431020 998144 431222 998200
rect 431278 998144 431283 998200
rect 431020 998142 431283 998144
rect 431217 998139 431283 998142
rect 432045 998066 432111 998069
rect 432045 998064 432308 998066
rect 432045 998008 432050 998064
rect 432106 998008 432308 998064
rect 432045 998006 432308 998008
rect 432045 998003 432111 998006
rect 417057 997799 417363 997893
rect 418245 997803 418551 997897
rect 430021 997794 430087 997797
rect 435357 997794 435423 997797
rect 524094 997796 524154 998550
rect 558821 998474 558887 998477
rect 558624 998472 558887 998474
rect 558624 998416 558826 998472
rect 558882 998416 558887 998472
rect 558624 998414 558887 998416
rect 558821 998411 558887 998414
rect 557993 998338 558059 998341
rect 557993 998336 558256 998338
rect 557993 998280 557998 998336
rect 558054 998280 558256 998336
rect 557993 998278 558256 998280
rect 557993 998275 558059 998278
rect 558821 998202 558887 998205
rect 558821 998200 559084 998202
rect 558821 998144 558826 998200
rect 558882 998144 559084 998200
rect 558821 998142 559084 998144
rect 558821 998139 558887 998142
rect 557993 998066 558059 998069
rect 557796 998064 558059 998066
rect 557796 998008 557998 998064
rect 558054 998008 558059 998064
rect 557796 998006 558059 998008
rect 557993 998003 558059 998006
rect 557625 997930 557691 997933
rect 560017 997930 560083 997933
rect 557428 997928 557691 997930
rect 557428 997872 557630 997928
rect 557686 997872 557691 997928
rect 557428 997870 557691 997872
rect 559820 997928 560083 997930
rect 559820 997872 560022 997928
rect 560078 997872 560083 997928
rect 559820 997870 560083 997872
rect 557625 997867 557691 997870
rect 560017 997867 560083 997870
rect 430021 997792 430284 997794
rect 430021 997736 430026 997792
rect 430082 997736 430284 997792
rect 430021 997734 430284 997736
rect 433136 997792 435423 997794
rect 433136 997736 435362 997792
rect 435418 997736 435423 997792
rect 433136 997734 435423 997736
rect 430021 997731 430087 997734
rect 435357 997731 435423 997734
rect 524086 997732 524092 997796
rect 524156 997732 524162 997796
rect 553945 997794 554011 997797
rect 553748 997792 554011 997794
rect 553748 997736 553950 997792
rect 554006 997736 554011 997792
rect 553748 997734 554011 997736
rect 553945 997731 554011 997734
rect 385902 997250 385908 997252
rect 383702 997190 385908 997250
rect 287900 997188 287906 997190
rect 302877 997187 302943 997190
rect 385902 997188 385908 997190
rect 385972 997188 385978 997252
rect 439681 997250 439747 997253
rect 488901 997250 488967 997253
rect 510981 997252 511047 997253
rect 510981 997250 511028 997252
rect 439681 997248 488967 997250
rect 439681 997192 439686 997248
rect 439742 997192 488906 997248
rect 488962 997192 488967 997248
rect 439681 997190 488967 997192
rect 510936 997248 511028 997250
rect 510936 997192 510986 997248
rect 510936 997190 511028 997192
rect 439681 997187 439747 997190
rect 488901 997187 488967 997190
rect 510981 997188 511028 997190
rect 511092 997188 511098 997252
rect 524045 997250 524111 997253
rect 532550 997250 532556 997252
rect 524045 997248 532556 997250
rect 524045 997192 524050 997248
rect 524106 997192 532556 997248
rect 524045 997190 532556 997192
rect 510981 997187 511047 997188
rect 524045 997187 524111 997190
rect 532550 997188 532556 997190
rect 532620 997188 532626 997252
rect 553526 997250 553532 997252
rect 553380 997190 553532 997250
rect 553526 997188 553532 997190
rect 553596 997188 553602 997252
rect 623681 997250 623747 997253
rect 630254 997250 630260 997252
rect 623681 997248 630260 997250
rect 623681 997192 623686 997248
rect 623742 997192 630260 997248
rect 623681 997190 630260 997192
rect 623681 997187 623747 997190
rect 630254 997188 630260 997190
rect 630324 997188 630330 997252
rect 295374 996916 295380 996980
rect 295444 996978 295450 996980
rect 299197 996978 299263 996981
rect 295444 996976 299263 996978
rect 295444 996920 299202 996976
rect 299258 996920 299263 996976
rect 295444 996918 299263 996920
rect 295444 996916 295450 996918
rect 299197 996915 299263 996918
rect 372521 996978 372587 996981
rect 399937 996978 400003 996981
rect 372521 996976 400003 996978
rect 372521 996920 372526 996976
rect 372582 996920 399942 996976
rect 399998 996920 400003 996976
rect 372521 996918 400003 996920
rect 372521 996915 372587 996918
rect 399937 996915 400003 996918
rect 439865 996978 439931 996981
rect 489085 996978 489151 996981
rect 439865 996976 489151 996978
rect 439865 996920 439870 996976
rect 439926 996920 489090 996976
rect 489146 996920 489151 996976
rect 439865 996918 489151 996920
rect 439865 996915 439931 996918
rect 489085 996915 489151 996918
rect 517053 996978 517119 996981
rect 540881 996978 540947 996981
rect 517053 996976 540947 996978
rect 517053 996920 517058 996976
rect 517114 996920 540886 996976
rect 540942 996920 540947 996976
rect 517053 996918 540947 996920
rect 517053 996915 517119 996918
rect 540881 996915 540947 996918
rect 590561 996978 590627 996981
rect 633934 996978 633940 996980
rect 590561 996976 633940 996978
rect 590561 996920 590566 996976
rect 590622 996920 633940 996976
rect 590561 996918 633940 996920
rect 590561 996915 590627 996918
rect 633934 996916 633940 996918
rect 634004 996916 634010 996980
rect 291510 996644 291516 996708
rect 291580 996706 291586 996708
rect 302233 996706 302299 996709
rect 291580 996704 302299 996706
rect 291580 996648 302238 996704
rect 302294 996648 302299 996704
rect 291580 996646 302299 996648
rect 291580 996644 291586 996646
rect 302233 996643 302299 996646
rect 372337 996706 372403 996709
rect 388662 996706 388668 996708
rect 372337 996704 388668 996706
rect 372337 996648 372342 996704
rect 372398 996648 388668 996704
rect 372337 996646 388668 996648
rect 372337 996643 372403 996646
rect 388662 996644 388668 996646
rect 388732 996644 388738 996708
rect 489729 996706 489795 996709
rect 489913 996706 489979 996709
rect 489729 996704 489979 996706
rect 489729 996648 489734 996704
rect 489790 996648 489918 996704
rect 489974 996648 489979 996704
rect 489729 996646 489979 996648
rect 489729 996643 489795 996646
rect 489913 996643 489979 996646
rect 523493 996706 523559 996709
rect 529790 996706 529796 996708
rect 523493 996704 529796 996706
rect 523493 996648 523498 996704
rect 523554 996648 529796 996704
rect 523493 996646 529796 996648
rect 523493 996643 523559 996646
rect 529790 996644 529796 996646
rect 529860 996644 529866 996708
rect 538254 996706 538260 996708
rect 536238 996646 538260 996706
rect 298461 996434 298527 996437
rect 238526 996374 248430 996434
rect 282686 996432 298527 996434
rect 282686 996376 298466 996432
rect 298522 996376 298527 996432
rect 282686 996374 298527 996376
rect 238526 995757 238586 996374
rect 247309 996026 247375 996029
rect 240550 996024 247375 996026
rect 240550 995968 247314 996024
rect 247370 995968 247375 996024
rect 240550 995966 247375 995968
rect 234478 995752 234587 995757
rect 234478 995696 234526 995752
rect 234582 995696 234587 995752
rect 234478 995694 234587 995696
rect 238526 995752 238635 995757
rect 238526 995696 238574 995752
rect 238630 995696 238635 995752
rect 238526 995694 238635 995696
rect 234521 995691 234587 995694
rect 238569 995691 238635 995694
rect 240041 995754 240107 995757
rect 240550 995754 240610 995966
rect 247309 995963 247375 995966
rect 282686 995757 282746 996374
rect 298461 996371 298527 996374
rect 396574 996372 396580 996436
rect 396644 996434 396650 996436
rect 414473 996434 414539 996437
rect 396644 996432 414539 996434
rect 396644 996376 414478 996432
rect 414534 996376 414539 996432
rect 396644 996374 414539 996376
rect 396644 996372 396650 996374
rect 414473 996371 414539 996374
rect 516685 996434 516751 996437
rect 524045 996434 524111 996437
rect 516685 996432 524111 996434
rect 516685 996376 516690 996432
rect 516746 996376 524050 996432
rect 524106 996376 524111 996432
rect 516685 996374 524111 996376
rect 516685 996371 516751 996374
rect 524045 996371 524111 996374
rect 381537 996298 381603 996301
rect 385350 996298 385356 996300
rect 381537 996296 385356 996298
rect 381537 996240 381542 996296
rect 381598 996240 385356 996296
rect 381537 996238 385356 996240
rect 381537 996235 381603 996238
rect 385350 996236 385356 996238
rect 385420 996236 385426 996300
rect 445017 996298 445083 996301
rect 471145 996298 471211 996301
rect 484342 996298 484348 996300
rect 445017 996296 471211 996298
rect 445017 996240 445022 996296
rect 445078 996240 471150 996296
rect 471206 996240 471211 996296
rect 445017 996238 471211 996240
rect 445017 996235 445083 996238
rect 471145 996235 471211 996238
rect 476070 996238 484348 996298
rect 292246 996162 292252 996164
rect 290782 996102 292252 996162
rect 240041 995752 240610 995754
rect 240041 995696 240046 995752
rect 240102 995696 240610 995752
rect 240041 995694 240610 995696
rect 243445 995756 243511 995757
rect 243813 995756 243879 995757
rect 243445 995752 243492 995756
rect 243556 995754 243562 995756
rect 243813 995754 243860 995756
rect 243445 995696 243450 995752
rect 240041 995691 240107 995694
rect 243445 995692 243492 995696
rect 243556 995694 243602 995754
rect 243768 995752 243860 995754
rect 243768 995696 243818 995752
rect 243768 995694 243860 995696
rect 243556 995692 243562 995694
rect 243813 995692 243860 995694
rect 243924 995692 243930 995756
rect 244089 995754 244155 995757
rect 246757 995754 246823 995757
rect 244089 995752 246823 995754
rect 244089 995696 244094 995752
rect 244150 995696 246762 995752
rect 246818 995696 246823 995752
rect 244089 995694 246823 995696
rect 282686 995752 282795 995757
rect 282686 995696 282734 995752
rect 282790 995696 282795 995752
rect 282686 995694 282795 995696
rect 243445 995691 243511 995692
rect 243813 995691 243879 995692
rect 244089 995691 244155 995694
rect 246757 995691 246823 995694
rect 282729 995691 282795 995694
rect 286777 995754 286843 995757
rect 290782 995754 290842 996102
rect 292246 996100 292252 996102
rect 292316 996100 292322 996164
rect 476070 996162 476130 996238
rect 484342 996236 484348 996238
rect 484412 996236 484418 996300
rect 298093 996026 298159 996029
rect 295014 996024 298159 996026
rect 295014 995968 298098 996024
rect 298154 995968 298159 996024
rect 295014 995966 298159 995968
rect 286777 995752 290842 995754
rect 286777 995696 286782 995752
rect 286838 995696 290842 995752
rect 286777 995694 290842 995696
rect 293585 995754 293651 995757
rect 295014 995754 295074 995966
rect 298093 995963 298159 995966
rect 295333 995756 295399 995757
rect 295333 995754 295380 995756
rect 293585 995752 295074 995754
rect 293585 995696 293590 995752
rect 293646 995696 295074 995752
rect 293585 995694 295074 995696
rect 295288 995752 295380 995754
rect 295288 995696 295338 995752
rect 295288 995694 295380 995696
rect 286777 995691 286843 995694
rect 293585 995691 293651 995694
rect 295333 995692 295380 995694
rect 295444 995692 295450 995756
rect 297265 995754 297331 995757
rect 298277 995754 298343 995757
rect 297265 995752 298343 995754
rect 297265 995696 297270 995752
rect 297326 995696 298282 995752
rect 298338 995696 298343 995752
rect 297265 995694 298343 995696
rect 295333 995691 295399 995692
rect 297265 995691 297331 995694
rect 298277 995691 298343 995694
rect 194317 995616 195119 995618
rect 194317 995560 194322 995616
rect 194378 995560 195058 995616
rect 195114 995560 195119 995616
rect 194317 995558 195119 995560
rect 192293 995555 192359 995556
rect 194317 995555 194383 995558
rect 195053 995555 195119 995558
rect 195286 995558 210710 995618
rect 240869 995618 240935 995621
rect 243261 995618 243327 995621
rect 240869 995616 243327 995618
rect 240869 995560 240874 995616
rect 240930 995560 243266 995616
rect 243322 995560 243327 995616
rect 240869 995558 243327 995560
rect 137369 995480 140698 995482
rect 137369 995424 137374 995480
rect 137430 995424 140698 995480
rect 137369 995422 140698 995424
rect 151770 995422 159282 995482
rect 137369 995419 137435 995422
rect 132401 995348 132467 995349
rect 132350 995346 132356 995348
rect 132310 995286 132356 995346
rect 132420 995344 132467 995348
rect 132462 995288 132467 995344
rect 132350 995284 132356 995286
rect 132420 995284 132467 995288
rect 140814 995284 140820 995348
rect 140884 995346 140890 995348
rect 151770 995346 151830 995422
rect 140884 995286 151830 995346
rect 177297 995346 177363 995349
rect 195286 995346 195346 995558
rect 240869 995555 240935 995558
rect 243261 995555 243327 995558
rect 292430 995556 292436 995620
rect 292500 995618 292506 995620
rect 293217 995618 293283 995621
rect 292500 995616 293283 995618
rect 292500 995560 293222 995616
rect 293278 995560 293283 995616
rect 292500 995558 293283 995560
rect 292500 995556 292506 995558
rect 293217 995555 293283 995558
rect 295517 995618 295583 995621
rect 296897 995618 296963 995621
rect 295517 995616 296963 995618
rect 295517 995560 295522 995616
rect 295578 995560 296902 995616
rect 296958 995560 296963 995616
rect 295517 995558 296963 995560
rect 295517 995555 295583 995558
rect 296897 995555 296963 995558
rect 298461 995618 298527 995621
rect 301497 995618 301563 995621
rect 298461 995616 301563 995618
rect 298461 995560 298466 995616
rect 298522 995560 301502 995616
rect 301558 995560 301563 995616
rect 298461 995558 301563 995560
rect 298461 995555 298527 995558
rect 301497 995555 301563 995558
rect 308765 995618 308831 995621
rect 311206 995618 311266 996132
rect 308765 995616 311266 995618
rect 308765 995560 308770 995616
rect 308826 995560 311266 995616
rect 308765 995558 311266 995560
rect 308765 995555 308831 995558
rect 177297 995344 195346 995346
rect 177297 995288 177302 995344
rect 177358 995288 195346 995344
rect 177297 995286 195346 995288
rect 195513 995346 195579 995349
rect 203149 995346 203215 995349
rect 241881 995346 241947 995349
rect 195513 995344 203215 995346
rect 195513 995288 195518 995344
rect 195574 995288 203154 995344
rect 203210 995288 203215 995344
rect 195513 995286 203215 995288
rect 140884 995284 140890 995286
rect 132401 995283 132467 995284
rect 177297 995283 177363 995286
rect 195513 995283 195579 995286
rect 203149 995283 203215 995286
rect 238710 995344 241947 995346
rect 238710 995288 241886 995344
rect 241942 995288 241947 995344
rect 238710 995286 241947 995288
rect 171041 995210 171107 995213
rect 171501 995210 171567 995213
rect 171041 995208 171567 995210
rect 171041 995152 171046 995208
rect 171102 995152 171506 995208
rect 171562 995152 171567 995208
rect 171041 995150 171567 995152
rect 171041 995147 171107 995150
rect 171501 995147 171567 995150
rect 80145 995072 103806 995074
rect 80145 995016 80150 995072
rect 80206 995016 103806 995072
rect 80145 995014 103806 995016
rect 124857 995074 124923 995077
rect 154297 995074 154363 995077
rect 124857 995072 154363 995074
rect 124857 995016 124862 995072
rect 124918 995016 154302 995072
rect 154358 995016 154363 995072
rect 124857 995014 154363 995016
rect 80145 995011 80211 995014
rect 124857 995011 124923 995014
rect 154297 995011 154363 995014
rect 173157 995074 173223 995077
rect 208393 995074 208459 995077
rect 173157 995072 208459 995074
rect 173157 995016 173162 995072
rect 173218 995016 208398 995072
rect 208454 995016 208459 995072
rect 173157 995014 208459 995016
rect 173157 995011 173223 995014
rect 208393 995011 208459 995014
rect 235901 995074 235967 995077
rect 238710 995074 238770 995286
rect 241881 995283 241947 995286
rect 242065 995346 242131 995349
rect 253381 995346 253447 995349
rect 242065 995344 253447 995346
rect 242065 995288 242070 995344
rect 242126 995288 253386 995344
rect 253442 995288 253447 995344
rect 242065 995286 253447 995288
rect 242065 995283 242131 995286
rect 253381 995283 253447 995286
rect 279417 995346 279483 995349
rect 312862 995346 312922 996132
rect 471286 996102 476130 996162
rect 373257 996026 373323 996029
rect 380893 996026 380959 996029
rect 466361 996026 466427 996029
rect 471286 996026 471346 996102
rect 373257 996024 379530 996026
rect 373257 995968 373262 996024
rect 373318 995968 379530 996024
rect 373257 995966 379530 995968
rect 373257 995963 373323 995966
rect 359457 995890 359523 995893
rect 364190 995890 364196 995892
rect 359457 995888 364196 995890
rect 359457 995832 359462 995888
rect 359518 995832 364196 995888
rect 359457 995830 364196 995832
rect 359457 995827 359523 995830
rect 364190 995828 364196 995830
rect 364260 995828 364266 995892
rect 279417 995344 312922 995346
rect 279417 995288 279422 995344
rect 279478 995288 312922 995344
rect 279417 995286 312922 995288
rect 279417 995283 279483 995286
rect 379470 995210 379530 995966
rect 380893 996024 393330 996026
rect 380893 995968 380898 996024
rect 380954 995968 393330 996024
rect 380893 995966 393330 995968
rect 380893 995963 380959 995966
rect 382273 995754 382339 995757
rect 388713 995756 388779 995757
rect 388478 995754 388484 995756
rect 382273 995752 388484 995754
rect 382273 995696 382278 995752
rect 382334 995696 388484 995752
rect 382273 995694 388484 995696
rect 382273 995691 382339 995694
rect 388478 995692 388484 995694
rect 388548 995692 388554 995756
rect 388662 995692 388668 995756
rect 388732 995754 388779 995756
rect 393270 995754 393330 995966
rect 466361 996024 471346 996026
rect 466361 995968 466366 996024
rect 466422 995968 471346 996024
rect 466361 995966 471346 995968
rect 479014 995966 489930 996026
rect 466361 995963 466427 995966
rect 471421 995890 471487 995893
rect 471421 995888 477970 995890
rect 471421 995832 471426 995888
rect 471482 995832 477970 995888
rect 471421 995830 477970 995832
rect 471421 995827 471487 995830
rect 416129 995754 416195 995757
rect 388732 995752 388824 995754
rect 388774 995696 388824 995752
rect 388732 995694 388824 995696
rect 393270 995752 416195 995754
rect 393270 995696 416134 995752
rect 416190 995696 416195 995752
rect 393270 995694 416195 995696
rect 477910 995754 477970 995830
rect 479014 995757 479074 995966
rect 478321 995754 478387 995757
rect 477910 995752 478387 995754
rect 477910 995696 478326 995752
rect 478382 995696 478387 995752
rect 477910 995694 478387 995696
rect 388732 995692 388779 995694
rect 388713 995691 388779 995692
rect 416129 995691 416195 995694
rect 478321 995691 478387 995694
rect 478965 995752 479074 995757
rect 478965 995696 478970 995752
rect 479026 995696 479074 995752
rect 478965 995694 479074 995696
rect 478965 995691 479031 995694
rect 484342 995692 484348 995756
rect 484412 995754 484418 995756
rect 485773 995754 485839 995757
rect 484412 995752 485839 995754
rect 484412 995696 485778 995752
rect 485834 995696 485839 995752
rect 484412 995694 485839 995696
rect 484412 995692 484418 995694
rect 485773 995691 485839 995694
rect 462957 995618 463023 995621
rect 477677 995618 477743 995621
rect 462957 995616 477743 995618
rect 462957 995560 462962 995616
rect 463018 995560 477682 995616
rect 477738 995560 477743 995616
rect 462957 995558 477743 995560
rect 462957 995555 463023 995558
rect 477677 995555 477743 995558
rect 383469 995482 383535 995485
rect 388161 995482 388227 995485
rect 392393 995482 392459 995485
rect 383469 995480 388227 995482
rect 383469 995424 383474 995480
rect 383530 995424 388166 995480
rect 388222 995424 388227 995480
rect 383469 995422 388227 995424
rect 383469 995419 383535 995422
rect 388161 995419 388227 995422
rect 389130 995480 392459 995482
rect 389130 995424 392398 995480
rect 392454 995424 392459 995480
rect 389130 995422 392459 995424
rect 389130 995346 389190 995422
rect 392393 995419 392459 995422
rect 393446 995420 393452 995484
rect 393516 995482 393522 995484
rect 393681 995482 393747 995485
rect 396533 995484 396599 995485
rect 396533 995482 396580 995484
rect 393516 995480 393747 995482
rect 393516 995424 393686 995480
rect 393742 995424 393747 995480
rect 393516 995422 393747 995424
rect 396488 995480 396580 995482
rect 396488 995424 396538 995480
rect 396488 995422 396580 995424
rect 393516 995420 393522 995422
rect 393681 995419 393747 995422
rect 396533 995420 396580 995422
rect 396644 995420 396650 995484
rect 415393 995482 415459 995485
rect 402930 995480 415459 995482
rect 402930 995424 415398 995480
rect 415454 995424 415459 995480
rect 402930 995422 415459 995424
rect 396533 995419 396599 995420
rect 388302 995286 389190 995346
rect 388302 995210 388362 995286
rect 379470 995150 388362 995210
rect 235901 995072 238770 995074
rect 235901 995016 235906 995072
rect 235962 995016 238770 995072
rect 235901 995014 238770 995016
rect 239581 995074 239647 995077
rect 246481 995074 246547 995077
rect 239581 995072 246547 995074
rect 239581 995016 239586 995072
rect 239642 995016 246486 995072
rect 246542 995016 246547 995072
rect 239581 995014 246547 995016
rect 235901 995011 235967 995014
rect 239581 995011 239647 995014
rect 246481 995011 246547 995014
rect 246665 995074 246731 995077
rect 250621 995074 250687 995077
rect 246665 995072 250687 995074
rect 246665 995016 246670 995072
rect 246726 995016 250626 995072
rect 250682 995016 250687 995072
rect 246665 995014 250687 995016
rect 246665 995011 246731 995014
rect 250621 995011 250687 995014
rect 270401 995074 270467 995077
rect 308765 995074 308831 995077
rect 270401 995072 308831 995074
rect 270401 995016 270406 995072
rect 270462 995016 308770 995072
rect 308826 995016 308831 995072
rect 385401 995042 385467 995043
rect 385350 995040 385356 995042
rect 270401 995014 308831 995016
rect 270401 995011 270467 995014
rect 308765 995011 308831 995014
rect 385310 994980 385356 995040
rect 385420 995038 385467 995042
rect 385462 994982 385467 995038
rect 388478 995012 388484 995076
rect 388548 995074 388554 995076
rect 402930 995074 402990 995422
rect 415393 995419 415459 995422
rect 485681 995482 485747 995485
rect 489269 995482 489335 995485
rect 485681 995480 489335 995482
rect 485681 995424 485686 995480
rect 485742 995424 489274 995480
rect 489330 995424 489335 995480
rect 485681 995422 489335 995424
rect 485681 995419 485747 995422
rect 489269 995419 489335 995422
rect 456793 995346 456859 995349
rect 480805 995346 480871 995349
rect 456793 995344 480871 995346
rect 456793 995288 456798 995344
rect 456854 995288 480810 995344
rect 480866 995288 480871 995344
rect 456793 995286 480871 995288
rect 489870 995346 489930 995966
rect 506430 995346 506490 996132
rect 489870 995286 506490 995346
rect 456793 995283 456859 995286
rect 480805 995283 480871 995286
rect 388548 995014 402990 995074
rect 469857 995074 469923 995077
rect 472249 995074 472315 995077
rect 469857 995072 472315 995074
rect 469857 995016 469862 995072
rect 469918 995016 472254 995072
rect 472310 995016 472315 995072
rect 469857 995014 472315 995016
rect 388548 995012 388554 995014
rect 469857 995011 469923 995014
rect 472249 995011 472315 995014
rect 472433 995074 472499 995077
rect 474733 995074 474799 995077
rect 472433 995072 474799 995074
rect 472433 995016 472438 995072
rect 472494 995016 474738 995072
rect 474794 995016 474799 995072
rect 472433 995014 474799 995016
rect 472433 995011 472499 995014
rect 474733 995011 474799 995014
rect 474917 995074 474983 995077
rect 476113 995074 476179 995077
rect 474917 995072 476179 995074
rect 474917 995016 474922 995072
rect 474978 995016 476118 995072
rect 476174 995016 476179 995072
rect 474917 995014 476179 995016
rect 474917 995011 474983 995014
rect 476113 995011 476179 995014
rect 476297 995074 476363 995077
rect 508822 995074 508882 996132
rect 520917 996026 520983 996029
rect 520917 996024 529306 996026
rect 520917 995968 520922 996024
rect 520978 995968 529306 996024
rect 520917 995966 529306 995968
rect 520917 995963 520983 995966
rect 516869 995754 516935 995757
rect 529013 995754 529079 995757
rect 516869 995752 529079 995754
rect 516869 995696 516874 995752
rect 516930 995696 529018 995752
rect 529074 995696 529079 995752
rect 516869 995694 529079 995696
rect 529246 995754 529306 995966
rect 529657 995754 529723 995757
rect 529246 995752 529723 995754
rect 529246 995696 529662 995752
rect 529718 995696 529723 995752
rect 529246 995694 529723 995696
rect 516869 995691 516935 995694
rect 529013 995691 529079 995694
rect 529657 995691 529723 995694
rect 531998 995692 532004 995756
rect 532068 995754 532074 995756
rect 532233 995754 532299 995757
rect 532068 995752 532299 995754
rect 532068 995696 532238 995752
rect 532294 995696 532299 995752
rect 532068 995694 532299 995696
rect 532068 995692 532074 995694
rect 532233 995691 532299 995694
rect 532550 995692 532556 995756
rect 532620 995754 532626 995756
rect 532785 995754 532851 995757
rect 532620 995752 532851 995754
rect 532620 995696 532790 995752
rect 532846 995696 532851 995752
rect 532620 995694 532851 995696
rect 532620 995692 532626 995694
rect 532785 995691 532851 995694
rect 534625 995754 534691 995757
rect 536238 995754 536298 996646
rect 538254 996644 538260 996646
rect 538324 996644 538330 996708
rect 590561 996706 590627 996709
rect 627862 996706 627868 996708
rect 590561 996704 627868 996706
rect 590561 996648 590566 996704
rect 590622 996648 627868 996704
rect 590561 996646 627868 996648
rect 590561 996643 590627 996646
rect 627862 996644 627868 996646
rect 627932 996644 627938 996708
rect 549437 996434 549503 996437
rect 536606 996432 549503 996434
rect 536606 996376 549442 996432
rect 549498 996376 549503 996432
rect 536606 996374 549503 996376
rect 536606 995757 536666 996374
rect 549437 996371 549503 996374
rect 590561 996434 590627 996437
rect 590561 996432 635290 996434
rect 590561 996376 590566 996432
rect 590622 996376 635290 996432
rect 590561 996374 635290 996376
rect 590561 996371 590627 996374
rect 534625 995752 536298 995754
rect 534625 995696 534630 995752
rect 534686 995696 536298 995752
rect 534625 995694 536298 995696
rect 536557 995752 536666 995757
rect 536557 995696 536562 995752
rect 536618 995696 536666 995752
rect 536557 995694 536666 995696
rect 534625 995691 534691 995694
rect 536557 995691 536623 995694
rect 529841 995620 529907 995621
rect 529790 995556 529796 995620
rect 529860 995618 529907 995620
rect 529860 995616 529952 995618
rect 529902 995560 529952 995616
rect 529860 995558 529952 995560
rect 529860 995556 529907 995558
rect 529841 995555 529907 995556
rect 517513 995346 517579 995349
rect 535637 995346 535703 995349
rect 517513 995344 535703 995346
rect 517513 995288 517518 995344
rect 517574 995288 535642 995344
rect 535698 995288 535703 995344
rect 517513 995286 535703 995288
rect 517513 995283 517579 995286
rect 535637 995283 535703 995286
rect 476297 995072 508882 995074
rect 476297 995016 476302 995072
rect 476358 995016 508882 995072
rect 476297 995014 508882 995016
rect 476297 995011 476363 995014
rect 522798 995012 522804 995076
rect 522868 995074 522874 995076
rect 527909 995074 527975 995077
rect 522868 995072 527975 995074
rect 522868 995016 527914 995072
rect 527970 995016 527975 995072
rect 522868 995014 527975 995016
rect 522868 995012 522874 995014
rect 527909 995011 527975 995014
rect 529657 995074 529723 995077
rect 559422 995074 559482 996132
rect 625429 996026 625495 996029
rect 625429 996024 629586 996026
rect 625429 995968 625434 996024
rect 625490 995968 629586 996024
rect 625429 995966 629586 995968
rect 625429 995963 625495 995966
rect 629526 995757 629586 995966
rect 635230 995757 635290 996374
rect 625613 995754 625679 995757
rect 627177 995754 627243 995757
rect 627913 995756 627979 995757
rect 625613 995752 627243 995754
rect 625613 995696 625618 995752
rect 625674 995696 627182 995752
rect 627238 995696 627243 995752
rect 625613 995694 627243 995696
rect 625613 995691 625679 995694
rect 627177 995691 627243 995694
rect 627862 995692 627868 995756
rect 627932 995754 627979 995756
rect 627932 995752 628024 995754
rect 627974 995696 628024 995752
rect 627932 995694 628024 995696
rect 629526 995752 629635 995757
rect 630305 995756 630371 995757
rect 633985 995756 634051 995757
rect 629526 995696 629574 995752
rect 629630 995696 629635 995752
rect 629526 995694 629635 995696
rect 627932 995692 627979 995694
rect 627913 995691 627979 995692
rect 629569 995691 629635 995694
rect 630254 995692 630260 995756
rect 630324 995754 630371 995756
rect 630324 995752 630416 995754
rect 630366 995696 630416 995752
rect 630324 995694 630416 995696
rect 630324 995692 630371 995694
rect 633934 995692 633940 995756
rect 634004 995754 634051 995756
rect 634004 995752 634096 995754
rect 634046 995696 634096 995752
rect 634004 995694 634096 995696
rect 635230 995752 635339 995757
rect 635230 995696 635278 995752
rect 635334 995696 635339 995752
rect 635230 995694 635339 995696
rect 634004 995692 634051 995694
rect 630305 995691 630371 995692
rect 633985 995691 634051 995692
rect 635273 995691 635339 995694
rect 636694 995692 636700 995756
rect 636764 995754 636770 995756
rect 637021 995754 637087 995757
rect 636764 995752 637087 995754
rect 636764 995696 637026 995752
rect 637082 995696 637087 995752
rect 636764 995694 637087 995696
rect 636764 995692 636770 995694
rect 637021 995691 637087 995694
rect 590745 995346 590811 995349
rect 634721 995346 634787 995349
rect 590745 995344 634787 995346
rect 590745 995288 590750 995344
rect 590806 995288 634726 995344
rect 634782 995288 634787 995344
rect 590745 995286 634787 995288
rect 590745 995283 590811 995286
rect 634721 995283 634787 995286
rect 529657 995072 559482 995074
rect 529657 995016 529662 995072
rect 529718 995016 559482 995072
rect 529657 995014 559482 995016
rect 590561 995074 590627 995077
rect 640977 995074 641043 995077
rect 590561 995072 641043 995074
rect 590561 995016 590566 995072
rect 590622 995016 640982 995072
rect 641038 995016 641043 995072
rect 590561 995014 641043 995016
rect 529657 995011 529723 995014
rect 590561 995011 590627 995014
rect 640977 995011 641043 995014
rect 385350 994978 385356 994980
rect 385420 994978 385467 994982
rect 385401 994977 385467 994978
rect 385953 994940 386019 994941
rect 385902 994876 385908 994940
rect 385972 994938 386019 994940
rect 385972 994936 386064 994938
rect 386014 994880 386064 994936
rect 385972 994878 386064 994880
rect 385972 994876 386019 994878
rect 385953 994875 386019 994876
rect 81985 994802 82051 994805
rect 93117 994802 93183 994805
rect 81985 994800 93183 994802
rect 81985 994744 81990 994800
rect 82046 994744 93122 994800
rect 93178 994744 93183 994800
rect 81985 994742 93183 994744
rect 81985 994739 82051 994742
rect 93117 994739 93183 994742
rect 132125 994802 132191 994805
rect 145557 994802 145623 994805
rect 132125 994800 145623 994802
rect 132125 994744 132130 994800
rect 132186 994744 145562 994800
rect 145618 994744 145623 994800
rect 132125 994742 145623 994744
rect 132125 994739 132191 994742
rect 145557 994739 145623 994742
rect 184841 994802 184907 994805
rect 184841 994800 188538 994802
rect 184841 994744 184846 994800
rect 184902 994744 188538 994800
rect 184841 994742 188538 994744
rect 184841 994739 184907 994742
rect 86309 994530 86375 994533
rect 97257 994530 97323 994533
rect 86309 994528 97323 994530
rect 86309 994472 86314 994528
rect 86370 994472 97262 994528
rect 97318 994472 97323 994528
rect 86309 994470 97323 994472
rect 86309 994467 86375 994470
rect 97257 994467 97323 994470
rect 142153 994530 142219 994533
rect 154573 994530 154639 994533
rect 142153 994528 154639 994530
rect 142153 994472 142158 994528
rect 142214 994472 154578 994528
rect 154634 994472 154639 994528
rect 142153 994470 154639 994472
rect 142153 994467 142219 994470
rect 154573 994467 154639 994470
rect 135897 994394 135963 994397
rect 141969 994394 142035 994397
rect 135897 994392 142035 994394
rect 135897 994336 135902 994392
rect 135958 994336 141974 994392
rect 142030 994336 142035 994392
rect 135897 994334 142035 994336
rect 135897 994331 135963 994334
rect 141969 994331 142035 994334
rect 186129 994394 186195 994397
rect 186497 994394 186563 994397
rect 186129 994392 186563 994394
rect 186129 994336 186134 994392
rect 186190 994336 186502 994392
rect 186558 994336 186563 994392
rect 186129 994334 186563 994336
rect 186129 994331 186195 994334
rect 186497 994331 186563 994334
rect 87873 994258 87939 994261
rect 95141 994258 95207 994261
rect 87873 994256 95207 994258
rect 87873 994200 87878 994256
rect 87934 994200 95146 994256
rect 95202 994200 95207 994256
rect 87873 994198 95207 994200
rect 87873 994195 87939 994198
rect 95141 994195 95207 994198
rect 142153 994258 142219 994261
rect 148501 994258 148567 994261
rect 142153 994256 148567 994258
rect 142153 994200 142158 994256
rect 142214 994200 148506 994256
rect 148562 994200 148567 994256
rect 142153 994198 148567 994200
rect 188478 994258 188538 994742
rect 191598 994740 191604 994804
rect 191668 994802 191674 994804
rect 195513 994802 195579 994805
rect 191668 994800 195579 994802
rect 191668 994744 195518 994800
rect 195574 994744 195579 994800
rect 191668 994742 195579 994744
rect 191668 994740 191674 994742
rect 195513 994739 195579 994742
rect 235257 994802 235323 994805
rect 253105 994802 253171 994805
rect 287789 994804 287855 994805
rect 291469 994804 291535 994805
rect 287789 994802 287836 994804
rect 235257 994800 253171 994802
rect 235257 994744 235262 994800
rect 235318 994744 253110 994800
rect 253166 994744 253171 994800
rect 235257 994742 253171 994744
rect 287744 994800 287836 994802
rect 287744 994744 287794 994800
rect 287744 994742 287836 994744
rect 235257 994739 235323 994742
rect 253105 994739 253171 994742
rect 287789 994740 287836 994742
rect 287900 994740 287906 994804
rect 291469 994802 291516 994804
rect 291424 994800 291516 994802
rect 291424 994744 291474 994800
rect 291424 994742 291516 994744
rect 291469 994740 291516 994742
rect 291580 994740 291586 994804
rect 309133 994802 309199 994805
rect 291702 994800 309199 994802
rect 291702 994744 309138 994800
rect 309194 994744 309199 994800
rect 291702 994742 309199 994744
rect 287789 994739 287855 994740
rect 291469 994739 291535 994740
rect 188797 994530 188863 994533
rect 200757 994530 200823 994533
rect 188797 994528 200823 994530
rect 188797 994472 188802 994528
rect 188858 994472 200762 994528
rect 200818 994472 200823 994528
rect 188797 994470 200823 994472
rect 188797 994467 188863 994470
rect 200757 994467 200823 994470
rect 241881 994530 241947 994533
rect 247861 994530 247927 994533
rect 241881 994528 247927 994530
rect 241881 994472 241886 994528
rect 241942 994472 247866 994528
rect 247922 994472 247927 994528
rect 241881 994470 247927 994472
rect 241881 994467 241947 994470
rect 247861 994467 247927 994470
rect 285949 994530 286015 994533
rect 291702 994530 291762 994742
rect 309133 994739 309199 994742
rect 464337 994802 464403 994805
rect 486601 994802 486667 994805
rect 464337 994800 486667 994802
rect 464337 994744 464342 994800
rect 464398 994744 486606 994800
rect 486662 994744 486667 994800
rect 464337 994742 486667 994744
rect 464337 994739 464403 994742
rect 486601 994739 486667 994742
rect 570413 994802 570479 994805
rect 630857 994802 630923 994805
rect 570413 994800 630923 994802
rect 570413 994744 570418 994800
rect 570474 994744 630862 994800
rect 630918 994744 630923 994800
rect 570413 994742 630923 994744
rect 570413 994739 570479 994742
rect 630857 994739 630923 994742
rect 304257 994530 304323 994533
rect 285949 994528 291762 994530
rect 285949 994472 285954 994528
rect 286010 994472 291762 994528
rect 285949 994470 291762 994472
rect 291886 994528 304323 994530
rect 291886 994472 304262 994528
rect 304318 994472 304323 994528
rect 291886 994470 304323 994472
rect 285949 994467 286015 994470
rect 196617 994258 196683 994261
rect 188478 994256 196683 994258
rect 188478 994200 196622 994256
rect 196678 994200 196683 994256
rect 188478 994198 196683 994200
rect 142153 994195 142219 994198
rect 148501 994195 148567 994198
rect 196617 994195 196683 994198
rect 287145 994258 287211 994261
rect 291886 994258 291946 994470
rect 304257 994467 304323 994470
rect 447777 994530 447843 994533
rect 482921 994530 482987 994533
rect 447777 994528 482987 994530
rect 447777 994472 447782 994528
rect 447838 994472 482926 994528
rect 482982 994472 482987 994528
rect 447777 994470 482987 994472
rect 447777 994467 447843 994470
rect 482921 994467 482987 994470
rect 538254 994468 538260 994532
rect 538324 994530 538330 994532
rect 538581 994530 538647 994533
rect 538324 994528 538647 994530
rect 538324 994472 538586 994528
rect 538642 994472 538647 994528
rect 538324 994470 538647 994472
rect 538324 994468 538330 994470
rect 538581 994467 538647 994470
rect 287145 994256 291946 994258
rect 287145 994200 287150 994256
rect 287206 994200 291946 994256
rect 287145 994198 291946 994200
rect 292113 994258 292179 994261
rect 300301 994258 300367 994261
rect 292113 994256 300367 994258
rect 292113 994200 292118 994256
rect 292174 994200 300306 994256
rect 300362 994200 300367 994256
rect 292113 994198 300367 994200
rect 287145 994195 287211 994198
rect 292113 994195 292179 994198
rect 300301 994195 300367 994198
rect 445661 994258 445727 994261
rect 481909 994258 481975 994261
rect 445661 994256 481975 994258
rect 445661 994200 445666 994256
rect 445722 994200 481914 994256
rect 481970 994200 481975 994256
rect 445661 994198 481975 994200
rect 445661 994195 445727 994198
rect 481909 994195 481975 994198
rect 133137 994122 133203 994125
rect 139209 994122 139275 994125
rect 133137 994120 139275 994122
rect 133137 994064 133142 994120
rect 133198 994064 139214 994120
rect 139270 994064 139275 994120
rect 133137 994062 139275 994064
rect 133137 994059 133203 994062
rect 139209 994059 139275 994062
rect 81065 993986 81131 993989
rect 94497 993986 94563 993989
rect 81065 993984 94563 993986
rect 81065 993928 81070 993984
rect 81126 993928 94502 993984
rect 94558 993928 94563 993984
rect 81065 993926 94563 993928
rect 81065 993923 81131 993926
rect 94497 993923 94563 993926
rect 139393 993986 139459 993989
rect 145741 993986 145807 993989
rect 139393 993984 145807 993986
rect 139393 993928 139398 993984
rect 139454 993928 145746 993984
rect 145802 993928 145807 993984
rect 139393 993926 145807 993928
rect 139393 993923 139459 993926
rect 145741 993923 145807 993926
rect 184289 993986 184355 993989
rect 186267 993986 186333 993989
rect 184289 993984 186333 993986
rect 184289 993928 184294 993984
rect 184350 993928 186272 993984
rect 186328 993928 186333 993984
rect 184289 993926 186333 993928
rect 184289 993923 184355 993926
rect 186267 993923 186333 993926
rect 132534 993788 132540 993852
rect 132604 993850 132610 993852
rect 137553 993850 137619 993853
rect 132604 993848 137619 993850
rect 132604 993792 137558 993848
rect 137614 993792 137619 993848
rect 132604 993790 137619 993792
rect 132604 993788 132610 993790
rect 137553 993787 137619 993790
rect 187417 993850 187483 993853
rect 195237 993850 195303 993853
rect 187417 993848 195303 993850
rect 187417 993792 187422 993848
rect 187478 993792 195242 993848
rect 195298 993792 195303 993848
rect 187417 993790 195303 993792
rect 187417 993787 187483 993790
rect 195237 993787 195303 993790
rect 137737 993714 137803 993717
rect 142153 993714 142219 993717
rect 137737 993712 142219 993714
rect 137737 993656 137742 993712
rect 137798 993656 142158 993712
rect 142214 993656 142219 993712
rect 137737 993654 142219 993656
rect 137737 993651 137803 993654
rect 142153 993651 142219 993654
rect 142337 993714 142403 993717
rect 152457 993714 152523 993717
rect 142337 993712 152523 993714
rect 142337 993656 142342 993712
rect 142398 993656 152462 993712
rect 152518 993656 152523 993712
rect 142337 993654 152523 993656
rect 142337 993651 142403 993654
rect 152457 993651 152523 993654
rect 139209 993442 139275 993445
rect 141918 993442 141924 993444
rect 139209 993440 141924 993442
rect 139209 993384 139214 993440
rect 139270 993384 141924 993440
rect 139209 993382 141924 993384
rect 139209 993379 139275 993382
rect 141918 993380 141924 993382
rect 141988 993380 141994 993444
rect 142286 993380 142292 993444
rect 142356 993442 142362 993444
rect 143809 993442 143875 993445
rect 142356 993440 143875 993442
rect 142356 993384 143814 993440
rect 143870 993384 143875 993440
rect 142356 993382 143875 993384
rect 142356 993380 142362 993382
rect 143809 993379 143875 993382
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 42149 967602 42215 967605
rect 42609 967602 42675 967605
rect 42149 967600 42675 967602
rect 42149 967544 42154 967600
rect 42210 967544 42614 967600
rect 42670 967544 42675 967600
rect 42149 967542 42675 967544
rect 42149 967539 42215 967542
rect 42609 967539 42675 967542
rect 41454 967132 41460 967196
rect 41524 967194 41530 967196
rect 41781 967194 41847 967197
rect 41524 967192 41847 967194
rect 41524 967136 41786 967192
rect 41842 967136 41847 967192
rect 41524 967134 41847 967136
rect 41524 967132 41530 967134
rect 41781 967131 41847 967134
rect 42149 967194 42215 967197
rect 43437 967194 43503 967197
rect 42149 967192 43503 967194
rect 42149 967136 42154 967192
rect 42210 967136 43442 967192
rect 43498 967136 43503 967192
rect 42149 967134 43503 967136
rect 42149 967131 42215 967134
rect 43437 967131 43503 967134
rect 674373 966106 674439 966109
rect 675201 966106 675267 966109
rect 674373 966104 675267 966106
rect 674373 966048 674378 966104
rect 674434 966048 675206 966104
rect 675262 966048 675267 966104
rect 674373 966046 675267 966048
rect 674373 966043 674439 966046
rect 675201 966043 675267 966046
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 42425 964746 42491 964749
rect 43437 964746 43503 964749
rect 42425 964744 43503 964746
rect 42425 964688 42430 964744
rect 42486 964688 43442 964744
rect 43498 964688 43503 964744
rect 42425 964686 43503 964688
rect 42425 964683 42491 964686
rect 43437 964683 43503 964686
rect 42425 963930 42491 963933
rect 43253 963930 43319 963933
rect 42425 963928 43319 963930
rect 42425 963872 42430 963928
rect 42486 963872 43258 963928
rect 43314 963872 43319 963928
rect 42425 963870 43319 963872
rect 42425 963867 42491 963870
rect 43253 963867 43319 963870
rect 675201 963658 675267 963661
rect 676622 963658 676628 963660
rect 675201 963656 676628 963658
rect 675201 963600 675206 963656
rect 675262 963600 676628 963656
rect 675201 963598 676628 963600
rect 675201 963595 675267 963598
rect 676622 963596 676628 963598
rect 676692 963596 676698 963660
rect 42425 963386 42491 963389
rect 43069 963386 43135 963389
rect 675385 963388 675451 963389
rect 675334 963386 675340 963388
rect 42425 963384 43135 963386
rect 42425 963328 42430 963384
rect 42486 963328 43074 963384
rect 43130 963328 43135 963384
rect 42425 963326 43135 963328
rect 675294 963326 675340 963386
rect 675404 963384 675451 963388
rect 675446 963328 675451 963384
rect 42425 963323 42491 963326
rect 43069 963323 43135 963326
rect 675334 963324 675340 963326
rect 675404 963324 675451 963328
rect 675385 963323 675451 963324
rect 42425 963114 42491 963117
rect 44265 963114 44331 963117
rect 42425 963112 44331 963114
rect 42425 963056 42430 963112
rect 42486 963056 44270 963112
rect 44326 963056 44331 963112
rect 42425 963054 44331 963056
rect 42425 963051 42491 963054
rect 44265 963051 44331 963054
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 673361 962842 673427 962845
rect 675477 962842 675543 962845
rect 673361 962840 675543 962842
rect 673361 962784 673366 962840
rect 673422 962784 675482 962840
rect 675538 962784 675543 962840
rect 673361 962782 675543 962784
rect 673361 962779 673427 962782
rect 675477 962779 675543 962782
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 673177 962570 673243 962573
rect 674925 962570 674991 962573
rect 673177 962568 674991 962570
rect 673177 962512 673182 962568
rect 673238 962512 674930 962568
rect 674986 962512 674991 962568
rect 673177 962510 674991 962512
rect 673177 962507 673243 962510
rect 674925 962507 674991 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 674649 962162 674715 962165
rect 675385 962162 675451 962165
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 674649 962160 675451 962162
rect 674649 962104 674654 962160
rect 674710 962104 675390 962160
rect 675446 962104 675451 962160
rect 674649 962102 675451 962104
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 674649 962099 674715 962102
rect 675385 962099 675451 962102
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 675201 959308 675267 959309
rect 675150 959306 675156 959308
rect 675110 959246 675156 959306
rect 675220 959304 675267 959308
rect 675262 959248 675267 959304
rect 675150 959244 675156 959246
rect 675220 959244 675267 959248
rect 675201 959243 675267 959244
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 42425 958762 42491 958765
rect 44449 958762 44515 958765
rect 42425 958760 44515 958762
rect 42425 958704 42430 958760
rect 42486 958704 44454 958760
rect 44510 958704 44515 958760
rect 42425 958702 44515 958704
rect 42425 958699 42491 958702
rect 44449 958699 44515 958702
rect 672993 958762 673059 958765
rect 675109 958762 675175 958765
rect 672993 958760 675175 958762
rect 672993 958704 672998 958760
rect 673054 958704 675114 958760
rect 675170 958704 675175 958760
rect 672993 958702 675175 958704
rect 672993 958699 673059 958702
rect 675109 958699 675175 958702
rect 41781 957812 41847 957813
rect 41781 957808 41828 957812
rect 41892 957810 41898 957812
rect 661677 957810 661743 957813
rect 675293 957810 675359 957813
rect 41781 957752 41786 957808
rect 41781 957748 41828 957752
rect 41892 957750 41938 957810
rect 661677 957808 675359 957810
rect 661677 957752 661682 957808
rect 661738 957752 675298 957808
rect 675354 957752 675359 957808
rect 661677 957750 675359 957752
rect 41892 957748 41898 957750
rect 41781 957747 41847 957748
rect 661677 957747 661743 957750
rect 675293 957747 675359 957750
rect 675753 957810 675819 957813
rect 676806 957810 676812 957812
rect 675753 957808 676812 957810
rect 675753 957752 675758 957808
rect 675814 957752 676812 957808
rect 675753 957750 676812 957752
rect 675753 957747 675819 957750
rect 676806 957748 676812 957750
rect 676876 957748 676882 957812
rect 674189 957130 674255 957133
rect 675477 957130 675543 957133
rect 674189 957128 675543 957130
rect 674189 957072 674194 957128
rect 674250 957072 675482 957128
rect 675538 957072 675543 957128
rect 674189 957070 675543 957072
rect 674189 957067 674255 957070
rect 675477 957067 675543 957070
rect 675753 956450 675819 956453
rect 676990 956450 676996 956452
rect 675753 956448 676996 956450
rect 675753 956392 675758 956448
rect 675814 956392 676996 956448
rect 675753 956390 676996 956392
rect 675753 956387 675819 956390
rect 676990 956388 676996 956390
rect 677060 956388 677066 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 41781 954680 41847 954685
rect 41781 954624 41786 954680
rect 41842 954624 41847 954680
rect 41781 954619 41847 954624
rect 41784 954413 41844 954619
rect 675017 954546 675083 954549
rect 675334 954546 675340 954548
rect 675017 954544 675340 954546
rect 675017 954488 675022 954544
rect 675078 954488 675340 954544
rect 675017 954486 675340 954488
rect 675017 954483 675083 954486
rect 675334 954484 675340 954486
rect 675404 954484 675410 954548
rect 41781 954408 41847 954413
rect 41781 954352 41786 954408
rect 41842 954352 41847 954408
rect 41781 954347 41847 954352
rect 674833 953458 674899 953461
rect 675385 953458 675451 953461
rect 674833 953456 675451 953458
rect 674833 953400 674838 953456
rect 674894 953400 675390 953456
rect 675446 953400 675451 953456
rect 674833 953398 675451 953400
rect 674833 953395 674899 953398
rect 675385 953395 675451 953398
rect 35157 952914 35223 952917
rect 41822 952914 41828 952916
rect 35157 952912 41828 952914
rect 35157 952856 35162 952912
rect 35218 952856 41828 952912
rect 35157 952854 41828 952856
rect 35157 952851 35223 952854
rect 41822 952852 41828 952854
rect 41892 952852 41898 952916
rect 37917 952506 37983 952509
rect 41454 952506 41460 952508
rect 37917 952504 41460 952506
rect 37917 952448 37922 952504
rect 37978 952448 41460 952504
rect 37917 952446 41460 952448
rect 37917 952443 37983 952446
rect 41454 952444 41460 952446
rect 41524 952444 41530 952508
rect 39297 952234 39363 952237
rect 41638 952234 41644 952236
rect 39297 952232 41644 952234
rect 39297 952176 39302 952232
rect 39358 952176 41644 952232
rect 39297 952174 41644 952176
rect 39297 952171 39363 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 40033 951690 40099 951693
rect 41270 951690 41276 951692
rect 40033 951688 41276 951690
rect 40033 951632 40038 951688
rect 40094 951632 41276 951688
rect 40033 951630 41276 951632
rect 40033 951627 40099 951630
rect 41270 951628 41276 951630
rect 41340 951628 41346 951692
rect 676622 951492 676628 951556
rect 676692 951554 676698 951556
rect 677501 951554 677567 951557
rect 676692 951552 677567 951554
rect 676692 951496 677506 951552
rect 677562 951496 677567 951552
rect 676692 951494 677567 951496
rect 676692 951492 676698 951494
rect 677501 951491 677567 951494
rect 675201 951418 675267 951421
rect 675845 951418 675911 951421
rect 675201 951416 675911 951418
rect 675201 951360 675206 951416
rect 675262 951360 675850 951416
rect 675906 951360 675911 951416
rect 675201 951358 675911 951360
rect 675201 951355 675267 951358
rect 675845 951355 675911 951358
rect 675201 951148 675267 951149
rect 675150 951146 675156 951148
rect 675110 951086 675156 951146
rect 675220 951144 675267 951148
rect 675262 951088 675267 951144
rect 675150 951084 675156 951086
rect 675220 951084 675267 951088
rect 675201 951083 675267 951084
rect 676070 950676 676076 950740
rect 676140 950738 676146 950740
rect 678237 950738 678303 950741
rect 676140 950736 678303 950738
rect 676140 950680 678242 950736
rect 678298 950680 678303 950736
rect 676140 950678 678303 950680
rect 676140 950676 676146 950678
rect 678237 950675 678303 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 664437 947338 664503 947341
rect 683113 947338 683179 947341
rect 664437 947336 683179 947338
rect 664437 947280 664442 947336
rect 664498 947280 683118 947336
rect 683174 947280 683179 947336
rect 664437 947278 683179 947280
rect 664437 947275 664503 947278
rect 683113 947275 683179 947278
rect 31753 946658 31819 946661
rect 46197 946658 46263 946661
rect 31753 946656 46263 946658
rect 31753 946600 31758 946656
rect 31814 946600 46202 946656
rect 46258 946600 46263 946656
rect 31753 946598 46263 946600
rect 31753 946595 31819 946598
rect 46197 946595 46263 946598
rect 40350 944012 40356 944076
rect 40420 944074 40426 944076
rect 42190 944074 42196 944076
rect 40420 944014 42196 944074
rect 40420 944012 40426 944014
rect 42190 944012 42196 944014
rect 42260 944012 42266 944076
rect 40718 943740 40724 943804
rect 40788 943802 40794 943804
rect 42006 943802 42012 943804
rect 40788 943742 42012 943802
rect 40788 943740 40794 943742
rect 42006 943740 42012 943742
rect 42076 943740 42082 943804
rect 45553 943530 45619 943533
rect 41492 943528 45619 943530
rect 41492 943472 45558 943528
rect 45614 943472 45619 943528
rect 41492 943470 45619 943472
rect 45553 943467 45619 943470
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 28717 942714 28783 942717
rect 28717 942712 28796 942714
rect 28717 942656 28722 942712
rect 28778 942656 28796 942712
rect 28717 942654 28796 942656
rect 28717 942651 28783 942654
rect 51717 942306 51783 942309
rect 41492 942304 51783 942306
rect 41492 942248 51722 942304
rect 51778 942248 51783 942304
rect 41492 942246 51783 942248
rect 51717 942243 51783 942246
rect 35801 941898 35867 941901
rect 35788 941896 35867 941898
rect 35788 941840 35806 941896
rect 35862 941840 35867 941896
rect 35788 941838 35867 941840
rect 35801 941835 35867 941838
rect 663057 941762 663123 941765
rect 676213 941762 676279 941765
rect 663057 941760 676279 941762
rect 663057 941704 663062 941760
rect 663118 941704 676218 941760
rect 676274 941704 676279 941760
rect 663057 941702 676279 941704
rect 663057 941699 663123 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 44633 941082 44699 941085
rect 41492 941080 44699 941082
rect 41492 941024 44638 941080
rect 44694 941024 44699 941080
rect 41492 941022 44699 941024
rect 44633 941019 44699 941022
rect 42057 940674 42123 940677
rect 41492 940672 42123 940674
rect 41492 940616 42062 940672
rect 42118 940616 42123 940672
rect 41492 940614 42123 940616
rect 42057 940611 42123 940614
rect 35801 940266 35867 940269
rect 35788 940264 35867 940266
rect 35788 940208 35806 940264
rect 35862 940208 35867 940264
rect 35788 940206 35867 940208
rect 35801 940203 35867 940206
rect 48957 940130 49023 940133
rect 41830 940128 49023 940130
rect 41830 940072 48962 940128
rect 49018 940072 49023 940128
rect 41830 940070 49023 940072
rect 41830 939858 41890 940070
rect 48957 940067 49023 940070
rect 41492 939798 41890 939858
rect 42057 939858 42123 939861
rect 50337 939858 50403 939861
rect 42057 939856 50403 939858
rect 42057 939800 42062 939856
rect 42118 939800 50342 939856
rect 50398 939800 50403 939856
rect 42057 939798 50403 939800
rect 42057 939795 42123 939798
rect 50337 939795 50403 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683113 939722 683179 939725
rect 683070 939720 683179 939722
rect 683070 939664 683118 939720
rect 683174 939664 683179 939720
rect 683070 939659 683179 939664
rect 683070 939556 683130 939659
rect 41822 939450 41828 939452
rect 41492 939390 41828 939450
rect 41822 939388 41828 939390
rect 41892 939388 41898 939452
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 36537 939042 36603 939045
rect 36524 939040 36603 939042
rect 36524 938984 36542 939040
rect 36598 938984 36603 939040
rect 36524 938982 36603 938984
rect 36537 938979 36603 938982
rect 37917 938634 37983 938637
rect 37917 938632 37996 938634
rect 37917 938576 37922 938632
rect 37978 938576 37996 938632
rect 37917 938574 37996 938576
rect 37917 938571 37983 938574
rect 668577 938498 668643 938501
rect 676262 938498 676322 938740
rect 668577 938496 676322 938498
rect 668577 938440 668582 938496
rect 668638 938440 676322 938496
rect 668577 938438 676322 938440
rect 668577 938435 668643 938438
rect 33777 938226 33843 938229
rect 33764 938224 33843 938226
rect 33764 938168 33782 938224
rect 33838 938168 33843 938224
rect 33764 938166 33843 938168
rect 33777 938163 33843 938166
rect 676446 938093 676506 938332
rect 672165 938090 672231 938093
rect 672165 938088 676322 938090
rect 672165 938032 672170 938088
rect 672226 938032 676322 938088
rect 672165 938030 676322 938032
rect 676446 938088 676555 938093
rect 676446 938032 676494 938088
rect 676550 938032 676555 938088
rect 676446 938030 676555 938032
rect 672165 938027 672231 938030
rect 676262 937924 676322 938030
rect 676489 938027 676555 938030
rect 35157 937818 35223 937821
rect 667197 937818 667263 937821
rect 672809 937818 672875 937821
rect 676029 937818 676095 937821
rect 35157 937816 35236 937818
rect 35157 937760 35162 937816
rect 35218 937760 35236 937816
rect 35157 937758 35236 937760
rect 667197 937816 672458 937818
rect 667197 937760 667202 937816
rect 667258 937760 672458 937816
rect 667197 937758 672458 937760
rect 35157 937755 35223 937758
rect 667197 937755 667263 937758
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 660297 937274 660363 937277
rect 672165 937274 672231 937277
rect 660297 937272 672231 937274
rect 660297 937216 660302 937272
rect 660358 937216 672170 937272
rect 672226 937216 672231 937272
rect 660297 937214 672231 937216
rect 672398 937274 672458 937758
rect 672809 937816 676095 937818
rect 672809 937760 672814 937816
rect 672870 937760 676034 937816
rect 676090 937760 676095 937816
rect 672809 937758 676095 937760
rect 672809 937755 672875 937758
rect 676029 937755 676095 937758
rect 672625 937546 672691 937549
rect 672625 937544 676292 937546
rect 672625 937488 672630 937544
rect 672686 937488 676292 937544
rect 672625 937486 676292 937488
rect 672625 937483 672691 937486
rect 672398 937214 676322 937274
rect 660297 937211 660363 937214
rect 672165 937211 672231 937214
rect 676262 937108 676322 937214
rect 42793 937002 42859 937005
rect 41492 937000 42859 937002
rect 41492 936944 42798 937000
rect 42854 936944 42859 937000
rect 41492 936942 42859 936944
rect 42793 936939 42859 936942
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 44449 936186 44515 936189
rect 41492 936184 44515 936186
rect 41492 936128 44454 936184
rect 44510 936128 44515 936184
rect 41492 936126 44515 936128
rect 44449 936123 44515 936126
rect 41822 935778 41828 935780
rect 41492 935718 41828 935778
rect 41822 935716 41828 935718
rect 41892 935716 41898 935780
rect 42057 935778 42123 935781
rect 64462 935778 64522 936836
rect 671797 936730 671863 936733
rect 671797 936728 676292 936730
rect 671797 936672 671802 936728
rect 671858 936672 676292 936728
rect 671797 936670 676292 936672
rect 671797 936667 671863 936670
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 42057 935776 64522 935778
rect 42057 935720 42062 935776
rect 42118 935720 64522 935776
rect 42057 935718 64522 935720
rect 671613 935778 671679 935781
rect 676262 935778 676322 935884
rect 671613 935776 676322 935778
rect 671613 935720 671618 935776
rect 671674 935720 676322 935776
rect 671613 935718 676322 935720
rect 42057 935715 42123 935718
rect 671613 935715 671679 935718
rect 678237 935642 678303 935645
rect 678237 935640 678346 935642
rect 678237 935584 678242 935640
rect 678298 935584 678346 935640
rect 678237 935579 678346 935584
rect 678286 935476 678346 935579
rect 43437 935370 43503 935373
rect 41492 935368 43503 935370
rect 41492 935312 43442 935368
rect 43498 935312 43503 935368
rect 41492 935310 43503 935312
rect 43437 935307 43503 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43069 934962 43135 934965
rect 41492 934960 43135 934962
rect 41492 934904 43074 934960
rect 43130 934904 43135 934960
rect 41492 934902 43135 934904
rect 43069 934899 43135 934902
rect 673177 934690 673243 934693
rect 673177 934688 676292 934690
rect 673177 934632 673182 934688
rect 673238 934632 676292 934688
rect 673177 934630 676292 934632
rect 673177 934627 673243 934630
rect 40033 934554 40099 934557
rect 40020 934552 40099 934554
rect 40020 934496 40038 934552
rect 40094 934496 40099 934552
rect 40020 934494 40099 934496
rect 40033 934491 40099 934494
rect 675017 934282 675083 934285
rect 675017 934280 676292 934282
rect 675017 934224 675022 934280
rect 675078 934224 676292 934280
rect 675017 934222 676292 934224
rect 675017 934219 675083 934222
rect 44265 934146 44331 934149
rect 41492 934144 44331 934146
rect 41492 934088 44270 934144
rect 44326 934088 44331 934144
rect 41492 934086 44331 934088
rect 44265 934083 44331 934086
rect 675201 933874 675267 933877
rect 675201 933872 676292 933874
rect 675201 933816 675206 933872
rect 675262 933816 676292 933872
rect 675201 933814 676292 933816
rect 675201 933811 675267 933814
rect 43253 933738 43319 933741
rect 41492 933736 43319 933738
rect 41492 933680 43258 933736
rect 43314 933680 43319 933736
rect 41492 933678 43319 933680
rect 43253 933675 43319 933678
rect 680997 933602 681063 933605
rect 680997 933600 681106 933602
rect 680997 933544 681002 933600
rect 681058 933544 681106 933600
rect 680997 933539 681106 933544
rect 681046 933436 681106 933539
rect 43345 933330 43411 933333
rect 41492 933328 43411 933330
rect 41492 933272 43350 933328
rect 43406 933272 43411 933328
rect 41492 933270 43411 933272
rect 43345 933267 43411 933270
rect 674373 933058 674439 933061
rect 674373 933056 676292 933058
rect 674373 933000 674378 933056
rect 674434 933000 676292 933056
rect 674373 932998 676292 933000
rect 674373 932995 674439 932998
rect 42241 932922 42307 932925
rect 41492 932920 42307 932922
rect 41492 932864 42246 932920
rect 42302 932864 42307 932920
rect 41492 932862 42307 932864
rect 42241 932859 42307 932862
rect 673361 932650 673427 932653
rect 673361 932648 676292 932650
rect 673361 932592 673366 932648
rect 673422 932592 676292 932648
rect 673361 932590 676292 932592
rect 673361 932587 673427 932590
rect 674649 932242 674715 932245
rect 674649 932240 676292 932242
rect 674649 932184 674654 932240
rect 674710 932184 676292 932240
rect 674649 932182 676292 932184
rect 674649 932179 674715 932182
rect 43529 932106 43595 932109
rect 41492 932104 43595 932106
rect 41492 932048 43534 932104
rect 43590 932048 43595 932104
rect 41492 932046 43595 932048
rect 43529 932043 43595 932046
rect 676990 931908 676996 931972
rect 677060 931908 677066 931972
rect 676998 931804 677058 931908
rect 676806 931500 676812 931564
rect 676876 931500 676882 931564
rect 676814 931396 676874 931500
rect 677501 931154 677567 931157
rect 677501 931152 677610 931154
rect 677501 931096 677506 931152
rect 677562 931096 677610 931152
rect 677501 931091 677610 931096
rect 677550 930988 677610 931091
rect 672993 930610 673059 930613
rect 672993 930608 676292 930610
rect 672993 930552 672998 930608
rect 673054 930552 676292 930608
rect 672993 930550 676292 930552
rect 672993 930547 673059 930550
rect 674189 930202 674255 930205
rect 674189 930200 676292 930202
rect 674189 930144 674194 930200
rect 674250 930144 676292 930200
rect 674189 930142 676292 930144
rect 674189 930139 674255 930142
rect 673361 929522 673427 929525
rect 676262 929522 676322 929764
rect 673361 929520 676322 929522
rect 673361 929464 673366 929520
rect 673422 929464 676322 929520
rect 673361 929462 676322 929464
rect 673361 929459 673427 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 671981 928298 672047 928301
rect 676262 928298 676322 928540
rect 671981 928296 676322 928298
rect 671981 928240 671986 928296
rect 672042 928240 676322 928296
rect 671981 928238 676322 928240
rect 671981 928235 672047 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 41689 911978 41755 911981
rect 42006 911978 42012 911980
rect 41689 911976 42012 911978
rect 41689 911920 41694 911976
rect 41750 911920 42012 911976
rect 41689 911918 42012 911920
rect 41689 911915 41755 911918
rect 42006 911916 42012 911918
rect 42076 911916 42082 911980
rect 41505 911706 41571 911709
rect 42190 911706 42196 911708
rect 41505 911704 42196 911706
rect 41505 911648 41510 911704
rect 41566 911648 42196 911704
rect 41505 911646 42196 911648
rect 41505 911643 41571 911646
rect 42190 911644 42196 911646
rect 42260 911644 42266 911708
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 44081 892802 44147 892805
rect 55857 892802 55923 892805
rect 44081 892800 55923 892802
rect 44081 892744 44086 892800
rect 44142 892744 55862 892800
rect 55918 892744 55923 892800
rect 44081 892742 55923 892744
rect 44081 892739 44147 892742
rect 55857 892739 55923 892742
rect 42931 892530 42997 892533
rect 54477 892530 54543 892533
rect 42931 892528 54543 892530
rect 42931 892472 42936 892528
rect 42992 892472 54482 892528
rect 54538 892472 54543 892528
rect 42931 892470 54543 892472
rect 42931 892467 42997 892470
rect 54477 892467 54543 892470
rect 43069 892258 43135 892261
rect 53281 892258 53347 892261
rect 43069 892256 53347 892258
rect 43069 892200 43074 892256
rect 43130 892200 53286 892256
rect 53342 892200 53347 892256
rect 43069 892198 53347 892200
rect 43069 892195 43135 892198
rect 53281 892195 53347 892198
rect 44081 891986 44147 891989
rect 47577 891986 47643 891989
rect 44081 891984 47643 891986
rect 44081 891928 44086 891984
rect 44142 891928 47582 891984
rect 47638 891928 47643 891984
rect 44081 891926 47643 891928
rect 44081 891923 44147 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 669221 879202 669287 879205
rect 675293 879202 675359 879205
rect 669221 879200 675359 879202
rect 669221 879144 669226 879200
rect 669282 879144 675298 879200
rect 675354 879144 675359 879200
rect 669221 879142 675359 879144
rect 669221 879139 669287 879142
rect 675293 879139 675359 879142
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 672533 873626 672599 873629
rect 675385 873626 675451 873629
rect 672533 873624 675451 873626
rect 672533 873568 672538 873624
rect 672594 873568 675390 873624
rect 675446 873568 675451 873624
rect 672533 873566 675451 873568
rect 672533 873563 672599 873566
rect 675385 873563 675451 873566
rect 673862 873156 673868 873220
rect 673932 873218 673938 873220
rect 675109 873218 675175 873221
rect 673932 873216 675175 873218
rect 673932 873160 675114 873216
rect 675170 873160 675175 873216
rect 673932 873158 675175 873160
rect 673932 873156 673938 873158
rect 675109 873155 675175 873158
rect 671153 872266 671219 872269
rect 675385 872266 675451 872269
rect 671153 872264 675451 872266
rect 671153 872208 671158 872264
rect 671214 872208 675390 872264
rect 675446 872208 675451 872264
rect 671153 872206 675451 872208
rect 671153 872203 671219 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 674925 870906 674991 870909
rect 676806 870906 676812 870908
rect 674925 870904 676812 870906
rect 674925 870848 674930 870904
rect 674986 870848 676812 870904
rect 674925 870846 676812 870848
rect 674925 870843 674991 870846
rect 676806 870844 676812 870846
rect 676876 870844 676882 870908
rect 672993 870090 673059 870093
rect 675109 870090 675175 870093
rect 672993 870088 675175 870090
rect 672993 870032 672998 870088
rect 673054 870032 675114 870088
rect 675170 870032 675175 870088
rect 672993 870030 675175 870032
rect 672993 870027 673059 870030
rect 675109 870027 675175 870030
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 664437 868730 664503 868733
rect 664437 868728 669330 868730
rect 664437 868672 664442 868728
rect 664498 868672 669330 868728
rect 664437 868670 669330 868672
rect 664437 868667 664503 868670
rect 669270 868458 669330 868670
rect 675293 868458 675359 868461
rect 669270 868456 675359 868458
rect 669270 868400 675298 868456
rect 675354 868400 675359 868456
rect 669270 868398 675359 868400
rect 675293 868395 675359 868398
rect 668209 868186 668275 868189
rect 674833 868186 674899 868189
rect 668209 868184 674899 868186
rect 668209 868128 668214 868184
rect 668270 868128 674838 868184
rect 674894 868128 674899 868184
rect 668209 868126 674899 868128
rect 668209 868123 668275 868126
rect 674833 868123 674899 868126
rect 670601 867914 670667 867917
rect 675477 867914 675543 867917
rect 670601 867912 675543 867914
rect 670601 867856 670606 867912
rect 670662 867856 675482 867912
rect 675538 867856 675543 867912
rect 670601 867854 675543 867856
rect 670601 867851 670667 867854
rect 675477 867851 675543 867854
rect 674833 867506 674899 867509
rect 675477 867506 675543 867509
rect 674833 867504 675543 867506
rect 674833 867448 674838 867504
rect 674894 867448 675482 867504
rect 675538 867448 675543 867504
rect 674833 867446 675543 867448
rect 674833 867443 674899 867446
rect 675477 867443 675543 867446
rect 673913 864922 673979 864925
rect 675385 864922 675451 864925
rect 673913 864920 675451 864922
rect 673913 864864 673918 864920
rect 673974 864864 675390 864920
rect 675446 864864 675451 864920
rect 673913 864862 675451 864864
rect 673913 864859 673979 864862
rect 675385 864859 675451 864862
rect 669773 864242 669839 864245
rect 675477 864242 675543 864245
rect 669773 864240 675543 864242
rect 669773 864184 669778 864240
rect 669834 864184 675482 864240
rect 675538 864184 675543 864240
rect 669773 864182 675543 864184
rect 669773 864179 669839 864182
rect 675477 864179 675543 864182
rect 675293 863156 675359 863157
rect 675293 863154 675340 863156
rect 675248 863152 675340 863154
rect 675248 863096 675298 863152
rect 675248 863094 675340 863096
rect 675293 863092 675340 863094
rect 675404 863092 675410 863156
rect 675293 863091 675359 863092
rect 62757 858666 62823 858669
rect 62757 858664 64492 858666
rect 62757 858608 62762 858664
rect 62818 858608 64492 858664
rect 62757 858606 64492 858608
rect 62757 858603 62823 858606
rect 652385 856354 652451 856357
rect 650164 856352 652451 856354
rect 650164 856296 652390 856352
rect 652446 856296 652451 856352
rect 650164 856294 652451 856296
rect 652385 856291 652451 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 652017 843026 652083 843029
rect 650164 843024 652083 843026
rect 650164 842968 652022 843024
rect 652078 842968 652083 843024
rect 650164 842966 652083 842968
rect 652017 842963 652083 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 35801 816506 35867 816509
rect 651465 816506 651531 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 35801 816443 35867 816446
rect 651465 816443 651531 816446
rect 44449 816098 44515 816101
rect 41492 816096 44515 816098
rect 41492 816040 44454 816096
rect 44510 816040 44515 816096
rect 41492 816038 44515 816040
rect 44449 816035 44515 816038
rect 44633 815690 44699 815693
rect 41492 815688 44699 815690
rect 41492 815632 44638 815688
rect 44694 815632 44699 815688
rect 41492 815630 44699 815632
rect 44633 815627 44699 815630
rect 44817 815282 44883 815285
rect 41492 815280 44883 815282
rect 41492 815224 44822 815280
rect 44878 815224 44883 815280
rect 41492 815222 44883 815224
rect 44817 815219 44883 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 44265 814466 44331 814469
rect 41492 814464 44331 814466
rect 41492 814408 44270 814464
rect 44326 814408 44331 814464
rect 41492 814406 44331 814408
rect 44265 814403 44331 814406
rect 39982 814234 39988 814298
rect 40052 814234 40058 814298
rect 39990 814028 40050 814234
rect 44633 813650 44699 813653
rect 41492 813648 44699 813650
rect 41492 813592 44638 813648
rect 44694 813592 44699 813648
rect 41492 813590 44699 813592
rect 44633 813587 44699 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 41321 812834 41387 812837
rect 41308 812832 41387 812834
rect 41308 812776 41326 812832
rect 41382 812776 41387 812832
rect 41308 812774 41387 812776
rect 41321 812771 41387 812774
rect 40953 812426 41019 812429
rect 40940 812424 41019 812426
rect 40940 812368 40958 812424
rect 41014 812368 41019 812424
rect 40940 812366 41019 812368
rect 40953 812363 41019 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 35157 811610 35223 811613
rect 35157 811608 35236 811610
rect 35157 811552 35162 811608
rect 35218 811552 35236 811608
rect 35157 811550 35236 811552
rect 35157 811547 35223 811550
rect 35893 811202 35959 811205
rect 35893 811200 35972 811202
rect 35893 811144 35898 811200
rect 35954 811144 35972 811200
rect 35893 811142 35972 811144
rect 35893 811139 35959 811142
rect 43161 810794 43227 810797
rect 41492 810792 43227 810794
rect 41492 810736 43166 810792
rect 43222 810736 43227 810792
rect 41492 810734 43227 810736
rect 43161 810731 43227 810734
rect 45001 810386 45067 810389
rect 41492 810384 45067 810386
rect 41492 810328 45006 810384
rect 45062 810328 45067 810384
rect 41492 810326 45067 810328
rect 45001 810323 45067 810326
rect 42793 809978 42859 809981
rect 41492 809976 42859 809978
rect 41492 809920 42798 809976
rect 42854 809920 42859 809976
rect 41492 809918 42859 809920
rect 42793 809915 42859 809918
rect 43897 809570 43963 809573
rect 41492 809568 43963 809570
rect 41492 809512 43902 809568
rect 43958 809512 43963 809568
rect 41492 809510 43963 809512
rect 43897 809507 43963 809510
rect 41781 809162 41847 809165
rect 41492 809160 41847 809162
rect 41492 809104 41786 809160
rect 41842 809104 41847 809160
rect 41492 809102 41847 809104
rect 41781 809099 41847 809102
rect 42190 808754 42196 808756
rect 41492 808694 42196 808754
rect 42190 808692 42196 808694
rect 42260 808692 42266 808756
rect 40585 808346 40651 808349
rect 40572 808344 40651 808346
rect 40572 808288 40590 808344
rect 40646 808288 40651 808344
rect 40572 808286 40651 808288
rect 40585 808283 40651 808286
rect 45185 807938 45251 807941
rect 41492 807936 45251 807938
rect 41492 807880 45190 807936
rect 45246 807880 45251 807936
rect 41492 807878 45251 807880
rect 45185 807875 45251 807878
rect 42977 807530 43043 807533
rect 41308 807528 43043 807530
rect 41308 807472 42982 807528
rect 43038 807472 43043 807528
rect 41308 807470 43043 807472
rect 42977 807467 43043 807470
rect 41462 806714 41522 807092
rect 42241 806714 42307 806717
rect 41462 806712 42307 806714
rect 41462 806684 42246 806712
rect 41492 806656 42246 806684
rect 42302 806656 42307 806712
rect 41492 806654 42307 806656
rect 42241 806651 42307 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43713 806306 43779 806309
rect 41492 806304 43779 806306
rect 41492 806248 43718 806304
rect 43774 806248 43779 806304
rect 41492 806246 43779 806248
rect 43713 806243 43779 806246
rect 41137 805626 41203 805629
rect 42006 805626 42012 805628
rect 41137 805624 42012 805626
rect 41137 805568 41142 805624
rect 41198 805568 42012 805624
rect 41137 805566 42012 805568
rect 41137 805563 41203 805566
rect 42006 805564 42012 805566
rect 42076 805564 42082 805628
rect 40769 805492 40835 805493
rect 40718 805490 40724 805492
rect 40678 805430 40724 805490
rect 40788 805488 40835 805492
rect 40830 805432 40835 805488
rect 40718 805428 40724 805430
rect 40788 805428 40835 805432
rect 40769 805427 40835 805428
rect 40953 805354 41019 805357
rect 41638 805354 41644 805356
rect 40953 805352 41644 805354
rect 40953 805296 40958 805352
rect 41014 805296 41644 805352
rect 40953 805294 41644 805296
rect 40953 805291 41019 805294
rect 41638 805292 41644 805294
rect 41708 805292 41714 805356
rect 40585 805082 40651 805085
rect 40902 805082 40908 805084
rect 40585 805080 40908 805082
rect 40585 805024 40590 805080
rect 40646 805024 40908 805080
rect 40585 805022 40908 805024
rect 40585 805019 40651 805022
rect 40902 805020 40908 805022
rect 40972 805020 40978 805084
rect 40534 804748 40540 804812
rect 40604 804810 40610 804812
rect 42190 804810 42196 804812
rect 40604 804750 42196 804810
rect 40604 804748 40610 804750
rect 42190 804748 42196 804750
rect 42260 804748 42266 804812
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41689 802498 41755 802501
rect 42517 802498 42583 802501
rect 41689 802496 42583 802498
rect 41689 802440 41694 802496
rect 41750 802440 42522 802496
rect 42578 802440 42583 802496
rect 41689 802438 42583 802440
rect 41689 802435 41755 802438
rect 42517 802435 42583 802438
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 53097 799098 53163 799101
rect 42566 799096 53163 799098
rect 42566 799040 53102 799096
rect 53158 799040 53163 799096
rect 42566 799038 53163 799040
rect 42566 798965 42626 799038
rect 53097 799035 53163 799038
rect 42517 798960 42626 798965
rect 42517 798904 42522 798960
rect 42578 798904 42626 798960
rect 42517 798902 42626 798904
rect 42517 798899 42583 798902
rect 42149 796242 42215 796245
rect 43897 796242 43963 796245
rect 42149 796240 43963 796242
rect 42149 796184 42154 796240
rect 42210 796184 43902 796240
rect 43958 796184 43963 796240
rect 42149 796182 43963 796184
rect 42149 796179 42215 796182
rect 43897 796179 43963 796182
rect 40902 795364 40908 795428
rect 40972 795426 40978 795428
rect 42517 795426 42583 795429
rect 40972 795424 42583 795426
rect 40972 795368 42522 795424
rect 42578 795368 42583 795424
rect 40972 795366 42583 795368
rect 40972 795364 40978 795366
rect 42517 795363 42583 795366
rect 42057 795018 42123 795021
rect 45185 795018 45251 795021
rect 42057 795016 45251 795018
rect 42057 794960 42062 795016
rect 42118 794960 45190 795016
rect 45246 794960 45251 795016
rect 42057 794958 45251 794960
rect 42057 794955 42123 794958
rect 45185 794955 45251 794958
rect 40718 794140 40724 794204
rect 40788 794202 40794 794204
rect 41781 794202 41847 794205
rect 40788 794200 41847 794202
rect 40788 794144 41786 794200
rect 41842 794144 41847 794200
rect 40788 794142 41847 794144
rect 40788 794140 40794 794142
rect 41781 794139 41847 794142
rect 62941 793658 63007 793661
rect 62941 793656 64492 793658
rect 62941 793600 62946 793656
rect 63002 793600 64492 793656
rect 62941 793598 64492 793600
rect 62941 793595 63007 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 669589 789442 669655 789445
rect 674925 789442 674991 789445
rect 669589 789440 674991 789442
rect 669589 789384 669594 789440
rect 669650 789384 674930 789440
rect 674986 789384 674991 789440
rect 669589 789382 674991 789384
rect 669589 789379 669655 789382
rect 674925 789379 674991 789382
rect 42149 789306 42215 789309
rect 45001 789306 45067 789309
rect 42149 789304 45067 789306
rect 42149 789248 42154 789304
rect 42210 789248 45006 789304
rect 45062 789248 45067 789304
rect 42149 789246 45067 789248
rect 42149 789243 42215 789246
rect 45001 789243 45067 789246
rect 41638 788972 41644 789036
rect 41708 789034 41714 789036
rect 42701 789034 42767 789037
rect 41708 789032 42767 789034
rect 41708 788976 42706 789032
rect 42762 788976 42767 789032
rect 41708 788974 42767 788976
rect 41708 788972 41714 788974
rect 42701 788971 42767 788974
rect 41781 788628 41847 788629
rect 41781 788624 41828 788628
rect 41892 788626 41898 788628
rect 42701 788626 42767 788629
rect 62757 788626 62823 788629
rect 41781 788568 41786 788624
rect 41781 788564 41828 788568
rect 41892 788566 41938 788626
rect 42701 788624 62823 788626
rect 42701 788568 42706 788624
rect 42762 788568 62762 788624
rect 62818 788568 62823 788624
rect 42701 788566 62823 788568
rect 41892 788564 41898 788566
rect 41781 788563 41847 788564
rect 42701 788563 42767 788566
rect 62757 788563 62823 788566
rect 42241 788218 42307 788221
rect 43161 788218 43227 788221
rect 42241 788216 43227 788218
rect 42241 788160 42246 788216
rect 42302 788160 43166 788216
rect 43222 788160 43227 788216
rect 42241 788158 43227 788160
rect 42241 788155 42307 788158
rect 43161 788155 43227 788158
rect 674465 788082 674531 788085
rect 675477 788082 675543 788085
rect 674465 788080 675543 788082
rect 674465 788024 674470 788080
rect 674526 788024 675482 788080
rect 675538 788024 675543 788080
rect 674465 788022 675543 788024
rect 674465 788019 674531 788022
rect 675477 788019 675543 788022
rect 674925 787538 674991 787541
rect 675477 787538 675543 787541
rect 674925 787536 675543 787538
rect 674925 787480 674930 787536
rect 674986 787480 675482 787536
rect 675538 787480 675543 787536
rect 674925 787478 675543 787480
rect 674925 787475 674991 787478
rect 675477 787475 675543 787478
rect 674833 787266 674899 787269
rect 675385 787266 675451 787269
rect 674833 787264 675451 787266
rect 674833 787208 674838 787264
rect 674894 787208 675390 787264
rect 675446 787208 675451 787264
rect 674833 787206 675451 787208
rect 674833 787203 674899 787206
rect 675385 787203 675451 787206
rect 41454 786796 41460 786860
rect 41524 786858 41530 786860
rect 41781 786858 41847 786861
rect 41524 786856 41847 786858
rect 41524 786800 41786 786856
rect 41842 786800 41847 786856
rect 41524 786798 41847 786800
rect 41524 786796 41530 786798
rect 41781 786795 41847 786798
rect 667749 786722 667815 786725
rect 675477 786722 675543 786725
rect 667749 786720 675543 786722
rect 667749 786664 667754 786720
rect 667810 786664 675482 786720
rect 675538 786664 675543 786720
rect 667749 786662 675543 786664
rect 667749 786659 667815 786662
rect 675477 786659 675543 786662
rect 672349 784410 672415 784413
rect 675477 784410 675543 784413
rect 672349 784408 675543 784410
rect 672349 784352 672354 784408
rect 672410 784352 675482 784408
rect 675538 784352 675543 784408
rect 672349 784350 675543 784352
rect 672349 784347 672415 784350
rect 675477 784347 675543 784350
rect 668393 783866 668459 783869
rect 675477 783866 675543 783869
rect 668393 783864 675543 783866
rect 668393 783808 668398 783864
rect 668454 783808 675482 783864
rect 675538 783808 675543 783864
rect 668393 783806 675543 783808
rect 668393 783803 668459 783806
rect 675477 783803 675543 783806
rect 670325 783050 670391 783053
rect 675477 783050 675543 783053
rect 670325 783048 675543 783050
rect 670325 782992 670330 783048
rect 670386 782992 675482 783048
rect 675538 782992 675543 783048
rect 670325 782990 675543 782992
rect 670325 782987 670391 782990
rect 675477 782987 675543 782990
rect 670969 781146 671035 781149
rect 675293 781146 675359 781149
rect 670969 781144 675359 781146
rect 670969 781088 670974 781144
rect 671030 781088 675298 781144
rect 675354 781088 675359 781144
rect 670969 781086 675359 781088
rect 670969 781083 671035 781086
rect 675293 781083 675359 781086
rect 670141 780602 670207 780605
rect 675477 780602 675543 780605
rect 670141 780600 675543 780602
rect 670141 780544 670146 780600
rect 670202 780544 675482 780600
rect 675538 780544 675543 780600
rect 670141 780542 675543 780544
rect 670141 780539 670207 780542
rect 675477 780539 675543 780542
rect 62757 780466 62823 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 62757 780403 62823 780406
rect 674281 779922 674347 779925
rect 675477 779922 675543 779925
rect 674281 779920 675543 779922
rect 674281 779864 674286 779920
rect 674342 779864 675482 779920
rect 675538 779864 675543 779920
rect 674281 779862 675543 779864
rect 674281 779859 674347 779862
rect 675477 779859 675543 779862
rect 673729 779242 673795 779245
rect 675477 779242 675543 779245
rect 673729 779240 675543 779242
rect 673729 779184 673734 779240
rect 673790 779184 675482 779240
rect 675538 779184 675543 779240
rect 673729 779182 675543 779184
rect 673729 779179 673795 779182
rect 675477 779179 675543 779182
rect 660297 778970 660363 778973
rect 660297 778968 669330 778970
rect 660297 778912 660302 778968
rect 660358 778912 669330 778968
rect 660297 778910 669330 778912
rect 660297 778907 660363 778910
rect 669270 778834 669330 778910
rect 675477 778834 675543 778837
rect 669270 778832 675543 778834
rect 669270 778776 675482 778832
rect 675538 778776 675543 778832
rect 669270 778774 675543 778776
rect 675477 778771 675543 778774
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 666277 777066 666343 777069
rect 675518 777066 675524 777068
rect 666277 777064 675524 777066
rect 666277 777008 666282 777064
rect 666338 777008 675524 777064
rect 666277 777006 675524 777008
rect 666277 777003 666343 777006
rect 675518 777004 675524 777006
rect 675588 777004 675594 777068
rect 651465 776658 651531 776661
rect 650164 776656 651531 776658
rect 650164 776600 651470 776656
rect 651526 776600 651531 776656
rect 650164 776598 651531 776600
rect 651465 776595 651531 776598
rect 675569 775708 675635 775709
rect 675518 775706 675524 775708
rect 675478 775646 675524 775706
rect 675588 775704 675635 775708
rect 675630 775648 675635 775704
rect 675518 775644 675524 775646
rect 675588 775644 675635 775648
rect 675569 775643 675635 775644
rect 675753 775572 675819 775573
rect 675702 775508 675708 775572
rect 675772 775570 675819 775572
rect 675772 775568 675864 775570
rect 675814 775512 675864 775568
rect 675772 775510 675864 775512
rect 675772 775508 675819 775510
rect 675753 775507 675819 775508
rect 675017 774618 675083 774621
rect 675017 774616 676230 774618
rect 675017 774560 675022 774616
rect 675078 774560 676230 774616
rect 675017 774558 676230 774560
rect 675017 774555 675083 774558
rect 676170 774482 676230 774558
rect 676990 774482 676996 774484
rect 41462 774346 41522 774452
rect 676170 774422 676996 774482
rect 676990 774420 676996 774422
rect 677060 774420 677066 774484
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 675109 774346 675175 774349
rect 675702 774346 675708 774348
rect 675109 774344 675708 774346
rect 675109 774288 675114 774344
rect 675170 774288 675708 774344
rect 675109 774286 675708 774288
rect 675109 774283 675175 774286
rect 675702 774284 675708 774286
rect 675772 774284 675778 774348
rect 41462 773938 41522 774044
rect 41462 773878 45570 773938
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 44449 773258 44515 773261
rect 41492 773256 44515 773258
rect 41492 773200 44454 773256
rect 44510 773200 44515 773256
rect 41492 773198 44515 773200
rect 44449 773195 44515 773198
rect 45093 772850 45159 772853
rect 41492 772848 45159 772850
rect 41492 772792 45098 772848
rect 45154 772792 45159 772848
rect 41492 772790 45159 772792
rect 45510 772850 45570 773878
rect 668945 773802 669011 773805
rect 675385 773802 675451 773805
rect 668945 773800 675451 773802
rect 668945 773744 668950 773800
rect 669006 773744 675390 773800
rect 675446 773744 675451 773800
rect 668945 773742 675451 773744
rect 668945 773739 669011 773742
rect 675385 773739 675451 773742
rect 55857 772850 55923 772853
rect 45510 772848 55923 772850
rect 45510 772792 55862 772848
rect 55918 772792 55923 772848
rect 45510 772790 55923 772792
rect 45093 772787 45159 772790
rect 55857 772787 55923 772790
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 682377 772714 682443 772717
rect 676140 772712 682443 772714
rect 676140 772656 682382 772712
rect 682438 772656 682443 772712
rect 676140 772654 682443 772656
rect 676140 772652 676146 772654
rect 682377 772651 682443 772654
rect 44817 772442 44883 772445
rect 41492 772440 44883 772442
rect 41492 772384 44822 772440
rect 44878 772384 44883 772440
rect 41492 772382 44883 772384
rect 44817 772379 44883 772382
rect 44449 772034 44515 772037
rect 41492 772032 44515 772034
rect 41492 771976 44454 772032
rect 44510 771976 44515 772032
rect 41492 771974 44515 771976
rect 44449 771971 44515 771974
rect 673913 772034 673979 772037
rect 683205 772034 683271 772037
rect 673913 772032 683271 772034
rect 673913 771976 673918 772032
rect 673974 771976 683210 772032
rect 683266 771976 683271 772032
rect 673913 771974 683271 771976
rect 673913 771971 673979 771974
rect 683205 771971 683271 771974
rect 44265 771626 44331 771629
rect 41492 771624 44331 771626
rect 41492 771568 44270 771624
rect 44326 771568 44331 771624
rect 41492 771566 44331 771568
rect 44265 771563 44331 771566
rect 44725 771218 44791 771221
rect 41492 771216 44791 771218
rect 41492 771160 44730 771216
rect 44786 771160 44791 771216
rect 41492 771158 44791 771160
rect 44725 771155 44791 771158
rect 673862 770884 673868 770948
rect 673932 770946 673938 770948
rect 683389 770946 683455 770949
rect 673932 770944 683455 770946
rect 673932 770888 683394 770944
rect 683450 770888 683455 770944
rect 673932 770886 683455 770888
rect 673932 770884 673938 770886
rect 683389 770883 683455 770886
rect 44909 770810 44975 770813
rect 41492 770808 44975 770810
rect 41492 770752 44914 770808
rect 44970 770752 44975 770808
rect 41492 770750 44975 770752
rect 44909 770747 44975 770750
rect 672165 770674 672231 770677
rect 683573 770674 683639 770677
rect 672165 770672 683639 770674
rect 672165 770616 672170 770672
rect 672226 770616 683578 770672
rect 683634 770616 683639 770672
rect 672165 770614 683639 770616
rect 672165 770611 672231 770614
rect 683573 770611 683639 770614
rect 44909 770402 44975 770405
rect 41492 770400 44975 770402
rect 41492 770344 44914 770400
rect 44970 770344 44975 770400
rect 41492 770342 44975 770344
rect 44909 770339 44975 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35574 769453 35634 769556
rect 35574 769448 35683 769453
rect 35574 769392 35622 769448
rect 35678 769392 35683 769448
rect 35574 769390 35683 769392
rect 35617 769387 35683 769390
rect 35390 769045 35450 769148
rect 35390 769040 35499 769045
rect 35801 769042 35867 769045
rect 35390 768984 35438 769040
rect 35494 768984 35499 769040
rect 35390 768982 35499 768984
rect 35433 768979 35499 768982
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 30974 768229 31034 768332
rect 30974 768224 31083 768229
rect 30974 768168 31022 768224
rect 31078 768168 31083 768224
rect 30974 768166 31083 768168
rect 31017 768163 31083 768166
rect 674833 768226 674899 768229
rect 675150 768226 675156 768228
rect 674833 768224 675156 768226
rect 674833 768168 674838 768224
rect 674894 768168 675156 768224
rect 674833 768166 675156 768168
rect 674833 768163 674899 768166
rect 675150 768164 675156 768166
rect 675220 768164 675226 768228
rect 35574 767821 35634 767924
rect 35525 767816 35634 767821
rect 35801 767818 35867 767821
rect 35525 767760 35530 767816
rect 35586 767760 35634 767816
rect 35525 767758 35634 767760
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35525 767755 35591 767758
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 44265 766730 44331 766733
rect 41492 766728 44331 766730
rect 41492 766672 44270 766728
rect 44326 766672 44331 766728
rect 41492 766670 44331 766672
rect 44265 766667 44331 766670
rect 675109 766594 675175 766597
rect 676070 766594 676076 766596
rect 675109 766592 676076 766594
rect 675109 766536 675114 766592
rect 675170 766536 676076 766592
rect 675109 766534 676076 766536
rect 675109 766531 675175 766534
rect 676070 766532 676076 766534
rect 676140 766532 676146 766596
rect 43161 766322 43227 766325
rect 41492 766320 43227 766322
rect 41492 766264 43166 766320
rect 43222 766264 43227 766320
rect 41492 766262 43227 766264
rect 43161 766259 43227 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 41321 765778 41387 765781
rect 42701 765778 42767 765781
rect 41321 765776 42767 765778
rect 41321 765720 41326 765776
rect 41382 765720 42706 765776
rect 42762 765720 42767 765776
rect 41321 765718 42767 765720
rect 41321 765715 41387 765718
rect 42701 765715 42767 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 45277 764826 45343 764829
rect 41462 764824 45343 764826
rect 41462 764768 45282 764824
rect 45338 764768 45343 764824
rect 41462 764766 45343 764768
rect 41462 764660 41522 764766
rect 45277 764763 45343 764766
rect 40033 764554 40099 764557
rect 41638 764554 41644 764556
rect 40033 764552 41644 764554
rect 40033 764496 40038 764552
rect 40094 764496 41644 764552
rect 40033 764494 41644 764496
rect 40033 764491 40099 764494
rect 41638 764492 41644 764494
rect 41708 764492 41714 764556
rect 45553 764282 45619 764285
rect 41492 764280 45619 764282
rect 41492 764224 45558 764280
rect 45614 764224 45619 764280
rect 41492 764222 45619 764224
rect 45553 764219 45619 764222
rect 37046 763333 37106 763844
rect 37046 763328 37155 763333
rect 651465 763330 651531 763333
rect 37046 763272 37094 763328
rect 37150 763272 37155 763328
rect 37046 763270 37155 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 37089 763267 37155 763270
rect 651465 763267 651531 763270
rect 46381 763058 46447 763061
rect 41492 763056 46447 763058
rect 41492 763000 46386 763056
rect 46442 763000 46447 763056
rect 41492 762998 46447 763000
rect 46381 762995 46447 762998
rect 671337 763058 671403 763061
rect 676029 763058 676095 763061
rect 671337 763056 676095 763058
rect 671337 763000 671342 763056
rect 671398 763000 676034 763056
rect 676090 763000 676095 763056
rect 671337 762998 676095 763000
rect 671337 762995 671403 762998
rect 676029 762995 676095 762998
rect 677041 761972 677107 761973
rect 676990 761908 676996 761972
rect 677060 761970 677107 761972
rect 677060 761968 677152 761970
rect 677102 761912 677152 761968
rect 677060 761910 677152 761912
rect 677060 761908 677107 761910
rect 677041 761907 677107 761908
rect 676765 761836 676831 761837
rect 676765 761832 676812 761836
rect 676876 761834 676882 761836
rect 676765 761776 676770 761832
rect 676765 761772 676812 761776
rect 676876 761774 676922 761834
rect 676876 761772 676882 761774
rect 676765 761771 676831 761772
rect 663750 761502 676292 761562
rect 663057 760882 663123 760885
rect 663750 760882 663810 761502
rect 663057 760880 663810 760882
rect 663057 760824 663062 760880
rect 663118 760824 663810 760880
rect 663057 760822 663810 760824
rect 669270 761094 676292 761154
rect 663057 760819 663123 760822
rect 661677 760474 661743 760477
rect 669270 760474 669330 761094
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 661677 760472 669330 760474
rect 661677 760416 661682 760472
rect 661738 760416 669330 760472
rect 661677 760414 669330 760416
rect 661677 760411 661743 760414
rect 672717 760338 672783 760341
rect 672717 760336 676292 760338
rect 672717 760280 672722 760336
rect 672778 760280 676292 760336
rect 672717 760278 676292 760280
rect 672717 760275 672783 760278
rect 672717 759930 672783 759933
rect 672717 759928 676292 759930
rect 672717 759872 672722 759928
rect 672778 759872 676292 759928
rect 672717 759870 676292 759872
rect 672717 759867 672783 759870
rect 683573 759522 683639 759525
rect 683573 759520 683652 759522
rect 683573 759464 683578 759520
rect 683634 759464 683652 759520
rect 683573 759462 683652 759464
rect 683573 759459 683639 759462
rect 673177 759114 673243 759117
rect 673177 759112 676292 759114
rect 673177 759056 673182 759112
rect 673238 759056 676292 759112
rect 673177 759054 676292 759056
rect 673177 759051 673243 759054
rect 671797 758706 671863 758709
rect 671797 758704 676292 758706
rect 671797 758648 671802 758704
rect 671858 758648 676292 758704
rect 671797 758646 676292 758648
rect 671797 758643 671863 758646
rect 671521 758298 671587 758301
rect 671521 758296 676292 758298
rect 671521 758240 671526 758296
rect 671582 758240 676292 758296
rect 671521 758238 676292 758240
rect 671521 758235 671587 758238
rect 40677 758162 40743 758165
rect 40677 758160 42028 758162
rect 40677 758104 40682 758160
rect 40738 758104 42028 758160
rect 40677 758102 42028 758104
rect 40677 758099 40743 758102
rect 41968 757890 42028 758102
rect 42793 757890 42859 757893
rect 41968 757888 42859 757890
rect 41968 757832 42798 757888
rect 42854 757832 42859 757888
rect 41968 757830 42859 757832
rect 42793 757827 42859 757830
rect 671705 757890 671771 757893
rect 671705 757888 676292 757890
rect 671705 757832 671710 757888
rect 671766 757832 676292 757888
rect 671705 757830 676292 757832
rect 671705 757827 671771 757830
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 671705 757482 671771 757485
rect 671705 757480 676292 757482
rect 671705 757424 671710 757480
rect 671766 757424 676292 757480
rect 671705 757422 676292 757424
rect 671705 757419 671771 757422
rect 39481 757346 39547 757349
rect 39481 757344 41844 757346
rect 39481 757288 39486 757344
rect 39542 757288 41844 757344
rect 39481 757286 41844 757288
rect 39481 757283 39547 757286
rect 41784 756669 41844 757286
rect 674649 757210 674715 757213
rect 676029 757210 676095 757213
rect 674649 757208 676095 757210
rect 674649 757152 674654 757208
rect 674710 757152 676034 757208
rect 676090 757152 676095 757208
rect 674649 757150 676095 757152
rect 674649 757147 674715 757150
rect 676029 757147 676095 757150
rect 682377 757074 682443 757077
rect 682364 757072 682443 757074
rect 682364 757016 682382 757072
rect 682438 757016 682443 757072
rect 682364 757014 682443 757016
rect 682377 757011 682443 757014
rect 41781 756664 41847 756669
rect 683297 756666 683363 756669
rect 41781 756608 41786 756664
rect 41842 756608 41847 756664
rect 41781 756603 41847 756608
rect 683284 756664 683363 756666
rect 683284 756608 683302 756664
rect 683358 756608 683363 756664
rect 683284 756606 683363 756608
rect 683297 756603 683363 756606
rect 42006 756332 42012 756396
rect 42076 756394 42082 756396
rect 46197 756394 46263 756397
rect 42076 756392 46263 756394
rect 42076 756336 46202 756392
rect 46258 756336 46263 756392
rect 42076 756334 46263 756336
rect 42076 756332 42082 756334
rect 46197 756331 46263 756334
rect 669270 756198 676292 756258
rect 669270 755173 669330 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 672993 755442 673059 755445
rect 672993 755440 676292 755442
rect 672993 755384 672998 755440
rect 673054 755384 676292 755440
rect 672993 755382 676292 755384
rect 672993 755379 673059 755382
rect 669221 755168 669330 755173
rect 669221 755112 669226 755168
rect 669282 755112 669330 755168
rect 669221 755110 669330 755112
rect 669221 755107 669287 755110
rect 677041 755034 677107 755037
rect 677028 755032 677107 755034
rect 677028 754976 677046 755032
rect 677102 754976 677107 755032
rect 677028 754974 677107 754976
rect 677041 754971 677107 754974
rect 40902 754836 40908 754900
rect 40972 754898 40978 754900
rect 40972 754838 42442 754898
rect 40972 754836 40978 754838
rect 42382 754221 42442 754838
rect 676765 754626 676831 754629
rect 676765 754624 676844 754626
rect 676765 754568 676770 754624
rect 676826 754568 676844 754624
rect 676765 754566 676844 754568
rect 676765 754563 676831 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 42333 754216 42442 754221
rect 42333 754160 42338 754216
rect 42394 754160 42442 754216
rect 42333 754158 42442 754160
rect 672533 754218 672599 754221
rect 672533 754216 676292 754218
rect 672533 754160 672538 754216
rect 672594 754160 676292 754216
rect 672533 754158 676292 754160
rect 42333 754155 42399 754158
rect 672533 754155 672599 754158
rect 41965 754084 42031 754085
rect 41965 754080 42012 754084
rect 42076 754082 42082 754084
rect 41965 754024 41970 754080
rect 41965 754020 42012 754024
rect 42076 754022 42122 754082
rect 42076 754020 42082 754022
rect 41965 754019 42031 754020
rect 683481 753810 683547 753813
rect 683468 753808 683547 753810
rect 683468 753752 683486 753808
rect 683542 753752 683547 753808
rect 683468 753750 683547 753752
rect 683481 753747 683547 753750
rect 45277 753538 45343 753541
rect 42198 753536 45343 753538
rect 42198 753480 45282 753536
rect 45338 753480 45343 753536
rect 42198 753478 45343 753480
rect 42198 753450 42304 753478
rect 45277 753475 45343 753478
rect 42244 753268 42304 753450
rect 42190 753204 42196 753268
rect 42260 753206 42304 753268
rect 669270 753342 676292 753402
rect 42260 753204 42266 753206
rect 42057 752994 42123 752997
rect 43161 752994 43227 752997
rect 42057 752992 43227 752994
rect 42057 752936 42062 752992
rect 42118 752936 43166 752992
rect 43222 752936 43227 752992
rect 42057 752934 43227 752936
rect 42057 752931 42123 752934
rect 43161 752931 43227 752934
rect 668209 752314 668275 752317
rect 669270 752314 669330 753342
rect 683113 752994 683179 752997
rect 683100 752992 683179 752994
rect 683100 752936 683118 752992
rect 683174 752936 683179 752992
rect 683100 752934 683179 752936
rect 683113 752931 683179 752934
rect 671153 752586 671219 752589
rect 671153 752584 676292 752586
rect 671153 752528 671158 752584
rect 671214 752528 676292 752584
rect 671153 752526 676292 752528
rect 671153 752523 671219 752526
rect 668209 752312 669330 752314
rect 668209 752256 668214 752312
rect 668270 752256 669330 752312
rect 668209 752254 669330 752256
rect 668209 752251 668275 752254
rect 673913 752178 673979 752181
rect 673913 752176 676292 752178
rect 673913 752120 673918 752176
rect 673974 752120 676292 752176
rect 673913 752118 676292 752120
rect 673913 752115 673979 752118
rect 42149 751772 42215 751773
rect 42149 751770 42196 751772
rect 42104 751768 42196 751770
rect 42104 751712 42154 751768
rect 42104 751710 42196 751712
rect 42149 751708 42196 751710
rect 42260 751708 42266 751772
rect 670601 751770 670667 751773
rect 670601 751768 676292 751770
rect 670601 751712 670606 751768
rect 670662 751712 676292 751768
rect 670601 751710 676292 751712
rect 42149 751707 42215 751708
rect 670601 751707 670667 751710
rect 672901 751362 672967 751365
rect 672901 751360 676292 751362
rect 672901 751304 672906 751360
rect 672962 751304 676292 751360
rect 672901 751302 676292 751304
rect 672901 751299 672967 751302
rect 669773 750954 669839 750957
rect 669773 750952 676292 750954
rect 669773 750896 669778 750952
rect 669834 750924 676292 750952
rect 669834 750896 676322 750924
rect 669773 750894 676322 750896
rect 669773 750891 669839 750894
rect 42241 750546 42307 750549
rect 42793 750546 42859 750549
rect 42241 750544 42859 750546
rect 42241 750488 42246 750544
rect 42302 750488 42798 750544
rect 42854 750488 42859 750544
rect 676262 750516 676322 750894
rect 42241 750486 42859 750488
rect 42241 750483 42307 750486
rect 42793 750483 42859 750486
rect 40718 750348 40724 750412
rect 40788 750410 40794 750412
rect 41781 750410 41847 750413
rect 40788 750408 41847 750410
rect 40788 750352 41786 750408
rect 41842 750352 41847 750408
rect 40788 750350 41847 750352
rect 40788 750348 40794 750350
rect 41781 750347 41847 750350
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 670785 750138 670851 750141
rect 670785 750136 676292 750138
rect 670785 750080 670790 750136
rect 670846 750080 676292 750136
rect 670785 750078 676292 750080
rect 670785 750075 670851 750078
rect 40534 747356 40540 747420
rect 40604 747418 40610 747420
rect 41781 747418 41847 747421
rect 40604 747416 41847 747418
rect 40604 747360 41786 747416
rect 41842 747360 41847 747416
rect 40604 747358 41847 747360
rect 40604 747356 40610 747358
rect 41781 747355 41847 747358
rect 42149 746738 42215 746741
rect 44265 746738 44331 746741
rect 42149 746736 44331 746738
rect 42149 746680 42154 746736
rect 42210 746680 44270 746736
rect 44326 746680 44331 746736
rect 42149 746678 44331 746680
rect 42149 746675 42215 746678
rect 44265 746675 44331 746678
rect 41638 745044 41644 745108
rect 41708 745106 41714 745108
rect 42425 745106 42491 745109
rect 41708 745104 42491 745106
rect 41708 745048 42430 745104
rect 42486 745048 42491 745104
rect 41708 745046 42491 745048
rect 41708 745044 41714 745046
rect 42425 745043 42491 745046
rect 41822 744772 41828 744836
rect 41892 744834 41898 744836
rect 42241 744834 42307 744837
rect 41892 744832 42307 744834
rect 41892 744776 42246 744832
rect 42302 744776 42307 744832
rect 41892 744774 42307 744776
rect 41892 744772 41898 744774
rect 42241 744771 42307 744774
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 667565 743202 667631 743205
rect 675109 743202 675175 743205
rect 667565 743200 675175 743202
rect 667565 743144 667570 743200
rect 667626 743144 675114 743200
rect 675170 743144 675175 743200
rect 667565 743142 675175 743144
rect 667565 743139 667631 743142
rect 675109 743139 675175 743142
rect 42609 743066 42675 743069
rect 62757 743066 62823 743069
rect 42609 743064 62823 743066
rect 42609 743008 42614 743064
rect 42670 743008 62762 743064
rect 62818 743008 62823 743064
rect 42609 743006 62823 743008
rect 42609 743003 42675 743006
rect 62757 743003 62823 743006
rect 666461 742794 666527 742797
rect 674925 742794 674991 742797
rect 666461 742792 674991 742794
rect 666461 742736 666466 742792
rect 666522 742736 674930 742792
rect 674986 742736 674991 742792
rect 666461 742734 674991 742736
rect 666461 742731 666527 742734
rect 674925 742731 674991 742734
rect 674414 742460 674420 742524
rect 674484 742522 674490 742524
rect 675385 742522 675451 742525
rect 674484 742520 675451 742522
rect 674484 742464 675390 742520
rect 675446 742464 675451 742520
rect 674484 742462 675451 742464
rect 674484 742460 674490 742462
rect 675385 742459 675451 742462
rect 42425 741706 42491 741709
rect 62941 741706 63007 741709
rect 42425 741704 63007 741706
rect 42425 741648 42430 741704
rect 42486 741648 62946 741704
rect 63002 741648 63007 741704
rect 42425 741646 63007 741648
rect 42425 741643 42491 741646
rect 62941 741643 63007 741646
rect 674230 741508 674236 741572
rect 674300 741570 674306 741572
rect 675109 741570 675175 741573
rect 674300 741568 675175 741570
rect 674300 741512 675114 741568
rect 675170 741512 675175 741568
rect 674300 741510 675175 741512
rect 674300 741508 674306 741510
rect 675109 741507 675175 741510
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 669405 741162 669471 741165
rect 674925 741162 674991 741165
rect 669405 741160 674991 741162
rect 669405 741104 669410 741160
rect 669466 741104 674930 741160
rect 674986 741104 674991 741160
rect 669405 741102 674991 741104
rect 669405 741099 669471 741102
rect 674925 741099 674991 741102
rect 674598 739604 674604 739668
rect 674668 739666 674674 739668
rect 675109 739666 675175 739669
rect 674668 739664 675175 739666
rect 674668 739608 675114 739664
rect 675170 739608 675175 739664
rect 674668 739606 675175 739608
rect 674668 739604 674674 739606
rect 675109 739603 675175 739606
rect 669773 738578 669839 738581
rect 675017 738578 675083 738581
rect 669773 738576 675083 738578
rect 669773 738520 669778 738576
rect 669834 738520 675022 738576
rect 675078 738520 675083 738576
rect 669773 738518 675083 738520
rect 669773 738515 669839 738518
rect 675017 738515 675083 738518
rect 675201 738374 675267 738377
rect 675158 738372 675267 738374
rect 675158 738316 675206 738372
rect 675262 738316 675267 738372
rect 675158 738311 675267 738316
rect 672533 738306 672599 738309
rect 675158 738306 675218 738311
rect 672533 738304 675218 738306
rect 672533 738248 672538 738304
rect 672594 738248 675218 738304
rect 672533 738246 675218 738248
rect 672533 738243 672599 738246
rect 671153 737082 671219 737085
rect 675109 737082 675175 737085
rect 671153 737080 675175 737082
rect 671153 737024 671158 737080
rect 671214 737024 675114 737080
rect 675170 737024 675175 737080
rect 671153 737022 675175 737024
rect 671153 737019 671219 737022
rect 675109 737019 675175 737022
rect 652569 736810 652635 736813
rect 650164 736808 652635 736810
rect 650164 736752 652574 736808
rect 652630 736752 652635 736808
rect 650164 736750 652635 736752
rect 652569 736747 652635 736750
rect 668761 734362 668827 734365
rect 674925 734362 674991 734365
rect 668761 734360 674991 734362
rect 668761 734304 668766 734360
rect 668822 734304 674930 734360
rect 674986 734304 674991 734360
rect 668761 734302 674991 734304
rect 668761 734299 668827 734302
rect 674925 734299 674991 734302
rect 672165 733954 672231 733957
rect 675109 733954 675175 733957
rect 672165 733952 675175 733954
rect 672165 733896 672170 733952
rect 672226 733896 675114 733952
rect 675170 733896 675175 733952
rect 672165 733894 675175 733896
rect 672165 733891 672231 733894
rect 675109 733891 675175 733894
rect 668209 733682 668275 733685
rect 675109 733682 675175 733685
rect 668209 733680 675175 733682
rect 668209 733624 668214 733680
rect 668270 733624 675114 733680
rect 675170 733624 675175 733680
rect 668209 733622 675175 733624
rect 668209 733619 668275 733622
rect 675109 733619 675175 733622
rect 671981 732868 672047 732869
rect 673361 732868 673427 732869
rect 671981 732864 672028 732868
rect 672092 732866 672098 732868
rect 673310 732866 673316 732868
rect 671981 732808 671986 732864
rect 671981 732804 672028 732808
rect 672092 732806 672138 732866
rect 673270 732806 673316 732866
rect 673380 732864 673427 732868
rect 673422 732808 673427 732864
rect 672092 732804 672098 732806
rect 673310 732804 673316 732806
rect 673380 732804 673427 732808
rect 671981 732803 672047 732804
rect 673361 732803 673427 732804
rect 668761 731506 668827 731509
rect 675109 731506 675175 731509
rect 668761 731504 675175 731506
rect 668761 731448 668766 731504
rect 668822 731448 675114 731504
rect 675170 731448 675175 731504
rect 668761 731446 675175 731448
rect 668761 731443 668827 731446
rect 675109 731443 675175 731446
rect 35617 731370 35683 731373
rect 35604 731368 35683 731370
rect 35604 731312 35622 731368
rect 35678 731312 35683 731368
rect 35604 731310 35683 731312
rect 35617 731307 35683 731310
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 671061 730554 671127 730557
rect 675477 730554 675543 730557
rect 671061 730552 675543 730554
rect 671061 730496 671066 730552
rect 671122 730496 675482 730552
rect 675538 730496 675543 730552
rect 671061 730494 675543 730496
rect 671061 730491 671127 730494
rect 675477 730491 675543 730494
rect 45093 730146 45159 730149
rect 41492 730144 45159 730146
rect 41492 730088 45098 730144
rect 45154 730088 45159 730144
rect 41492 730086 45159 730088
rect 45093 730083 45159 730086
rect 673361 730146 673427 730149
rect 675293 730146 675359 730149
rect 673361 730144 675359 730146
rect 673361 730088 673366 730144
rect 673422 730088 675298 730144
rect 675354 730088 675359 730144
rect 673361 730086 675359 730088
rect 673361 730083 673427 730086
rect 675293 730083 675359 730086
rect 675886 729948 675892 730012
rect 675956 730010 675962 730012
rect 676806 730010 676812 730012
rect 675956 729950 676812 730010
rect 675956 729948 675962 729950
rect 676806 729948 676812 729950
rect 676876 729948 676882 730012
rect 44265 729738 44331 729741
rect 41492 729736 44331 729738
rect 41492 729680 44270 729736
rect 44326 729680 44331 729736
rect 41492 729678 44331 729680
rect 44265 729675 44331 729678
rect 44449 729330 44515 729333
rect 41492 729328 44515 729330
rect 41492 729272 44454 729328
rect 44510 729272 44515 729328
rect 41492 729270 44515 729272
rect 44449 729267 44515 729270
rect 44541 728922 44607 728925
rect 41492 728920 44607 728922
rect 41492 728864 44546 728920
rect 44602 728864 44607 728920
rect 41492 728862 44607 728864
rect 44541 728859 44607 728862
rect 44725 728514 44791 728517
rect 673361 728516 673427 728517
rect 41492 728512 44791 728514
rect 41492 728456 44730 728512
rect 44786 728456 44791 728512
rect 41492 728454 44791 728456
rect 44725 728451 44791 728454
rect 673310 728452 673316 728516
rect 673380 728514 673427 728516
rect 673380 728512 673472 728514
rect 673422 728456 673472 728512
rect 673380 728454 673472 728456
rect 673380 728452 673427 728454
rect 673361 728451 673427 728452
rect 62757 728242 62823 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 62757 728179 62823 728182
rect 672022 728180 672028 728244
rect 672092 728242 672098 728244
rect 673821 728242 673887 728245
rect 672092 728240 673887 728242
rect 672092 728184 673826 728240
rect 673882 728184 673887 728240
rect 672092 728182 673887 728184
rect 672092 728180 672098 728182
rect 673821 728179 673887 728182
rect 44725 728106 44791 728109
rect 41492 728104 44791 728106
rect 41492 728048 44730 728104
rect 44786 728048 44791 728104
rect 41492 728046 44791 728048
rect 44725 728043 44791 728046
rect 670785 727970 670851 727973
rect 674143 727970 674209 727973
rect 670785 727968 674209 727970
rect 670785 727912 670790 727968
rect 670846 727912 674148 727968
rect 674204 727912 674209 727968
rect 670785 727910 674209 727912
rect 670785 727907 670851 727910
rect 674143 727907 674209 727910
rect 44909 727698 44975 727701
rect 41492 727696 44975 727698
rect 41492 727640 44914 727696
rect 44970 727640 44975 727696
rect 41492 727638 44975 727640
rect 44909 727635 44975 727638
rect 673821 727698 673887 727701
rect 674741 727698 674807 727701
rect 673821 727696 674807 727698
rect 673821 727640 673826 727696
rect 673882 727640 674746 727696
rect 674802 727640 674807 727696
rect 673821 727638 674807 727640
rect 673821 727635 673887 727638
rect 674741 727635 674807 727638
rect 45093 727290 45159 727293
rect 41492 727288 45159 727290
rect 41492 727232 45098 727288
rect 45154 727232 45159 727288
rect 41492 727230 45159 727232
rect 45093 727227 45159 727230
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 674281 726882 674347 726885
rect 683481 726882 683547 726885
rect 674281 726880 683547 726882
rect 674281 726824 674286 726880
rect 674342 726824 683486 726880
rect 683542 726824 683547 726880
rect 674281 726822 683547 726824
rect 674281 726819 674347 726822
rect 683481 726819 683547 726822
rect 674005 726610 674071 726613
rect 674557 726610 674623 726613
rect 674005 726608 674114 726610
rect 674005 726552 674010 726608
rect 674066 726552 674114 726608
rect 674005 726547 674114 726552
rect 674557 726608 674666 726610
rect 674557 726552 674562 726608
rect 674618 726552 674666 726608
rect 674557 726547 674666 726552
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 41321 726411 41387 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 674054 725522 674114 726547
rect 674606 726474 674666 726547
rect 683665 726474 683731 726477
rect 674606 726472 683731 726474
rect 674606 726416 683670 726472
rect 683726 726416 683731 726472
rect 674606 726414 683731 726416
rect 683665 726411 683731 726414
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 682377 725794 682443 725797
rect 676140 725792 682443 725794
rect 676140 725736 682382 725792
rect 682438 725736 682443 725792
rect 676140 725734 682443 725736
rect 676140 725732 676146 725734
rect 682377 725731 682443 725734
rect 683849 725522 683915 725525
rect 674054 725520 683915 725522
rect 674054 725464 683854 725520
rect 683910 725464 683915 725520
rect 674054 725462 683915 725464
rect 683849 725459 683915 725462
rect 31017 725250 31083 725253
rect 31004 725248 31083 725250
rect 31004 725192 31022 725248
rect 31078 725192 31083 725248
rect 31004 725190 31083 725192
rect 31017 725187 31083 725190
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 40677 724434 40743 724437
rect 40677 724432 40756 724434
rect 40677 724376 40682 724432
rect 40738 724376 40756 724432
rect 40677 724374 40756 724376
rect 40677 724371 40743 724374
rect 673545 724162 673611 724165
rect 683297 724162 683363 724165
rect 673545 724160 683363 724162
rect 673545 724104 673550 724160
rect 673606 724104 683302 724160
rect 683358 724104 683363 724160
rect 673545 724102 683363 724104
rect 673545 724099 673611 724102
rect 683297 724099 683363 724102
rect 33041 724026 33107 724029
rect 33028 724024 33107 724026
rect 33028 723968 33046 724024
rect 33102 723968 33107 724024
rect 33028 723966 33107 723968
rect 33041 723963 33107 723966
rect 43161 723618 43227 723621
rect 41492 723616 43227 723618
rect 41492 723560 43166 723616
rect 43222 723560 43227 723616
rect 41492 723558 43227 723560
rect 43161 723555 43227 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 33777 723210 33843 723213
rect 33764 723208 33843 723210
rect 33764 723152 33782 723208
rect 33838 723152 33843 723208
rect 33764 723150 33843 723152
rect 33777 723147 33843 723150
rect 44173 722802 44239 722805
rect 41492 722800 44239 722802
rect 41492 722744 44178 722800
rect 44234 722744 44239 722800
rect 41492 722742 44239 722744
rect 44173 722739 44239 722742
rect 41822 722394 41828 722396
rect 41492 722334 41828 722394
rect 41822 722332 41828 722334
rect 41892 722332 41898 722396
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 43897 721578 43963 721581
rect 41492 721576 43963 721578
rect 41492 721520 43902 721576
rect 43958 721520 43963 721576
rect 41492 721518 43963 721520
rect 43897 721515 43963 721518
rect 44725 721170 44791 721173
rect 41492 721168 44791 721170
rect 41492 721112 44730 721168
rect 44786 721112 44791 721168
rect 41492 721110 44791 721112
rect 44725 721107 44791 721110
rect 41321 720354 41387 720357
rect 41308 720352 41387 720354
rect 41308 720296 41326 720352
rect 41382 720296 41387 720352
rect 41308 720294 41387 720296
rect 41321 720291 41387 720294
rect 46933 719946 46999 719949
rect 41492 719944 46999 719946
rect 41492 719888 46938 719944
rect 46994 719888 46999 719944
rect 41492 719886 46999 719888
rect 46933 719883 46999 719886
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41822 718586 41828 718588
rect 40604 718526 41828 718586
rect 40604 718524 40610 718526
rect 41822 718524 41828 718526
rect 41892 718524 41898 718588
rect 652017 718314 652083 718317
rect 676029 718314 676095 718317
rect 652017 718312 676095 718314
rect 652017 718256 652022 718312
rect 652078 718256 676034 718312
rect 676090 718256 676095 718312
rect 652017 718254 676095 718256
rect 652017 718251 652083 718254
rect 676029 718251 676095 718254
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 663750 716078 676292 716138
rect 658917 716002 658983 716005
rect 663750 716002 663810 716078
rect 658917 716000 663810 716002
rect 658917 715944 658922 716000
rect 658978 715944 663810 716000
rect 658917 715942 663810 715944
rect 658917 715939 658983 715942
rect 41597 715866 41663 715869
rect 42701 715866 42767 715869
rect 41597 715864 42767 715866
rect 41597 715808 41602 715864
rect 41658 715808 42706 715864
rect 42762 715808 42767 715864
rect 41597 715806 42767 715808
rect 41597 715803 41663 715806
rect 42701 715803 42767 715806
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 41873 715594 41939 715597
rect 42609 715594 42675 715597
rect 41873 715592 42675 715594
rect 41873 715536 41878 715592
rect 41934 715536 42614 715592
rect 42670 715536 42675 715592
rect 41873 715534 42675 715536
rect 41873 715531 41939 715534
rect 42609 715531 42675 715534
rect 62113 715322 62179 715325
rect 672809 715322 672875 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 672809 715320 676292 715322
rect 672809 715264 672814 715320
rect 672870 715264 676292 715320
rect 672809 715262 676292 715264
rect 62113 715259 62179 715262
rect 672809 715259 672875 715262
rect 672809 714914 672875 714917
rect 672809 714912 676292 714914
rect 672809 714856 672814 714912
rect 672870 714856 676292 714912
rect 672809 714854 676292 714856
rect 672809 714851 672875 714854
rect 40677 714778 40743 714781
rect 42006 714778 42012 714780
rect 40677 714776 42012 714778
rect 40677 714720 40682 714776
rect 40738 714720 42012 714776
rect 40677 714718 42012 714720
rect 40677 714715 40743 714718
rect 42006 714716 42012 714718
rect 42076 714716 42082 714780
rect 41822 714444 41828 714508
rect 41892 714506 41898 714508
rect 42057 714506 42123 714509
rect 41892 714504 42123 714506
rect 41892 714448 42062 714504
rect 42118 714448 42123 714504
rect 41892 714446 42123 714448
rect 41892 714444 41898 714446
rect 42057 714443 42123 714446
rect 673177 714506 673243 714509
rect 673177 714504 676292 714506
rect 673177 714448 673182 714504
rect 673238 714448 676292 714504
rect 673177 714446 676292 714448
rect 673177 714443 673243 714446
rect 41321 714236 41387 714237
rect 41270 714172 41276 714236
rect 41340 714234 41387 714236
rect 41340 714232 41432 714234
rect 41382 714176 41432 714232
rect 41340 714174 41432 714176
rect 41340 714172 41387 714174
rect 41321 714171 41387 714172
rect 672993 714098 673059 714101
rect 672993 714096 676292 714098
rect 672993 714040 672998 714096
rect 673054 714040 676292 714096
rect 672993 714038 676292 714040
rect 672993 714035 673059 714038
rect 41781 713962 41847 713965
rect 41781 713960 41890 713962
rect 41781 713904 41786 713960
rect 41842 713904 41890 713960
rect 41781 713899 41890 713904
rect 41830 713557 41890 713899
rect 671521 713690 671587 713693
rect 671521 713688 676292 713690
rect 671521 713632 671526 713688
rect 671582 713632 676292 713688
rect 671521 713630 676292 713632
rect 671521 713627 671587 713630
rect 41781 713552 41890 713557
rect 41781 713496 41786 713552
rect 41842 713496 41890 713552
rect 41781 713494 41890 713496
rect 41781 713491 41847 713494
rect 42057 713282 42123 713285
rect 42374 713282 42380 713284
rect 42057 713280 42380 713282
rect 42057 713224 42062 713280
rect 42118 713224 42380 713280
rect 42057 713222 42380 713224
rect 42057 713219 42123 713222
rect 42374 713220 42380 713222
rect 42444 713220 42450 713284
rect 671521 713282 671587 713285
rect 671521 713280 676292 713282
rect 671521 713224 671526 713280
rect 671582 713224 676292 713280
rect 671521 713222 676292 713224
rect 671521 713219 671587 713222
rect 671705 712874 671771 712877
rect 671705 712872 676292 712874
rect 671705 712816 671710 712872
rect 671766 712816 676292 712872
rect 671705 712814 676292 712816
rect 671705 712811 671771 712814
rect 670785 712466 670851 712469
rect 670785 712464 676292 712466
rect 670785 712408 670790 712464
rect 670846 712408 676292 712464
rect 670785 712406 676292 712408
rect 670785 712403 670851 712406
rect 41270 712132 41276 712196
rect 41340 712194 41346 712196
rect 41781 712194 41847 712197
rect 47577 712194 47643 712197
rect 41340 712192 41847 712194
rect 41340 712136 41786 712192
rect 41842 712136 41847 712192
rect 41340 712134 41847 712136
rect 41340 712132 41346 712134
rect 41781 712131 41847 712134
rect 42198 712192 47643 712194
rect 42198 712136 47582 712192
rect 47638 712136 47643 712192
rect 42198 712134 47643 712136
rect 42198 710837 42258 712134
rect 47577 712131 47643 712134
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 682377 711650 682443 711653
rect 682364 711648 682443 711650
rect 682364 711592 682382 711648
rect 682438 711592 682443 711648
rect 682364 711590 682443 711592
rect 682377 711587 682443 711590
rect 683665 711242 683731 711245
rect 683652 711240 683731 711242
rect 683652 711184 683670 711240
rect 683726 711184 683731 711240
rect 683652 711182 683731 711184
rect 683665 711179 683731 711182
rect 42701 711106 42767 711109
rect 43897 711106 43963 711109
rect 42701 711104 43963 711106
rect 42701 711048 42706 711104
rect 42762 711048 43902 711104
rect 43958 711048 43963 711104
rect 42701 711046 43963 711048
rect 42701 711043 42767 711046
rect 43897 711043 43963 711046
rect 42149 710832 42258 710837
rect 42149 710776 42154 710832
rect 42210 710776 42258 710832
rect 42149 710774 42258 710776
rect 667749 710834 667815 710837
rect 667749 710832 676292 710834
rect 667749 710776 667754 710832
rect 667810 710776 676292 710832
rect 667749 710774 676292 710776
rect 42149 710771 42215 710774
rect 667749 710771 667815 710774
rect 670141 710426 670207 710429
rect 670141 710424 676292 710426
rect 670141 710368 670146 710424
rect 670202 710368 676292 710424
rect 670141 710366 676292 710368
rect 670141 710363 670207 710366
rect 652569 710290 652635 710293
rect 650164 710288 652635 710290
rect 650164 710232 652574 710288
rect 652630 710232 652635 710288
rect 650164 710230 652635 710232
rect 652569 710227 652635 710230
rect 668945 710018 669011 710021
rect 668945 710016 676292 710018
rect 668945 709960 668950 710016
rect 669006 709960 676292 710016
rect 668945 709958 676292 709960
rect 668945 709955 669011 709958
rect 41873 709884 41939 709885
rect 41822 709820 41828 709884
rect 41892 709882 41939 709884
rect 41892 709880 41984 709882
rect 41934 709824 41984 709880
rect 41892 709822 41984 709824
rect 41892 709820 41939 709822
rect 41873 709819 41939 709820
rect 669589 709610 669655 709613
rect 669589 709608 676292 709610
rect 669589 709552 669594 709608
rect 669650 709552 676292 709608
rect 669589 709550 676292 709552
rect 669589 709547 669655 709550
rect 672349 709202 672415 709205
rect 672349 709200 676292 709202
rect 672349 709144 672354 709200
rect 672410 709144 676292 709200
rect 672349 709142 676292 709144
rect 672349 709139 672415 709142
rect 668393 708794 668459 708797
rect 668393 708792 676292 708794
rect 668393 708736 668398 708792
rect 668454 708736 676292 708792
rect 668393 708734 676292 708736
rect 668393 708731 668459 708734
rect 42701 708658 42767 708661
rect 42198 708656 42767 708658
rect 42198 708600 42706 708656
rect 42762 708600 42767 708656
rect 42198 708598 42767 708600
rect 42198 708525 42258 708598
rect 42701 708595 42767 708598
rect 42149 708520 42258 708525
rect 42149 708464 42154 708520
rect 42210 708464 42258 708520
rect 42149 708462 42258 708464
rect 42149 708459 42215 708462
rect 683849 708386 683915 708389
rect 683836 708384 683915 708386
rect 683836 708328 683854 708384
rect 683910 708328 683915 708384
rect 683836 708326 683915 708328
rect 683849 708323 683915 708326
rect 683297 707978 683363 707981
rect 683284 707976 683363 707978
rect 683284 707920 683302 707976
rect 683358 707920 683363 707976
rect 683284 707918 683363 707920
rect 683297 707915 683363 707918
rect 42057 707706 42123 707709
rect 44173 707706 44239 707709
rect 42057 707704 44239 707706
rect 42057 707648 42062 707704
rect 42118 707648 44178 707704
rect 44234 707648 44239 707704
rect 42057 707646 44239 707648
rect 42057 707643 42123 707646
rect 44173 707643 44239 707646
rect 670325 707570 670391 707573
rect 670325 707568 676292 707570
rect 670325 707512 670330 707568
rect 670386 707512 676292 707568
rect 670325 707510 676292 707512
rect 670325 707507 670391 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 42374 707372 42380 707436
rect 42444 707434 42450 707436
rect 42701 707434 42767 707437
rect 42444 707432 42767 707434
rect 42444 707376 42706 707432
rect 42762 707376 42767 707432
rect 42444 707374 42767 707376
rect 42444 707372 42450 707374
rect 42701 707371 42767 707374
rect 683481 707162 683547 707165
rect 683468 707160 683547 707162
rect 683468 707104 683486 707160
rect 683542 707104 683547 707160
rect 683468 707102 683547 707104
rect 683481 707099 683547 707102
rect 42057 706754 42123 706757
rect 42517 706754 42583 706757
rect 42057 706752 42583 706754
rect 42057 706696 42062 706752
rect 42118 706696 42522 706752
rect 42578 706696 42583 706752
rect 42057 706694 42583 706696
rect 42057 706691 42123 706694
rect 42517 706691 42583 706694
rect 670969 706754 671035 706757
rect 670969 706752 676292 706754
rect 670969 706696 670974 706752
rect 671030 706696 676292 706752
rect 670969 706694 676292 706696
rect 670969 706691 671035 706694
rect 40534 706420 40540 706484
rect 40604 706482 40610 706484
rect 42241 706482 42307 706485
rect 40604 706480 42307 706482
rect 40604 706424 42246 706480
rect 42302 706424 42307 706480
rect 40604 706422 42307 706424
rect 40604 706420 40610 706422
rect 42241 706419 42307 706422
rect 674373 706346 674439 706349
rect 674373 706344 676292 706346
rect 674373 706288 674378 706344
rect 674434 706288 676292 706344
rect 674373 706286 676292 706288
rect 674373 706283 674439 706286
rect 666277 705530 666343 705533
rect 676262 705530 676322 705908
rect 666277 705528 676322 705530
rect 666277 705472 666282 705528
rect 666338 705500 676322 705528
rect 666338 705472 676292 705500
rect 666277 705470 676292 705472
rect 666277 705467 666343 705470
rect 669221 705122 669287 705125
rect 669221 705120 676292 705122
rect 669221 705064 669226 705120
rect 669282 705064 676292 705120
rect 669221 705062 676292 705064
rect 669221 705059 669287 705062
rect 42057 703490 42123 703493
rect 43161 703490 43227 703493
rect 42057 703488 43227 703490
rect 42057 703432 42062 703488
rect 42118 703432 43166 703488
rect 43222 703432 43227 703488
rect 42057 703430 43227 703432
rect 42057 703427 42123 703430
rect 43161 703427 43227 703430
rect 42057 702810 42123 702813
rect 42701 702810 42767 702813
rect 42057 702808 42767 702810
rect 42057 702752 42062 702808
rect 42118 702752 42706 702808
rect 42762 702752 42767 702808
rect 42057 702750 42767 702752
rect 42057 702747 42123 702750
rect 42701 702747 42767 702750
rect 41638 702340 41644 702404
rect 41708 702402 41714 702404
rect 42609 702402 42675 702405
rect 41708 702400 42675 702402
rect 41708 702344 42614 702400
rect 42670 702344 42675 702400
rect 41708 702342 42675 702344
rect 41708 702340 41714 702342
rect 42609 702339 42675 702342
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 42149 699956 42215 699957
rect 42149 699954 42196 699956
rect 42104 699952 42196 699954
rect 42104 699896 42154 699952
rect 42104 699894 42196 699896
rect 42149 699892 42196 699894
rect 42260 699892 42266 699956
rect 42149 699891 42215 699892
rect 670601 699818 670667 699821
rect 674925 699818 674991 699821
rect 670601 699816 674991 699818
rect 670601 699760 670606 699816
rect 670662 699760 674930 699816
rect 674986 699760 674991 699816
rect 670601 699758 674991 699760
rect 670601 699755 670667 699758
rect 674925 699755 674991 699758
rect 673177 698322 673243 698325
rect 675109 698322 675175 698325
rect 673177 698320 675175 698322
rect 673177 698264 673182 698320
rect 673238 698264 675114 698320
rect 675170 698264 675175 698320
rect 673177 698262 675175 698264
rect 673177 698259 673243 698262
rect 675109 698259 675175 698262
rect 41689 697914 41755 697917
rect 62757 697914 62823 697917
rect 41689 697912 62823 697914
rect 41689 697856 41694 697912
rect 41750 697856 62762 697912
rect 62818 697856 62823 697912
rect 41689 697854 62823 697856
rect 41689 697851 41755 697854
rect 62757 697851 62823 697854
rect 652385 696962 652451 696965
rect 650164 696960 652451 696962
rect 650164 696904 652390 696960
rect 652446 696904 652451 696960
rect 650164 696902 652451 696904
rect 652385 696899 652451 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 669589 695194 669655 695197
rect 675109 695194 675175 695197
rect 669589 695192 675175 695194
rect 669589 695136 669594 695192
rect 669650 695136 675114 695192
rect 675170 695136 675175 695192
rect 669589 695134 675175 695136
rect 669589 695131 669655 695134
rect 675109 695131 675175 695134
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676990 694106 676996 694108
rect 675894 694046 676996 694106
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 674005 693562 674071 693565
rect 675109 693562 675175 693565
rect 674005 693560 675175 693562
rect 674005 693504 674010 693560
rect 674066 693504 675114 693560
rect 675170 693504 675175 693560
rect 674005 693502 675175 693504
rect 674005 693499 674071 693502
rect 675109 693499 675175 693502
rect 668393 692882 668459 692885
rect 675109 692882 675175 692885
rect 668393 692880 675175 692882
rect 668393 692824 668398 692880
rect 668454 692824 675114 692880
rect 675170 692824 675175 692880
rect 668393 692822 675175 692824
rect 668393 692819 668459 692822
rect 675109 692819 675175 692822
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 674189 690162 674255 690165
rect 675385 690162 675451 690165
rect 674189 690160 675451 690162
rect 674189 690104 674194 690160
rect 674250 690104 675390 690160
rect 675446 690104 675451 690160
rect 674189 690102 675451 690104
rect 674189 690099 674255 690102
rect 675385 690099 675451 690102
rect 673545 689618 673611 689621
rect 675293 689618 675359 689621
rect 673545 689616 675359 689618
rect 673545 689560 673550 689616
rect 673606 689560 675298 689616
rect 675354 689560 675359 689616
rect 673545 689558 675359 689560
rect 673545 689555 673611 689558
rect 675293 689555 675359 689558
rect 663057 689346 663123 689349
rect 663057 689344 675172 689346
rect 663057 689288 663062 689344
rect 663118 689288 675172 689344
rect 663057 689286 675172 689288
rect 663057 689283 663123 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 667749 688938 667815 688941
rect 674925 688938 674991 688941
rect 667749 688936 674991 688938
rect 667749 688880 667754 688936
rect 667810 688880 674930 688936
rect 674986 688880 674991 688936
rect 667749 688878 674991 688880
rect 675112 688938 675172 689286
rect 675293 688938 675359 688941
rect 675112 688936 675359 688938
rect 675112 688880 675298 688936
rect 675354 688880 675359 688936
rect 675112 688878 675359 688880
rect 667749 688875 667815 688878
rect 674925 688875 674991 688878
rect 675293 688875 675359 688878
rect 671981 688666 672047 688669
rect 675109 688666 675175 688669
rect 671981 688664 675175 688666
rect 671981 688608 671986 688664
rect 672042 688608 675114 688664
rect 675170 688608 675175 688664
rect 671981 688606 675175 688608
rect 671981 688603 672047 688606
rect 675109 688603 675175 688606
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 670325 687442 670391 687445
rect 675477 687442 675543 687445
rect 670325 687440 675543 687442
rect 670325 687384 670330 687440
rect 670386 687384 675482 687440
rect 675538 687384 675543 687440
rect 670325 687382 675543 687384
rect 670325 687379 670391 687382
rect 675477 687379 675543 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 44357 686898 44423 686901
rect 41492 686896 44423 686898
rect 41492 686840 44362 686896
rect 44418 686840 44423 686896
rect 41492 686838 44423 686840
rect 44357 686835 44423 686838
rect 44357 686490 44423 686493
rect 41492 686488 44423 686490
rect 41492 686432 44362 686488
rect 44418 686432 44423 686488
rect 41492 686430 44423 686432
rect 44357 686427 44423 686430
rect 674833 686490 674899 686493
rect 675334 686490 675340 686492
rect 674833 686488 675340 686490
rect 674833 686432 674838 686488
rect 674894 686432 675340 686488
rect 674833 686430 675340 686432
rect 674833 686427 674899 686430
rect 675334 686428 675340 686430
rect 675404 686428 675410 686492
rect 44541 686082 44607 686085
rect 41492 686080 44607 686082
rect 41492 686024 44546 686080
rect 44602 686024 44607 686080
rect 41492 686022 44607 686024
rect 44541 686019 44607 686022
rect 672993 685810 673059 685813
rect 675477 685810 675543 685813
rect 672993 685808 675543 685810
rect 672993 685752 672998 685808
rect 673054 685752 675482 685808
rect 675538 685752 675543 685808
rect 672993 685750 675543 685752
rect 672993 685747 673059 685750
rect 675477 685747 675543 685750
rect 45369 685674 45435 685677
rect 41492 685672 45435 685674
rect 41492 685616 45374 685672
rect 45430 685616 45435 685672
rect 41492 685614 45435 685616
rect 45369 685611 45435 685614
rect 670969 685538 671035 685541
rect 675201 685538 675267 685541
rect 670969 685536 675267 685538
rect 670969 685480 670974 685536
rect 671030 685480 675206 685536
rect 675262 685480 675267 685536
rect 670969 685478 675267 685480
rect 670969 685475 671035 685478
rect 675201 685475 675267 685478
rect 44909 685266 44975 685269
rect 41492 685264 44975 685266
rect 41492 685208 44914 685264
rect 44970 685208 44975 685264
rect 41492 685206 44975 685208
rect 44909 685203 44975 685206
rect 45277 684858 45343 684861
rect 41492 684856 45343 684858
rect 41492 684800 45282 684856
rect 45338 684800 45343 684856
rect 41492 684798 45343 684800
rect 45277 684795 45343 684798
rect 45093 684450 45159 684453
rect 41492 684448 45159 684450
rect 41492 684392 45098 684448
rect 45154 684392 45159 684448
rect 41492 684390 45159 684392
rect 45093 684387 45159 684390
rect 44909 684042 44975 684045
rect 41492 684040 44975 684042
rect 41492 683984 44914 684040
rect 44970 683984 44975 684040
rect 41492 683982 44975 683984
rect 44909 683979 44975 683982
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 652017 683634 652083 683637
rect 650164 683632 652083 683634
rect 650164 683576 652022 683632
rect 652078 683576 652083 683632
rect 650164 683574 652083 683576
rect 652017 683571 652083 683574
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35433 682818 35499 682821
rect 35420 682816 35499 682818
rect 35420 682760 35438 682816
rect 35494 682760 35499 682816
rect 35420 682758 35499 682760
rect 35433 682755 35499 682758
rect 674414 682620 674420 682684
rect 674484 682682 674490 682684
rect 683205 682682 683271 682685
rect 674484 682680 683271 682682
rect 674484 682624 683210 682680
rect 683266 682624 683271 682680
rect 674484 682622 683271 682624
rect 674484 682620 674490 682622
rect 683205 682619 683271 682622
rect 35617 682410 35683 682413
rect 35604 682408 35683 682410
rect 35604 682352 35622 682408
rect 35678 682352 35683 682408
rect 35604 682350 35683 682352
rect 35617 682347 35683 682350
rect 674230 682348 674236 682412
rect 674300 682410 674306 682412
rect 683665 682410 683731 682413
rect 674300 682408 683731 682410
rect 674300 682352 683670 682408
rect 683726 682352 683731 682408
rect 674300 682350 683731 682352
rect 674300 682348 674306 682350
rect 683665 682347 683731 682350
rect 35801 682002 35867 682005
rect 35788 682000 35867 682002
rect 35788 681944 35806 682000
rect 35862 681944 35867 682000
rect 35788 681942 35867 681944
rect 35801 681939 35867 681942
rect 35617 681594 35683 681597
rect 35604 681592 35683 681594
rect 35604 681536 35622 681592
rect 35678 681536 35683 681592
rect 35604 681534 35683 681536
rect 35617 681531 35683 681534
rect 35801 681186 35867 681189
rect 35788 681184 35867 681186
rect 35788 681128 35806 681184
rect 35862 681128 35867 681184
rect 35788 681126 35867 681128
rect 35801 681123 35867 681126
rect 41781 681052 41847 681053
rect 41781 681050 41828 681052
rect 41736 681048 41828 681050
rect 41736 680992 41786 681048
rect 41736 680990 41828 680992
rect 41781 680988 41828 680990
rect 41892 680988 41898 681052
rect 673729 681050 673795 681053
rect 683481 681050 683547 681053
rect 673729 681048 683547 681050
rect 673729 680992 673734 681048
rect 673790 680992 683486 681048
rect 683542 680992 683547 681048
rect 673729 680990 683547 680992
rect 41781 680987 41847 680988
rect 673729 680987 673795 680990
rect 683481 680987 683547 680990
rect 35157 680778 35223 680781
rect 35157 680776 35236 680778
rect 35157 680720 35162 680776
rect 35218 680720 35236 680776
rect 35157 680718 35236 680720
rect 35157 680715 35223 680718
rect 44173 680370 44239 680373
rect 41492 680368 44239 680370
rect 41492 680312 44178 680368
rect 44234 680312 44239 680368
rect 41492 680310 44239 680312
rect 44173 680307 44239 680310
rect 42793 679962 42859 679965
rect 41492 679960 42859 679962
rect 41492 679904 42798 679960
rect 42854 679904 42859 679960
rect 41492 679902 42859 679904
rect 42793 679899 42859 679902
rect 44357 679554 44423 679557
rect 41492 679552 44423 679554
rect 41492 679496 44362 679552
rect 44418 679496 44423 679552
rect 41492 679494 44423 679496
rect 44357 679491 44423 679494
rect 43161 679146 43227 679149
rect 41492 679144 43227 679146
rect 41492 679088 43166 679144
rect 43222 679088 43227 679144
rect 41492 679086 43227 679088
rect 43161 679083 43227 679086
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678990 40794 678992
rect 40788 678930 41844 678990
rect 40788 678928 40794 678930
rect 40542 678708 40602 678928
rect 41784 678330 41844 678930
rect 41492 678270 41844 678330
rect 47209 677922 47275 677925
rect 41492 677920 47275 677922
rect 41492 677864 47214 677920
rect 47270 677864 47275 677920
rect 41492 677862 47275 677864
rect 47209 677859 47275 677862
rect 39990 677109 40050 677484
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 45737 676698 45803 676701
rect 41492 676696 45803 676698
rect 41492 676640 45742 676696
rect 45798 676640 45803 676696
rect 41492 676638 45803 676640
rect 45737 676635 45803 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 42057 673162 42123 673165
rect 42558 673162 42564 673164
rect 42057 673160 42564 673162
rect 42057 673104 42062 673160
rect 42118 673104 42564 673160
rect 42057 673102 42564 673104
rect 42057 673099 42123 673102
rect 42558 673100 42564 673102
rect 42628 673100 42634 673164
rect 669957 673162 670023 673165
rect 676489 673162 676555 673165
rect 669957 673160 676555 673162
rect 669957 673104 669962 673160
rect 670018 673104 676494 673160
rect 676550 673104 676555 673160
rect 669957 673102 676555 673104
rect 669957 673099 670023 673102
rect 676489 673099 676555 673102
rect 42374 672828 42380 672892
rect 42444 672890 42450 672892
rect 42793 672890 42859 672893
rect 42444 672888 42859 672890
rect 42444 672832 42798 672888
rect 42854 672832 42859 672888
rect 42444 672830 42859 672832
rect 42444 672828 42450 672830
rect 42793 672827 42859 672830
rect 40493 672618 40559 672621
rect 42793 672618 42859 672621
rect 40493 672616 42859 672618
rect 40493 672560 40498 672616
rect 40554 672560 42798 672616
rect 42854 672560 42859 672616
rect 40493 672558 42859 672560
rect 40493 672555 40559 672558
rect 42793 672555 42859 672558
rect 41505 672346 41571 672349
rect 42241 672346 42307 672349
rect 41505 672344 42307 672346
rect 41505 672288 41510 672344
rect 41566 672288 42246 672344
rect 42302 672288 42307 672344
rect 41505 672286 42307 672288
rect 41505 672283 41571 672286
rect 42241 672283 42307 672286
rect 37917 671258 37983 671261
rect 41822 671258 41828 671260
rect 37917 671256 41828 671258
rect 37917 671200 37922 671256
rect 37978 671200 41828 671256
rect 37917 671198 41828 671200
rect 37917 671195 37983 671198
rect 41822 671196 41828 671198
rect 41892 671196 41898 671260
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 676489 671122 676555 671125
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 676446 671120 676555 671122
rect 676446 671064 676494 671120
rect 676550 671064 676555 671120
rect 667197 671059 667263 671062
rect 676446 671059 676555 671064
rect 676446 670956 676506 671059
rect 668577 670578 668643 670581
rect 668577 670576 676292 670578
rect 668577 670520 668582 670576
rect 668638 670520 676292 670576
rect 668577 670518 676292 670520
rect 668577 670515 668643 670518
rect 651465 670442 651531 670445
rect 650164 670440 651531 670442
rect 650164 670384 651470 670440
rect 651526 670384 651531 670440
rect 650164 670382 651531 670384
rect 651465 670379 651531 670382
rect 672441 670170 672507 670173
rect 674598 670170 674604 670172
rect 672441 670168 674604 670170
rect 672441 670112 672446 670168
rect 672502 670112 674604 670168
rect 672441 670110 674604 670112
rect 672441 670107 672507 670110
rect 674598 670108 674604 670110
rect 674668 670108 674674 670172
rect 674833 670170 674899 670173
rect 674833 670168 676292 670170
rect 674833 670112 674838 670168
rect 674894 670112 676292 670168
rect 674833 670110 676292 670112
rect 674833 670107 674899 670110
rect 672441 669898 672507 669901
rect 672441 669896 676322 669898
rect 672441 669840 672446 669896
rect 672502 669840 676322 669896
rect 672441 669838 676322 669840
rect 672441 669835 672507 669838
rect 676262 669732 676322 669838
rect 672809 669490 672875 669493
rect 674833 669490 674899 669493
rect 672809 669488 674899 669490
rect 672809 669432 672814 669488
rect 672870 669432 674838 669488
rect 674894 669432 674899 669488
rect 672809 669430 674899 669432
rect 672809 669427 672875 669430
rect 674833 669427 674899 669430
rect 42190 669292 42196 669356
rect 42260 669354 42266 669356
rect 48957 669354 49023 669357
rect 42260 669352 49023 669354
rect 42260 669296 48962 669352
rect 49018 669296 49023 669352
rect 42260 669294 49023 669296
rect 42260 669292 42266 669294
rect 48957 669291 49023 669294
rect 674966 669292 674972 669356
rect 675036 669354 675042 669356
rect 675036 669294 676292 669354
rect 675036 669292 675042 669294
rect 672809 668946 672875 668949
rect 672809 668944 676292 668946
rect 672809 668888 672814 668944
rect 672870 668888 676292 668944
rect 672809 668886 676292 668888
rect 672809 668883 672875 668886
rect 42057 668538 42123 668541
rect 42558 668538 42564 668540
rect 42057 668536 42564 668538
rect 42057 668480 42062 668536
rect 42118 668480 42564 668536
rect 42057 668478 42564 668480
rect 42057 668475 42123 668478
rect 42558 668476 42564 668478
rect 42628 668476 42634 668540
rect 671613 668538 671679 668541
rect 671613 668536 676292 668538
rect 671613 668480 671618 668536
rect 671674 668480 676292 668536
rect 671613 668478 676292 668480
rect 671613 668475 671679 668478
rect 40718 668204 40724 668268
rect 40788 668266 40794 668268
rect 42241 668266 42307 668269
rect 40788 668264 42307 668266
rect 40788 668208 42246 668264
rect 42302 668208 42307 668264
rect 40788 668206 42307 668208
rect 40788 668204 40794 668206
rect 42241 668203 42307 668206
rect 671797 668130 671863 668133
rect 671797 668128 676292 668130
rect 671797 668072 671802 668128
rect 671858 668072 676292 668128
rect 671797 668070 676292 668072
rect 671797 668067 671863 668070
rect 41965 667724 42031 667725
rect 41965 667722 42012 667724
rect 41920 667720 42012 667722
rect 41920 667664 41970 667720
rect 41920 667662 42012 667664
rect 41965 667660 42012 667662
rect 42076 667660 42082 667724
rect 670785 667722 670851 667725
rect 670785 667720 676292 667722
rect 670785 667664 670790 667720
rect 670846 667664 676292 667720
rect 670785 667662 676292 667664
rect 41965 667659 42031 667660
rect 670785 667659 670851 667662
rect 671521 667314 671587 667317
rect 671521 667312 676292 667314
rect 671521 667256 671526 667312
rect 671582 667256 676292 667312
rect 671521 667254 676292 667256
rect 671521 667251 671587 667254
rect 683665 667042 683731 667045
rect 683622 667040 683731 667042
rect 683622 666984 683670 667040
rect 683726 666984 683731 667040
rect 683622 666979 683731 666984
rect 683622 666876 683682 666979
rect 42057 666634 42123 666637
rect 42374 666634 42380 666636
rect 42057 666632 42380 666634
rect 42057 666576 42062 666632
rect 42118 666576 42380 666632
rect 42057 666574 42380 666576
rect 42057 666571 42123 666574
rect 42374 666572 42380 666574
rect 42444 666572 42450 666636
rect 673361 666498 673427 666501
rect 673361 666496 676292 666498
rect 673361 666440 673366 666496
rect 673422 666440 676292 666496
rect 673361 666438 676292 666440
rect 673361 666435 673427 666438
rect 669773 666226 669839 666229
rect 676489 666226 676555 666229
rect 669773 666224 676555 666226
rect 669773 666168 669778 666224
rect 669834 666168 676494 666224
rect 676550 666168 676555 666224
rect 669773 666166 676555 666168
rect 669773 666163 669839 666166
rect 676489 666163 676555 666166
rect 667565 665954 667631 665957
rect 676262 665954 676322 666060
rect 667565 665952 676322 665954
rect 667565 665896 667570 665952
rect 667626 665896 676322 665952
rect 667565 665894 676322 665896
rect 667565 665891 667631 665894
rect 666461 665410 666527 665413
rect 676262 665410 676322 665652
rect 676489 665410 676555 665413
rect 666461 665408 676322 665410
rect 666461 665352 666466 665408
rect 666522 665352 676322 665408
rect 666461 665350 676322 665352
rect 676446 665408 676555 665410
rect 676446 665352 676494 665408
rect 676550 665352 676555 665408
rect 666461 665347 666527 665350
rect 676446 665347 676555 665352
rect 676446 665244 676506 665347
rect 42241 664866 42307 664869
rect 44357 664866 44423 664869
rect 42241 664864 44423 664866
rect 42241 664808 42246 664864
rect 42302 664808 44362 664864
rect 44418 664808 44423 664864
rect 42241 664806 44423 664808
rect 42241 664803 42307 664806
rect 44357 664803 44423 664806
rect 668761 664594 668827 664597
rect 676262 664594 676322 664836
rect 668761 664592 676322 664594
rect 668761 664536 668766 664592
rect 668822 664536 676322 664592
rect 668761 664534 676322 664536
rect 683205 664594 683271 664597
rect 683205 664592 683314 664594
rect 683205 664536 683210 664592
rect 683266 664536 683314 664592
rect 668761 664531 668827 664534
rect 683205 664531 683314 664536
rect 683254 664428 683314 664531
rect 40534 663988 40540 664052
rect 40604 664050 40610 664052
rect 41781 664050 41847 664053
rect 40604 664048 41847 664050
rect 40604 663992 41786 664048
rect 41842 663992 41847 664048
rect 40604 663990 41847 663992
rect 40604 663988 40610 663990
rect 41781 663987 41847 663990
rect 674414 663988 674420 664052
rect 674484 664050 674490 664052
rect 674484 663990 676292 664050
rect 674484 663988 674490 663990
rect 669405 663642 669471 663645
rect 669405 663640 676292 663642
rect 669405 663584 669410 663640
rect 669466 663584 676292 663640
rect 669405 663582 676292 663584
rect 669405 663579 669471 663582
rect 42425 663506 42491 663509
rect 44173 663506 44239 663509
rect 42425 663504 44239 663506
rect 42425 663448 42430 663504
rect 42486 663448 44178 663504
rect 44234 663448 44239 663504
rect 42425 663446 44239 663448
rect 42425 663443 42491 663446
rect 44173 663443 44239 663446
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 676262 662962 676322 663204
rect 683481 662962 683547 662965
rect 669270 662902 676322 662962
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 42241 662690 42307 662693
rect 43161 662690 43227 662693
rect 42241 662688 43227 662690
rect 42241 662632 42246 662688
rect 42302 662632 43166 662688
rect 43222 662632 43227 662688
rect 42241 662630 43227 662632
rect 42241 662627 42307 662630
rect 43161 662627 43227 662630
rect 668209 662554 668275 662557
rect 669270 662554 669330 662902
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 668209 662552 669330 662554
rect 668209 662496 668214 662552
rect 668270 662496 669330 662552
rect 668209 662494 669330 662496
rect 668209 662491 668275 662494
rect 671153 662416 671219 662421
rect 671153 662360 671158 662416
rect 671214 662360 671219 662416
rect 671153 662355 671219 662360
rect 672625 662418 672691 662421
rect 672625 662416 676292 662418
rect 672625 662360 672630 662416
rect 672686 662360 676292 662416
rect 672625 662358 676292 662360
rect 672625 662355 672691 662358
rect 671156 662146 671216 662355
rect 671156 662086 676322 662146
rect 676262 661980 676322 662086
rect 672165 661602 672231 661605
rect 672165 661600 676292 661602
rect 672165 661544 672170 661600
rect 672226 661544 676292 661600
rect 672165 661542 676292 661544
rect 672165 661539 672231 661542
rect 672625 661194 672691 661197
rect 672625 661192 676292 661194
rect 672625 661136 672630 661192
rect 672686 661136 676292 661192
rect 672625 661134 676292 661136
rect 672625 661131 672691 661134
rect 673361 660786 673427 660789
rect 673361 660784 676292 660786
rect 673361 660728 673366 660784
rect 673422 660756 676292 660784
rect 673422 660728 676322 660756
rect 673361 660726 676322 660728
rect 673361 660723 673427 660726
rect 676262 660348 676322 660726
rect 673361 659970 673427 659973
rect 673361 659968 676292 659970
rect 673361 659912 673366 659968
rect 673422 659912 676292 659968
rect 673361 659910 676292 659912
rect 673361 659907 673427 659910
rect 41454 659636 41460 659700
rect 41524 659698 41530 659700
rect 42609 659698 42675 659701
rect 41524 659696 42675 659698
rect 41524 659640 42614 659696
rect 42670 659640 42675 659696
rect 41524 659638 42675 659640
rect 41524 659636 41530 659638
rect 42609 659635 42675 659638
rect 42057 659154 42123 659157
rect 42793 659154 42859 659157
rect 42057 659152 42859 659154
rect 42057 659096 42062 659152
rect 42118 659096 42798 659152
rect 42854 659096 42859 659152
rect 42057 659094 42859 659096
rect 42057 659091 42123 659094
rect 42793 659091 42859 659094
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42425 658610 42491 658613
rect 41708 658608 42491 658610
rect 41708 658552 42430 658608
rect 42486 658552 42491 658608
rect 41708 658550 42491 658552
rect 41708 658548 41714 658550
rect 42425 658547 42491 658550
rect 41822 658276 41828 658340
rect 41892 658338 41898 658340
rect 42241 658338 42307 658341
rect 41892 658336 42307 658338
rect 41892 658280 42246 658336
rect 42302 658280 42307 658336
rect 41892 658278 42307 658280
rect 41892 658276 41898 658278
rect 42241 658275 42307 658278
rect 42057 657386 42123 657389
rect 42609 657386 42675 657389
rect 42057 657384 42675 657386
rect 42057 657328 42062 657384
rect 42118 657328 42614 657384
rect 42670 657328 42675 657384
rect 42057 657326 42675 657328
rect 42057 657323 42123 657326
rect 42609 657323 42675 657326
rect 651465 657114 651531 657117
rect 650164 657112 651531 657114
rect 650164 657056 651470 657112
rect 651526 657056 651531 657112
rect 650164 657054 651531 657056
rect 651465 657051 651531 657054
rect 668209 654258 668275 654261
rect 675385 654258 675451 654261
rect 668209 654256 675451 654258
rect 668209 654200 668214 654256
rect 668270 654200 675390 654256
rect 675446 654200 675451 654256
rect 668209 654198 675451 654200
rect 668209 654195 668275 654198
rect 675385 654195 675451 654198
rect 44214 653108 44220 653172
rect 44284 653170 44290 653172
rect 44725 653170 44791 653173
rect 44284 653168 44791 653170
rect 44284 653112 44730 653168
rect 44786 653112 44791 653168
rect 44284 653110 44791 653112
rect 44284 653108 44290 653110
rect 44725 653107 44791 653110
rect 675334 652836 675340 652900
rect 675404 652898 675410 652900
rect 675569 652898 675635 652901
rect 675404 652896 675635 652898
rect 675404 652840 675574 652896
rect 675630 652840 675635 652896
rect 675404 652838 675635 652840
rect 675404 652836 675410 652838
rect 675569 652835 675635 652838
rect 674966 651476 674972 651540
rect 675036 651538 675042 651540
rect 675385 651538 675451 651541
rect 675036 651536 675451 651538
rect 675036 651480 675390 651536
rect 675446 651480 675451 651536
rect 675036 651478 675451 651480
rect 675036 651476 675042 651478
rect 675385 651475 675451 651478
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 675201 649772 675267 649773
rect 675150 649770 675156 649772
rect 675110 649710 675156 649770
rect 675220 649768 675267 649772
rect 675262 649712 675267 649768
rect 675150 649708 675156 649710
rect 675220 649708 675267 649712
rect 675201 649707 675267 649708
rect 674414 648892 674420 648956
rect 674484 648954 674490 648956
rect 675385 648954 675451 648957
rect 674484 648952 675451 648954
rect 674484 648896 675390 648952
rect 675446 648896 675451 648952
rect 674484 648894 675451 648896
rect 674484 648892 674490 648894
rect 675385 648891 675451 648894
rect 669037 648682 669103 648685
rect 675477 648682 675543 648685
rect 669037 648680 675543 648682
rect 669037 648624 669042 648680
rect 669098 648624 675482 648680
rect 675538 648624 675543 648680
rect 669037 648622 675543 648624
rect 669037 648619 669103 648622
rect 675477 648619 675543 648622
rect 673729 647866 673795 647869
rect 675477 647866 675543 647869
rect 673729 647864 675543 647866
rect 673729 647808 673734 647864
rect 673790 647808 675482 647864
rect 675538 647808 675543 647864
rect 673729 647806 675543 647808
rect 673729 647803 673795 647806
rect 675477 647803 675543 647806
rect 674465 647596 674531 647597
rect 674414 647532 674420 647596
rect 674484 647594 674531 647596
rect 674833 647594 674899 647597
rect 675150 647594 675156 647596
rect 674484 647592 674576 647594
rect 674526 647536 674576 647592
rect 674484 647534 674576 647536
rect 674833 647592 675156 647594
rect 674833 647536 674838 647592
rect 674894 647536 675156 647592
rect 674833 647534 675156 647536
rect 674484 647532 674531 647534
rect 674465 647531 674531 647532
rect 674833 647531 674899 647534
rect 675150 647532 675156 647534
rect 675220 647532 675226 647596
rect 675017 647324 675083 647325
rect 674966 647260 674972 647324
rect 675036 647322 675083 647324
rect 675036 647320 675128 647322
rect 675078 647264 675128 647320
rect 675036 647262 675128 647264
rect 675036 647260 675083 647262
rect 675017 647259 675083 647260
rect 35801 646778 35867 646781
rect 35801 646776 35910 646778
rect 35801 646720 35806 646776
rect 35862 646720 35910 646776
rect 35801 646715 35910 646720
rect 35850 646642 35910 646715
rect 51717 646642 51783 646645
rect 35850 646640 51783 646642
rect 35850 646584 51722 646640
rect 51778 646584 51783 646640
rect 35850 646582 51783 646584
rect 51717 646579 51783 646582
rect 669773 645418 669839 645421
rect 675477 645418 675543 645421
rect 669773 645416 675543 645418
rect 669773 645360 669778 645416
rect 669834 645360 675482 645416
rect 675538 645360 675543 645416
rect 669773 645358 675543 645360
rect 669773 645355 669839 645358
rect 675477 645355 675543 645358
rect 674046 645084 674052 645148
rect 674116 645146 674122 645148
rect 674373 645146 674439 645149
rect 674116 645144 674439 645146
rect 674116 645088 674378 645144
rect 674434 645088 674439 645144
rect 674116 645086 674439 645088
rect 674116 645084 674122 645086
rect 674373 645083 674439 645086
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 669957 644874 670023 644877
rect 675385 644874 675451 644877
rect 669957 644872 675451 644874
rect 669957 644816 669962 644872
rect 670018 644816 675390 644872
rect 675446 644816 675451 644872
rect 669957 644814 675451 644816
rect 669957 644811 670023 644814
rect 675385 644811 675451 644814
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 35758 644504 35818 644675
rect 675753 644330 675819 644333
rect 676806 644330 676812 644332
rect 675753 644328 676812 644330
rect 675753 644272 675758 644328
rect 675814 644272 676812 644328
rect 675753 644270 676812 644272
rect 675753 644267 675819 644270
rect 676806 644268 676812 644270
rect 676876 644268 676882 644332
rect 41462 643922 41522 644096
rect 675201 644060 675267 644061
rect 675150 643996 675156 644060
rect 675220 644058 675267 644060
rect 675220 644056 675312 644058
rect 675262 644000 675312 644056
rect 675220 643998 675312 644000
rect 675220 643996 675267 643998
rect 675201 643995 675267 643996
rect 41462 643862 45570 643922
rect 41462 643650 41522 643688
rect 44541 643650 44607 643653
rect 41462 643648 44607 643650
rect 41462 643592 44546 643648
rect 44602 643592 44607 643648
rect 41462 643590 44607 643592
rect 44541 643587 44607 643590
rect 44725 643378 44791 643381
rect 41462 643376 44791 643378
rect 41462 643320 44730 643376
rect 44786 643320 44791 643376
rect 41462 643318 44791 643320
rect 41462 643280 41522 643318
rect 44725 643315 44791 643318
rect 45510 643242 45570 643862
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 661861 643786 661927 643789
rect 675201 643786 675267 643789
rect 661861 643784 675267 643786
rect 661861 643728 661866 643784
rect 661922 643728 675206 643784
rect 675262 643728 675267 643784
rect 661861 643726 675267 643728
rect 661861 643723 661927 643726
rect 675201 643723 675267 643726
rect 671470 643452 671476 643516
rect 671540 643514 671546 643516
rect 675477 643514 675543 643517
rect 671540 643512 675543 643514
rect 671540 643456 675482 643512
rect 675538 643456 675543 643512
rect 671540 643454 675543 643456
rect 671540 643452 671546 643454
rect 675477 643451 675543 643454
rect 55857 643242 55923 643245
rect 45510 643240 55923 643242
rect 45510 643184 55862 643240
rect 55918 643184 55923 643240
rect 45510 643182 55923 643184
rect 55857 643179 55923 643182
rect 45369 643106 45435 643109
rect 41462 643104 45435 643106
rect 41462 643048 45374 643104
rect 45430 643048 45435 643104
rect 41462 643046 45435 643048
rect 41462 642872 41522 643046
rect 45369 643043 45435 643046
rect 44449 642562 44515 642565
rect 41462 642560 44515 642562
rect 41462 642504 44454 642560
rect 44510 642504 44515 642560
rect 41462 642502 44515 642504
rect 41462 642464 41522 642502
rect 44449 642499 44515 642502
rect 45185 642290 45251 642293
rect 41462 642288 45251 642290
rect 41462 642232 45190 642288
rect 45246 642232 45251 642288
rect 41462 642230 45251 642232
rect 41462 642056 41522 642230
rect 45185 642227 45251 642230
rect 674189 641746 674255 641749
rect 675293 641746 675359 641749
rect 674189 641744 675359 641746
rect 674189 641688 674194 641744
rect 674250 641688 675298 641744
rect 675354 641688 675359 641744
rect 674189 641686 675359 641688
rect 674189 641683 674255 641686
rect 675293 641683 675359 641686
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 44909 641474 44975 641477
rect 41462 641472 44975 641474
rect 41462 641416 44914 641472
rect 44970 641416 44975 641472
rect 41462 641414 44975 641416
rect 41462 641240 41522 641414
rect 44909 641411 44975 641414
rect 41781 641202 41847 641205
rect 45001 641202 45067 641205
rect 41781 641200 45067 641202
rect 41781 641144 41786 641200
rect 41842 641144 45006 641200
rect 45062 641144 45067 641200
rect 41781 641142 45067 641144
rect 41781 641139 41847 641142
rect 45001 641139 45067 641142
rect 45369 640930 45435 640933
rect 41462 640928 45435 640930
rect 41462 640872 45374 640928
rect 45430 640872 45435 640928
rect 41462 640870 45435 640872
rect 41462 640832 41522 640870
rect 45369 640867 45435 640870
rect 674833 640794 674899 640797
rect 674833 640792 676230 640794
rect 674833 640736 674838 640792
rect 674894 640736 676230 640792
rect 674833 640734 676230 640736
rect 674833 640731 674899 640734
rect 41638 640658 41644 640660
rect 41462 640598 41644 640658
rect 41462 640424 41522 640598
rect 41638 640596 41644 640598
rect 41708 640596 41714 640660
rect 671153 640522 671219 640525
rect 675385 640522 675451 640525
rect 671153 640520 675451 640522
rect 671153 640464 671158 640520
rect 671214 640464 675390 640520
rect 675446 640464 675451 640520
rect 671153 640462 675451 640464
rect 671153 640459 671219 640462
rect 675385 640459 675451 640462
rect 676170 640250 676230 640734
rect 676622 640250 676628 640252
rect 676170 640190 676628 640250
rect 676622 640188 676628 640190
rect 676692 640188 676698 640252
rect 35758 639845 35818 640016
rect 35758 639840 35867 639845
rect 35758 639784 35806 639840
rect 35862 639784 35867 639840
rect 35758 639782 35867 639784
rect 35801 639779 35867 639782
rect 41462 639436 41522 639608
rect 41454 639372 41460 639436
rect 41524 639372 41530 639436
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35758 638621 35818 638792
rect 672165 638754 672231 638757
rect 675477 638754 675543 638757
rect 672165 638752 675543 638754
rect 672165 638696 672170 638752
rect 672226 638696 675482 638752
rect 675538 638696 675543 638752
rect 672165 638694 675543 638696
rect 672165 638691 672231 638694
rect 675477 638691 675543 638694
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 41781 638210 41847 638213
rect 47393 638210 47459 638213
rect 41781 638208 47459 638210
rect 41781 638152 41786 638208
rect 41842 638152 47398 638208
rect 47454 638152 47459 638208
rect 41781 638150 47459 638152
rect 32397 638147 32463 638150
rect 41781 638147 41847 638150
rect 47393 638147 47459 638150
rect 675150 638012 675156 638076
rect 675220 638074 675226 638076
rect 675385 638074 675451 638077
rect 675220 638072 675451 638074
rect 675220 638016 675390 638072
rect 675446 638016 675451 638072
rect 675220 638014 675451 638016
rect 675220 638012 675226 638014
rect 675385 638011 675451 638014
rect 41462 637802 41522 637976
rect 676622 637876 676628 637940
rect 676692 637938 676698 637940
rect 677501 637938 677567 637941
rect 676692 637936 677567 637938
rect 676692 637880 677506 637936
rect 677562 637880 677567 637936
rect 676692 637878 677567 637880
rect 676692 637876 676698 637878
rect 677501 637875 677567 637878
rect 46013 637802 46079 637805
rect 41462 637800 46079 637802
rect 41462 637744 46018 637800
rect 46074 637744 46079 637800
rect 41462 637742 46079 637744
rect 46013 637739 46079 637742
rect 675334 637604 675340 637668
rect 675404 637666 675410 637668
rect 675753 637666 675819 637669
rect 675404 637664 675819 637666
rect 675404 637608 675758 637664
rect 675814 637608 675819 637664
rect 675404 637606 675819 637608
rect 675404 637604 675410 637606
rect 675753 637603 675819 637606
rect 41781 637598 41847 637601
rect 41492 637596 41847 637598
rect 41492 637540 41786 637596
rect 41842 637540 41847 637596
rect 41492 637538 41847 637540
rect 41781 637535 41847 637538
rect 40033 637394 40099 637397
rect 41822 637394 41828 637396
rect 40033 637392 41828 637394
rect 40033 637336 40038 637392
rect 40094 637336 41828 637392
rect 40033 637334 41828 637336
rect 40033 637331 40099 637334
rect 41822 637332 41828 637334
rect 41892 637332 41898 637396
rect 41462 637122 41522 637160
rect 46197 637122 46263 637125
rect 41462 637120 46263 637122
rect 41462 637064 46202 637120
rect 46258 637064 46263 637120
rect 41462 637062 46263 637064
rect 46197 637059 46263 637062
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 673545 636850 673611 636853
rect 683297 636850 683363 636853
rect 673545 636848 683363 636850
rect 673545 636792 673550 636848
rect 673606 636792 683302 636848
rect 683358 636792 683363 636848
rect 673545 636790 683363 636792
rect 673545 636787 673611 636790
rect 683297 636787 683363 636790
rect 41462 636578 41522 636752
rect 45185 636578 45251 636581
rect 41462 636576 45251 636578
rect 41462 636520 45190 636576
rect 45246 636520 45251 636576
rect 41462 636518 45251 636520
rect 45185 636515 45251 636518
rect 41462 636306 41522 636344
rect 43161 636306 43227 636309
rect 41462 636304 43227 636306
rect 41462 636248 43166 636304
rect 43222 636248 43227 636304
rect 41462 636246 43227 636248
rect 43161 636243 43227 636246
rect 41462 635762 41522 635936
rect 44909 635762 44975 635765
rect 41462 635760 44975 635762
rect 41462 635704 44914 635760
rect 44970 635704 44975 635760
rect 41462 635702 44975 635704
rect 44909 635699 44975 635702
rect 41462 635354 41522 635528
rect 672809 635490 672875 635493
rect 683665 635490 683731 635493
rect 672809 635488 683731 635490
rect 672809 635432 672814 635488
rect 672870 635432 683670 635488
rect 683726 635432 683731 635488
rect 672809 635430 683731 635432
rect 672809 635427 672875 635430
rect 683665 635427 683731 635430
rect 43897 635354 43963 635357
rect 41462 635352 43963 635354
rect 41462 635296 43902 635352
rect 43958 635296 43963 635352
rect 41462 635294 43963 635296
rect 43897 635291 43963 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 40542 634540 40602 634712
rect 40534 634476 40540 634540
rect 40604 634476 40610 634540
rect 41462 633858 41522 634304
rect 42517 633858 42583 633861
rect 41462 633856 42583 633858
rect 41462 633800 42522 633856
rect 42578 633800 42583 633856
rect 41462 633798 42583 633800
rect 42517 633795 42583 633798
rect 41462 633450 41522 633488
rect 44265 633450 44331 633453
rect 41462 633448 44331 633450
rect 41462 633392 44270 633448
rect 44326 633392 44331 633448
rect 41462 633390 44331 633392
rect 44265 633387 44331 633390
rect 674925 631410 674991 631413
rect 675334 631410 675340 631412
rect 674925 631408 675340 631410
rect 674925 631352 674930 631408
rect 674986 631352 675340 631408
rect 674925 631350 675340 631352
rect 674925 631347 674991 631350
rect 675334 631348 675340 631350
rect 675404 631348 675410 631412
rect 675753 631410 675819 631413
rect 676070 631410 676076 631412
rect 675753 631408 676076 631410
rect 675753 631352 675758 631408
rect 675814 631352 676076 631408
rect 675753 631350 676076 631352
rect 675753 631347 675819 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 651465 630594 651531 630597
rect 650164 630592 651531 630594
rect 650164 630536 651470 630592
rect 651526 630536 651531 630592
rect 650164 630534 651531 630536
rect 651465 630531 651531 630534
rect 671337 627874 671403 627877
rect 675845 627874 675911 627877
rect 671337 627872 675911 627874
rect 671337 627816 671342 627872
rect 671398 627816 675850 627872
rect 675906 627816 675911 627872
rect 671337 627814 675911 627816
rect 671337 627811 671403 627814
rect 675845 627811 675911 627814
rect 41413 627738 41479 627741
rect 42701 627738 42767 627741
rect 41413 627736 42767 627738
rect 41413 627680 41418 627736
rect 41474 627680 42706 627736
rect 42762 627680 42767 627736
rect 41413 627678 42767 627680
rect 41413 627675 41479 627678
rect 42701 627675 42767 627678
rect 42558 626588 42564 626652
rect 42628 626650 42634 626652
rect 50337 626650 50403 626653
rect 42628 626648 50403 626650
rect 42628 626592 50342 626648
rect 50398 626592 50403 626648
rect 42628 626590 50403 626592
rect 42628 626588 42634 626590
rect 50337 626587 50403 626590
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 42057 625834 42123 625837
rect 42517 625834 42583 625837
rect 42057 625832 42583 625834
rect 42057 625776 42062 625832
rect 42118 625776 42522 625832
rect 42578 625776 42583 625832
rect 42057 625774 42583 625776
rect 42057 625771 42123 625774
rect 42517 625771 42583 625774
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 669270 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 42190 625228 42196 625292
rect 42260 625290 42266 625292
rect 45277 625290 45343 625293
rect 42260 625288 45343 625290
rect 42260 625232 45282 625288
rect 45338 625232 45343 625288
rect 42260 625230 45343 625232
rect 42260 625228 42266 625230
rect 45277 625227 45343 625230
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 672441 625154 672507 625157
rect 672441 625152 676292 625154
rect 672441 625096 672446 625152
rect 672502 625096 676292 625152
rect 672441 625094 676292 625096
rect 672441 625091 672507 625094
rect 42517 625020 42583 625021
rect 42517 625018 42564 625020
rect 42472 625016 42564 625018
rect 42472 624960 42522 625016
rect 42472 624958 42564 624960
rect 42517 624956 42564 624958
rect 42628 624956 42634 625020
rect 42517 624955 42583 624956
rect 674373 624882 674439 624885
rect 683113 624882 683179 624885
rect 674373 624880 683179 624882
rect 674373 624824 674378 624880
rect 674434 624824 683118 624880
rect 683174 624824 683179 624880
rect 674373 624822 683179 624824
rect 674373 624819 674439 624822
rect 683113 624819 683179 624822
rect 671613 624474 671679 624477
rect 676262 624474 676322 624716
rect 683665 624474 683731 624477
rect 671613 624472 676322 624474
rect 671613 624416 671618 624472
rect 671674 624416 676322 624472
rect 671613 624414 676322 624416
rect 683622 624472 683731 624474
rect 683622 624416 683670 624472
rect 683726 624416 683731 624472
rect 671613 624411 671679 624414
rect 683622 624411 683731 624416
rect 683622 624308 683682 624411
rect 42241 624066 42307 624069
rect 43161 624066 43227 624069
rect 42241 624064 43227 624066
rect 42241 624008 42246 624064
rect 42302 624008 43166 624064
rect 43222 624008 43227 624064
rect 42241 624006 43227 624008
rect 42241 624003 42307 624006
rect 43161 624003 43227 624006
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 670785 623930 670851 623933
rect 670785 623928 676292 623930
rect 670785 623872 670790 623928
rect 670846 623872 676292 623928
rect 670785 623870 676292 623872
rect 670785 623867 670851 623870
rect 671797 623522 671863 623525
rect 671797 623520 676292 623522
rect 671797 623464 671802 623520
rect 671858 623464 676292 623520
rect 671797 623462 676292 623464
rect 671797 623459 671863 623462
rect 41965 623386 42031 623389
rect 42190 623386 42196 623388
rect 41965 623384 42196 623386
rect 41965 623328 41970 623384
rect 42026 623328 42196 623384
rect 41965 623326 42196 623328
rect 41965 623323 42031 623326
rect 42190 623324 42196 623326
rect 42260 623324 42266 623388
rect 42425 623386 42491 623389
rect 43897 623386 43963 623389
rect 42425 623384 43963 623386
rect 42425 623328 42430 623384
rect 42486 623328 43902 623384
rect 43958 623328 43963 623384
rect 42425 623326 43963 623328
rect 42425 623323 42491 623326
rect 43897 623323 43963 623326
rect 671705 623114 671771 623117
rect 671705 623112 676292 623114
rect 671705 623056 671710 623112
rect 671766 623056 676292 623112
rect 671705 623054 676292 623056
rect 671705 623051 671771 623054
rect 671429 622706 671495 622709
rect 671429 622704 676292 622706
rect 671429 622648 671434 622704
rect 671490 622648 676292 622704
rect 671429 622646 676292 622648
rect 671429 622643 671495 622646
rect 672809 622298 672875 622301
rect 672809 622296 676292 622298
rect 672809 622240 672814 622296
rect 672870 622240 676292 622296
rect 672809 622238 676292 622240
rect 672809 622235 672875 622238
rect 40718 622100 40724 622164
rect 40788 622162 40794 622164
rect 41781 622162 41847 622165
rect 40788 622160 41847 622162
rect 40788 622104 41786 622160
rect 41842 622104 41847 622160
rect 40788 622102 41847 622104
rect 40788 622100 40794 622102
rect 41781 622099 41847 622102
rect 677501 622026 677567 622029
rect 677501 622024 677610 622026
rect 677501 621968 677506 622024
rect 677562 621968 677610 622024
rect 677501 621963 677610 621968
rect 677550 621860 677610 621963
rect 674606 621422 676292 621482
rect 667749 621210 667815 621213
rect 674606 621210 674666 621422
rect 667749 621208 674666 621210
rect 667749 621152 667754 621208
rect 667810 621152 674666 621208
rect 667749 621150 674666 621152
rect 667749 621147 667815 621150
rect 674790 621014 676292 621074
rect 673177 620938 673243 620941
rect 674790 620938 674850 621014
rect 673177 620936 674850 620938
rect 673177 620880 673182 620936
rect 673238 620880 674850 620936
rect 673177 620878 674850 620880
rect 673177 620875 673243 620878
rect 669589 620666 669655 620669
rect 669589 620664 676292 620666
rect 669589 620608 669594 620664
rect 669650 620608 676292 620664
rect 669589 620606 676292 620608
rect 669589 620603 669655 620606
rect 668393 620258 668459 620261
rect 668393 620256 676292 620258
rect 668393 620200 668398 620256
rect 668454 620200 676292 620256
rect 668393 620198 676292 620200
rect 668393 620195 668459 620198
rect 42517 620122 42583 620125
rect 44909 620122 44975 620125
rect 42517 620120 44975 620122
rect 42517 620064 42522 620120
rect 42578 620064 44914 620120
rect 44970 620064 44975 620120
rect 42517 620062 44975 620064
rect 42517 620059 42583 620062
rect 44909 620059 44975 620062
rect 40534 619788 40540 619852
rect 40604 619850 40610 619852
rect 42701 619850 42767 619853
rect 40604 619848 42767 619850
rect 40604 619792 42706 619848
rect 42762 619792 42767 619848
rect 40604 619790 42767 619792
rect 40604 619788 40610 619790
rect 42701 619787 42767 619790
rect 670969 619850 671035 619853
rect 670969 619848 676292 619850
rect 670969 619792 670974 619848
rect 671030 619792 676292 619848
rect 670969 619790 676292 619792
rect 670969 619787 671035 619790
rect 670417 619442 670483 619445
rect 670417 619440 676292 619442
rect 670417 619384 670422 619440
rect 670478 619384 676292 619440
rect 670417 619382 676292 619384
rect 670417 619379 670483 619382
rect 676990 619108 676996 619172
rect 677060 619108 677066 619172
rect 676998 619004 677058 619108
rect 42425 618898 42491 618901
rect 47393 618898 47459 618901
rect 42425 618896 47459 618898
rect 42425 618840 42430 618896
rect 42486 618840 47398 618896
rect 47454 618840 47459 618896
rect 42425 618838 47459 618840
rect 42425 618835 42491 618838
rect 47393 618835 47459 618838
rect 673913 618626 673979 618629
rect 673913 618624 676292 618626
rect 673913 618568 673918 618624
rect 673974 618568 676292 618624
rect 673913 618566 676292 618568
rect 673913 618563 673979 618566
rect 42425 618490 42491 618493
rect 46197 618490 46263 618493
rect 42425 618488 46263 618490
rect 42425 618432 42430 618488
rect 42486 618432 46202 618488
rect 46258 618432 46263 618488
rect 42425 618430 46263 618432
rect 42425 618427 42491 618430
rect 46197 618427 46263 618430
rect 670417 618218 670483 618221
rect 670417 618216 676292 618218
rect 670417 618160 670422 618216
rect 670478 618160 676292 618216
rect 670417 618158 676292 618160
rect 670417 618155 670483 618158
rect 683297 617946 683363 617949
rect 683254 617944 683363 617946
rect 683254 617888 683302 617944
rect 683358 617888 683363 617944
rect 683254 617883 683363 617888
rect 683254 617780 683314 617883
rect 674741 617402 674807 617405
rect 674741 617400 676292 617402
rect 674741 617344 674746 617400
rect 674802 617344 676292 617400
rect 674741 617342 676292 617344
rect 674741 617339 674807 617342
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683113 617130 683179 617133
rect 683070 617128 683179 617130
rect 683070 617072 683118 617128
rect 683174 617072 683179 617128
rect 683070 617067 683179 617072
rect 683070 616964 683130 617067
rect 672073 616722 672139 616725
rect 672073 616720 676230 616722
rect 672073 616664 672078 616720
rect 672134 616664 676230 616720
rect 672073 616662 676230 616664
rect 672073 616659 672139 616662
rect 676170 616586 676230 616662
rect 676170 616526 676292 616586
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 42057 615908 42123 615909
rect 42006 615906 42012 615908
rect 41966 615846 42012 615906
rect 42076 615904 42123 615908
rect 42118 615848 42123 615904
rect 42006 615844 42012 615846
rect 42076 615844 42123 615848
rect 42057 615843 42123 615844
rect 672993 615770 673059 615773
rect 672993 615768 676292 615770
rect 672993 615712 672998 615768
rect 673054 615740 676292 615768
rect 673054 615712 676322 615740
rect 672993 615710 676322 615712
rect 672993 615707 673059 615710
rect 46013 615634 46079 615637
rect 42704 615632 46079 615634
rect 42704 615576 46018 615632
rect 46074 615576 46079 615632
rect 42704 615574 46079 615576
rect 41454 615436 41460 615500
rect 41524 615498 41530 615500
rect 42425 615498 42491 615501
rect 41524 615496 42491 615498
rect 41524 615440 42430 615496
rect 42486 615440 42491 615496
rect 41524 615438 42491 615440
rect 41524 615436 41530 615438
rect 42425 615435 42491 615438
rect 42057 615226 42123 615229
rect 42704 615226 42764 615574
rect 46013 615571 46079 615574
rect 676262 615332 676322 615710
rect 42057 615224 42764 615226
rect 42057 615168 42062 615224
rect 42118 615168 42764 615224
rect 42057 615166 42764 615168
rect 42057 615163 42123 615166
rect 672073 614954 672139 614957
rect 672073 614952 676292 614954
rect 672073 614896 672078 614952
rect 672134 614896 676292 614952
rect 672073 614894 676292 614896
rect 672073 614891 672139 614894
rect 41873 614140 41939 614141
rect 41822 614138 41828 614140
rect 41782 614078 41828 614138
rect 41892 614136 41939 614140
rect 41934 614080 41939 614136
rect 41822 614076 41828 614078
rect 41892 614076 41939 614080
rect 41873 614075 41939 614076
rect 43989 614138 44055 614141
rect 44214 614138 44220 614140
rect 43989 614136 44220 614138
rect 43989 614080 43994 614136
rect 44050 614080 44220 614136
rect 43989 614078 44220 614080
rect 43989 614075 44055 614078
rect 44214 614076 44220 614078
rect 44284 614076 44290 614140
rect 42977 612370 43043 612373
rect 43575 612370 43641 612373
rect 42977 612368 43641 612370
rect 42977 612312 42982 612368
rect 43038 612312 43580 612368
rect 43636 612312 43641 612368
rect 42977 612310 43641 612312
rect 42977 612307 43043 612310
rect 43575 612307 43641 612310
rect 42701 611010 42767 611013
rect 44817 611010 44883 611013
rect 42701 611008 44883 611010
rect 42701 610952 42706 611008
rect 42762 610952 44822 611008
rect 44878 610952 44883 611008
rect 42701 610950 44883 610952
rect 42701 610947 42767 610950
rect 44817 610947 44883 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 675477 607748 675543 607749
rect 675477 607744 675524 607748
rect 675588 607746 675594 607748
rect 675477 607688 675482 607744
rect 675477 607684 675524 607688
rect 675588 607686 675634 607746
rect 675588 607684 675594 607686
rect 675477 607683 675543 607684
rect 670601 607338 670667 607341
rect 675477 607338 675543 607341
rect 670601 607336 675543 607338
rect 670601 607280 670606 607336
rect 670662 607280 675482 607336
rect 675538 607280 675543 607336
rect 670601 607278 675543 607280
rect 670601 607275 670667 607278
rect 675477 607275 675543 607278
rect 674373 606522 674439 606525
rect 675477 606522 675543 606525
rect 674373 606520 675543 606522
rect 674373 606464 674378 606520
rect 674434 606464 675482 606520
rect 675538 606464 675543 606520
rect 674373 606462 675543 606464
rect 674373 606459 674439 606462
rect 675477 606459 675543 606462
rect 673085 604618 673151 604621
rect 675477 604618 675543 604621
rect 673085 604616 675543 604618
rect 673085 604560 673090 604616
rect 673146 604560 675482 604616
rect 675538 604560 675543 604616
rect 673085 604558 675543 604560
rect 673085 604555 673151 604558
rect 675477 604555 675543 604558
rect 672441 604346 672507 604349
rect 675477 604346 675543 604349
rect 672441 604344 675543 604346
rect 672441 604288 672446 604344
rect 672502 604288 675482 604344
rect 675538 604288 675543 604344
rect 672441 604286 675543 604288
rect 672441 604283 672507 604286
rect 675477 604283 675543 604286
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 673545 603530 673611 603533
rect 675477 603530 675543 603533
rect 673545 603528 675543 603530
rect 673545 603472 673550 603528
rect 673606 603472 675482 603528
rect 675538 603472 675543 603528
rect 673545 603470 675543 603472
rect 673545 603467 673611 603470
rect 675477 603467 675543 603470
rect 674833 603258 674899 603261
rect 669270 603256 674899 603258
rect 669270 603200 674838 603256
rect 674894 603200 674899 603256
rect 669270 603198 674899 603200
rect 666461 603122 666527 603125
rect 669270 603122 669330 603198
rect 674833 603195 674899 603198
rect 666461 603120 669330 603122
rect 666461 603064 666466 603120
rect 666522 603064 669330 603120
rect 666461 603062 669330 603064
rect 666461 603059 666527 603062
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675477 602986 675543 602989
rect 674484 602984 675543 602986
rect 674484 602928 675482 602984
rect 675538 602928 675543 602984
rect 674484 602926 675543 602928
rect 674484 602924 674490 602926
rect 675477 602923 675543 602926
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 668393 601762 668459 601765
rect 675017 601762 675083 601765
rect 668393 601760 675083 601762
rect 668393 601704 668398 601760
rect 668454 601704 675022 601760
rect 675078 601704 675083 601760
rect 668393 601702 675083 601704
rect 668393 601699 668459 601702
rect 675017 601699 675083 601702
rect 48957 601354 49023 601357
rect 41492 601352 49023 601354
rect 41492 601296 48962 601352
rect 49018 601296 49023 601352
rect 41492 601294 49023 601296
rect 48957 601291 49023 601294
rect 674833 601082 674899 601085
rect 675477 601082 675543 601085
rect 674833 601080 675543 601082
rect 674833 601024 674838 601080
rect 674894 601024 675482 601080
rect 675538 601024 675543 601080
rect 674833 601022 675543 601024
rect 674833 601019 674899 601022
rect 675477 601019 675543 601022
rect 54477 600946 54543 600949
rect 41492 600944 54543 600946
rect 41492 600888 54482 600944
rect 54538 600888 54543 600944
rect 41492 600886 54543 600888
rect 54477 600883 54543 600886
rect 44725 600538 44791 600541
rect 41492 600536 44791 600538
rect 41492 600480 44730 600536
rect 44786 600480 44791 600536
rect 41492 600478 44791 600480
rect 44725 600475 44791 600478
rect 675017 600538 675083 600541
rect 675477 600538 675543 600541
rect 675017 600536 675543 600538
rect 675017 600480 675022 600536
rect 675078 600480 675482 600536
rect 675538 600480 675543 600536
rect 675017 600478 675543 600480
rect 675017 600475 675083 600478
rect 675477 600475 675543 600478
rect 44909 600130 44975 600133
rect 41492 600128 44975 600130
rect 41492 600072 44914 600128
rect 44970 600072 44975 600128
rect 41492 600070 44975 600072
rect 44909 600067 44975 600070
rect 44449 599722 44515 599725
rect 675017 599722 675083 599725
rect 41492 599720 44515 599722
rect 41492 599664 44454 599720
rect 44510 599664 44515 599720
rect 41492 599662 44515 599664
rect 44449 599659 44515 599662
rect 663750 599720 675083 599722
rect 663750 599664 675022 599720
rect 675078 599664 675083 599720
rect 663750 599662 675083 599664
rect 660297 599586 660363 599589
rect 663750 599586 663810 599662
rect 675017 599659 675083 599662
rect 660297 599584 663810 599586
rect 660297 599528 660302 599584
rect 660358 599528 663810 599584
rect 660297 599526 663810 599528
rect 660297 599523 660363 599526
rect 44725 599314 44791 599317
rect 41492 599312 44791 599314
rect 41492 599256 44730 599312
rect 44786 599256 44791 599312
rect 41492 599254 44791 599256
rect 44725 599251 44791 599254
rect 674005 599178 674071 599181
rect 675477 599178 675543 599181
rect 674005 599176 675543 599178
rect 674005 599120 674010 599176
rect 674066 599120 675482 599176
rect 675538 599120 675543 599176
rect 674005 599118 675543 599120
rect 674005 599115 674071 599118
rect 675477 599115 675543 599118
rect 45093 598906 45159 598909
rect 41492 598904 45159 598906
rect 41492 598848 45098 598904
rect 45154 598848 45159 598904
rect 41492 598846 45159 598848
rect 45093 598843 45159 598846
rect 670325 598906 670391 598909
rect 674833 598906 674899 598909
rect 670325 598904 674899 598906
rect 670325 598848 670330 598904
rect 670386 598848 674838 598904
rect 674894 598848 674899 598904
rect 670325 598846 674899 598848
rect 670325 598843 670391 598846
rect 674833 598843 674899 598846
rect 45093 598498 45159 598501
rect 41492 598496 45159 598498
rect 41492 598440 45098 598496
rect 45154 598440 45159 598496
rect 41492 598438 45159 598440
rect 45093 598435 45159 598438
rect 673821 598498 673887 598501
rect 675477 598498 675543 598501
rect 673821 598496 675543 598498
rect 673821 598440 673826 598496
rect 673882 598440 675482 598496
rect 675538 598440 675543 598496
rect 673821 598438 675543 598440
rect 673821 598435 673887 598438
rect 675477 598435 675543 598438
rect 45369 598090 45435 598093
rect 41492 598088 45435 598090
rect 41492 598032 45374 598088
rect 45430 598032 45435 598088
rect 41492 598030 45435 598032
rect 45369 598027 45435 598030
rect 674833 598090 674899 598093
rect 675477 598090 675543 598093
rect 674833 598088 675543 598090
rect 674833 598032 674838 598088
rect 674894 598032 675482 598088
rect 675538 598032 675543 598088
rect 674833 598030 675543 598032
rect 674833 598027 674899 598030
rect 675477 598027 675543 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41492 597622 42994 597682
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 42934 597005 42994 597622
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 41045 596866 41111 596869
rect 675017 596866 675083 596869
rect 675477 596866 675543 596869
rect 41045 596864 41124 596866
rect 41045 596808 41050 596864
rect 41106 596808 41124 596864
rect 41045 596806 41124 596808
rect 675017 596864 675543 596866
rect 675017 596808 675022 596864
rect 675078 596808 675482 596864
rect 675538 596808 675543 596864
rect 675017 596806 675543 596808
rect 41045 596803 41111 596806
rect 675017 596803 675083 596806
rect 675477 596803 675543 596806
rect 41822 596458 41828 596460
rect 41492 596398 41828 596458
rect 41822 596396 41828 596398
rect 41892 596396 41898 596460
rect 41229 596050 41295 596053
rect 41229 596048 41308 596050
rect 41229 595992 41234 596048
rect 41290 595992 41308 596048
rect 41229 595990 41308 595992
rect 41229 595987 41295 595990
rect 32397 595642 32463 595645
rect 32397 595640 32476 595642
rect 32397 595584 32402 595640
rect 32458 595584 32476 595640
rect 32397 595582 32476 595584
rect 32397 595579 32463 595582
rect 674925 595506 674991 595509
rect 675385 595506 675451 595509
rect 674925 595504 675451 595506
rect 674925 595448 674930 595504
rect 674986 595448 675390 595504
rect 675446 595448 675451 595504
rect 674925 595446 675451 595448
rect 674925 595443 674991 595446
rect 675385 595443 675451 595446
rect 36537 595234 36603 595237
rect 36524 595232 36603 595234
rect 36524 595176 36542 595232
rect 36598 595176 36603 595232
rect 36524 595174 36603 595176
rect 36537 595171 36603 595174
rect 37917 594826 37983 594829
rect 671245 594826 671311 594829
rect 675477 594826 675543 594829
rect 37917 594824 37996 594826
rect 37917 594768 37922 594824
rect 37978 594768 37996 594824
rect 37917 594766 37996 594768
rect 671245 594824 675543 594826
rect 671245 594768 671250 594824
rect 671306 594768 675482 594824
rect 675538 594768 675543 594824
rect 671245 594766 675543 594768
rect 37917 594763 37983 594766
rect 671245 594763 671311 594766
rect 675477 594763 675543 594766
rect 35157 594418 35223 594421
rect 35157 594416 35236 594418
rect 35157 594360 35162 594416
rect 35218 594360 35236 594416
rect 35157 594358 35236 594360
rect 35157 594355 35223 594358
rect 41321 594010 41387 594013
rect 41308 594008 41387 594010
rect 41308 593952 41326 594008
rect 41382 593952 41387 594008
rect 41308 593950 41387 593952
rect 41321 593947 41387 593950
rect 668853 593738 668919 593741
rect 675385 593738 675451 593741
rect 668853 593736 675451 593738
rect 668853 593680 668858 593736
rect 668914 593680 675390 593736
rect 675446 593680 675451 593736
rect 668853 593678 675451 593680
rect 668853 593675 668919 593678
rect 675385 593675 675451 593678
rect 40677 593602 40743 593605
rect 40677 593600 40756 593602
rect 40677 593544 40682 593600
rect 40738 593544 40756 593600
rect 40677 593542 40756 593544
rect 40677 593539 40743 593542
rect 676070 593404 676076 593468
rect 676140 593466 676146 593468
rect 676990 593466 676996 593468
rect 676140 593406 676996 593466
rect 676140 593404 676146 593406
rect 676990 593404 676996 593406
rect 677060 593404 677066 593468
rect 41822 593194 41828 593196
rect 41492 593134 41828 593194
rect 41822 593132 41828 593134
rect 41892 593132 41898 593196
rect 674189 592922 674255 592925
rect 683297 592922 683363 592925
rect 674189 592920 683363 592922
rect 674189 592864 674194 592920
rect 674250 592864 683302 592920
rect 683358 592864 683363 592920
rect 674189 592862 683363 592864
rect 674189 592859 674255 592862
rect 683297 592859 683363 592862
rect 41873 592786 41939 592789
rect 41492 592784 41939 592786
rect 41492 592728 41878 592784
rect 41934 592728 41939 592784
rect 41492 592726 41939 592728
rect 41873 592723 41939 592726
rect 674557 592650 674623 592653
rect 683113 592650 683179 592653
rect 674557 592648 683179 592650
rect 674557 592592 674562 592648
rect 674618 592592 683118 592648
rect 683174 592592 683179 592648
rect 674557 592590 683179 592592
rect 674557 592587 674623 592590
rect 683113 592587 683179 592590
rect 42190 592378 42196 592380
rect 41492 592318 42196 592378
rect 42190 592316 42196 592318
rect 42260 592316 42266 592380
rect 675334 592316 675340 592380
rect 675404 592378 675410 592380
rect 675753 592378 675819 592381
rect 675404 592376 675819 592378
rect 675404 592320 675758 592376
rect 675814 592320 675819 592376
rect 675404 592318 675819 592320
rect 675404 592316 675410 592318
rect 675753 592315 675819 592318
rect 675569 592108 675635 592109
rect 675518 592106 675524 592108
rect 675478 592046 675524 592106
rect 675588 592104 675635 592108
rect 675630 592048 675635 592104
rect 675518 592044 675524 592046
rect 675588 592044 675635 592048
rect 675569 592043 675635 592044
rect 44449 591970 44515 591973
rect 41492 591968 44515 591970
rect 41492 591912 44454 591968
rect 44510 591912 44515 591968
rect 41492 591910 44515 591912
rect 44449 591907 44515 591910
rect 43846 591562 43852 591564
rect 41492 591502 43852 591562
rect 43846 591500 43852 591502
rect 43916 591500 43922 591564
rect 673729 591154 673795 591157
rect 683481 591154 683547 591157
rect 673729 591152 683547 591154
rect 39990 590749 40050 591124
rect 673729 591096 673734 591152
rect 673790 591096 683486 591152
rect 683542 591096 683547 591152
rect 673729 591094 683547 591096
rect 673729 591091 673795 591094
rect 683481 591091 683547 591094
rect 39941 590744 40050 590749
rect 651465 590746 651531 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 651531 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 651470 590744
rect 651526 590688 651531 590744
rect 650164 590686 651531 590688
rect 39941 590683 40007 590686
rect 651465 590683 651531 590686
rect 43437 590338 43503 590341
rect 41492 590336 43503 590338
rect 41492 590280 43442 590336
rect 43498 590280 43503 590336
rect 41492 590278 43503 590280
rect 43437 590275 43503 590278
rect 40493 589660 40559 589661
rect 40493 589658 40540 589660
rect 40448 589656 40540 589658
rect 40448 589600 40498 589656
rect 40448 589598 40540 589600
rect 40493 589596 40540 589598
rect 40604 589596 40610 589660
rect 40718 589596 40724 589660
rect 40788 589658 40794 589660
rect 41822 589658 41828 589660
rect 40788 589598 41828 589658
rect 40788 589596 40794 589598
rect 41822 589596 41828 589598
rect 41892 589596 41898 589660
rect 40493 589595 40559 589596
rect 40902 589324 40908 589388
rect 40972 589386 40978 589388
rect 42190 589386 42196 589388
rect 40972 589326 42196 589386
rect 40972 589324 40978 589326
rect 42190 589324 42196 589326
rect 42260 589324 42266 589388
rect 675569 586258 675635 586261
rect 676070 586258 676076 586260
rect 675569 586256 676076 586258
rect 675569 586200 675574 586256
rect 675630 586200 676076 586256
rect 675569 586198 676076 586200
rect 675569 586195 675635 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 41689 586122 41755 586125
rect 42517 586122 42583 586125
rect 41689 586120 42583 586122
rect 41689 586064 41694 586120
rect 41750 586064 42522 586120
rect 42578 586064 42583 586120
rect 41689 586062 42583 586064
rect 41689 586059 41755 586062
rect 42517 586059 42583 586062
rect 41873 585850 41939 585853
rect 42425 585850 42491 585853
rect 41873 585848 42491 585850
rect 41873 585792 41878 585848
rect 41934 585792 42430 585848
rect 42486 585792 42491 585848
rect 41873 585790 42491 585792
rect 41873 585787 41939 585790
rect 42425 585787 42491 585790
rect 41505 585442 41571 585445
rect 42006 585442 42012 585444
rect 41505 585440 42012 585442
rect 41505 585384 41510 585440
rect 41566 585384 42012 585440
rect 41505 585382 42012 585384
rect 41505 585379 41571 585382
rect 42006 585380 42012 585382
rect 42076 585380 42082 585444
rect 37917 585170 37983 585173
rect 41822 585170 41828 585172
rect 37917 585168 41828 585170
rect 37917 585112 37922 585168
rect 37978 585112 41828 585168
rect 37917 585110 41828 585112
rect 37917 585107 37983 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 39941 584898 40007 584901
rect 42149 584898 42215 584901
rect 39941 584896 42215 584898
rect 39941 584840 39946 584896
rect 40002 584840 42154 584896
rect 42210 584840 42215 584896
rect 39941 584838 42215 584840
rect 39941 584835 40007 584838
rect 42149 584835 42215 584838
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40677 584626 40743 584629
rect 41086 584626 41092 584628
rect 40677 584624 41092 584626
rect 40677 584568 40682 584624
rect 40738 584568 41092 584624
rect 40677 584566 41092 584568
rect 40677 584563 40743 584566
rect 41086 584564 41092 584566
rect 41156 584564 41162 584628
rect 652017 582994 652083 582997
rect 676029 582994 676095 582997
rect 652017 582992 676095 582994
rect 652017 582936 652022 582992
rect 652078 582936 676034 582992
rect 676090 582936 676095 582992
rect 652017 582934 676095 582936
rect 652017 582931 652083 582934
rect 676029 582931 676095 582934
rect 47577 582450 47643 582453
rect 42014 582448 47643 582450
rect 42014 582392 47582 582448
rect 47638 582392 47643 582448
rect 42014 582390 47643 582392
rect 42014 581498 42074 582390
rect 47577 582387 47643 582390
rect 42241 581498 42307 581501
rect 42014 581496 42307 581498
rect 42014 581440 42246 581496
rect 42302 581440 42307 581496
rect 42014 581438 42307 581440
rect 42241 581435 42307 581438
rect 44449 581090 44515 581093
rect 42198 581088 44515 581090
rect 42198 581032 44454 581088
rect 44510 581032 44515 581088
rect 42198 581030 44515 581032
rect 42198 580821 42258 581030
rect 44449 581027 44515 581030
rect 661677 581090 661743 581093
rect 661677 581088 676292 581090
rect 661677 581032 661682 581088
rect 661738 581032 676292 581088
rect 661677 581030 676292 581032
rect 661677 581027 661743 581030
rect 42198 580816 42307 580821
rect 42198 580760 42246 580816
rect 42302 580760 42307 580816
rect 42198 580758 42307 580760
rect 42241 580755 42307 580758
rect 42006 580484 42012 580548
rect 42076 580546 42082 580548
rect 42425 580546 42491 580549
rect 676262 580546 676322 580652
rect 42076 580544 42491 580546
rect 42076 580488 42430 580544
rect 42486 580488 42491 580544
rect 42076 580486 42491 580488
rect 42076 580484 42082 580486
rect 42425 580483 42491 580486
rect 669270 580486 676322 580546
rect 41086 580212 41092 580276
rect 41156 580274 41162 580276
rect 41781 580274 41847 580277
rect 41156 580272 41847 580274
rect 41156 580216 41786 580272
rect 41842 580216 41847 580272
rect 41156 580214 41847 580216
rect 41156 580212 41162 580214
rect 41781 580211 41847 580214
rect 664437 579730 664503 579733
rect 669270 579730 669330 580486
rect 676029 580274 676095 580277
rect 676029 580272 676292 580274
rect 676029 580216 676034 580272
rect 676090 580216 676292 580272
rect 676029 580214 676292 580216
rect 676029 580211 676095 580214
rect 671429 579866 671495 579869
rect 671429 579864 676292 579866
rect 671429 579808 671434 579864
rect 671490 579808 676292 579864
rect 671429 579806 676292 579808
rect 671429 579803 671495 579806
rect 664437 579728 669330 579730
rect 664437 579672 664442 579728
rect 664498 579672 669330 579728
rect 664437 579670 669330 579672
rect 664437 579667 664503 579670
rect 671521 579458 671587 579461
rect 671521 579456 676292 579458
rect 671521 579400 671526 579456
rect 671582 579400 676292 579456
rect 671521 579398 676292 579400
rect 671521 579395 671587 579398
rect 670785 579050 670851 579053
rect 670785 579048 676292 579050
rect 670785 578992 670790 579048
rect 670846 578992 676292 579048
rect 670785 578990 676292 578992
rect 670785 578987 670851 578990
rect 670785 578642 670851 578645
rect 670785 578640 676292 578642
rect 670785 578584 670790 578640
rect 670846 578584 676292 578640
rect 670785 578582 676292 578584
rect 670785 578579 670851 578582
rect 40718 578172 40724 578236
rect 40788 578234 40794 578236
rect 41781 578234 41847 578237
rect 40788 578232 41847 578234
rect 40788 578176 41786 578232
rect 41842 578176 41847 578232
rect 40788 578174 41847 578176
rect 40788 578172 40794 578174
rect 41781 578171 41847 578174
rect 671705 578234 671771 578237
rect 671705 578232 676292 578234
rect 671705 578176 671710 578232
rect 671766 578176 676292 578232
rect 671705 578174 676292 578176
rect 671705 578171 671771 578174
rect 671061 577826 671127 577829
rect 671061 577824 676292 577826
rect 671061 577768 671066 577824
rect 671122 577768 676292 577824
rect 671061 577766 676292 577768
rect 671061 577763 671127 577766
rect 40902 577492 40908 577556
rect 40972 577554 40978 577556
rect 41781 577554 41847 577557
rect 40972 577552 41847 577554
rect 40972 577496 41786 577552
rect 41842 577496 41847 577552
rect 40972 577494 41847 577496
rect 40972 577492 40978 577494
rect 41781 577491 41847 577494
rect 42425 577420 42491 577421
rect 42374 577418 42380 577420
rect 42334 577358 42380 577418
rect 42444 577416 42491 577420
rect 651465 577418 651531 577421
rect 42486 577360 42491 577416
rect 42374 577356 42380 577358
rect 42444 577356 42491 577360
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 42425 577355 42491 577356
rect 651465 577355 651531 577358
rect 672809 577418 672875 577421
rect 672809 577416 676292 577418
rect 672809 577360 672814 577416
rect 672870 577360 676292 577416
rect 672809 577358 676292 577360
rect 672809 577355 672875 577358
rect 672809 577010 672875 577013
rect 672809 577008 676292 577010
rect 672809 576952 672814 577008
rect 672870 576952 676292 577008
rect 672809 576950 676292 576952
rect 672809 576947 672875 576950
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 42241 576874 42307 576877
rect 40604 576872 42307 576874
rect 40604 576816 42246 576872
rect 42302 576816 42307 576872
rect 40604 576814 42307 576816
rect 40604 576812 40610 576814
rect 42241 576811 42307 576814
rect 675753 576602 675819 576605
rect 675753 576600 676292 576602
rect 675753 576544 675758 576600
rect 675814 576544 676292 576600
rect 675753 576542 676292 576544
rect 675753 576539 675819 576542
rect 671705 576194 671771 576197
rect 671705 576192 676292 576194
rect 671705 576136 671710 576192
rect 671766 576136 676292 576192
rect 671705 576134 676292 576136
rect 671705 576131 671771 576134
rect 676990 575996 676996 576060
rect 677060 575996 677066 576060
rect 676998 575756 677058 575996
rect 682377 575650 682443 575653
rect 682334 575648 682443 575650
rect 682334 575592 682382 575648
rect 682438 575592 682443 575648
rect 682334 575587 682443 575592
rect 682334 575348 682394 575587
rect 669773 574970 669839 574973
rect 669773 574968 676292 574970
rect 669773 574912 669778 574968
rect 669834 574912 676292 574968
rect 669773 574910 676292 574912
rect 669773 574907 669839 574910
rect 672165 574562 672231 574565
rect 672165 574560 676292 574562
rect 672165 574504 672170 574560
rect 672226 574504 676292 574560
rect 672165 574502 676292 574504
rect 672165 574499 672231 574502
rect 668209 574154 668275 574157
rect 668209 574152 676292 574154
rect 668209 574096 668214 574152
rect 668270 574096 676292 574152
rect 668209 574094 676292 574096
rect 668209 574091 668275 574094
rect 683113 574018 683179 574021
rect 683070 574016 683179 574018
rect 683070 573960 683118 574016
rect 683174 573960 683179 574016
rect 683070 573955 683179 573960
rect 42149 573882 42215 573885
rect 42701 573882 42767 573885
rect 42149 573880 42767 573882
rect 42149 573824 42154 573880
rect 42210 573824 42706 573880
rect 42762 573824 42767 573880
rect 42149 573822 42767 573824
rect 42149 573819 42215 573822
rect 42701 573819 42767 573822
rect 683070 573716 683130 573955
rect 669037 573202 669103 573205
rect 676262 573202 676322 573308
rect 683297 573202 683363 573205
rect 669037 573200 676322 573202
rect 669037 573144 669042 573200
rect 669098 573144 676322 573200
rect 669037 573142 676322 573144
rect 683254 573200 683363 573202
rect 683254 573144 683302 573200
rect 683358 573144 683363 573200
rect 669037 573139 669103 573142
rect 683254 573139 683363 573144
rect 683254 572900 683314 573139
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 42057 572658 42123 572661
rect 42374 572658 42380 572660
rect 42057 572656 42380 572658
rect 42057 572600 42062 572656
rect 42118 572600 42380 572656
rect 42057 572598 42380 572600
rect 42057 572595 42123 572598
rect 42374 572596 42380 572598
rect 42444 572596 42450 572660
rect 676814 572492 676874 572732
rect 683481 572386 683547 572389
rect 683438 572384 683547 572386
rect 683438 572328 683486 572384
rect 683542 572328 683547 572384
rect 683438 572323 683547 572328
rect 41822 572188 41828 572252
rect 41892 572250 41898 572252
rect 42241 572250 42307 572253
rect 41892 572248 42307 572250
rect 41892 572192 42246 572248
rect 42302 572192 42307 572248
rect 41892 572190 42307 572192
rect 41892 572188 41898 572190
rect 42241 572187 42307 572190
rect 683438 572084 683498 572323
rect 41454 571916 41460 571980
rect 41524 571978 41530 571980
rect 42609 571978 42675 571981
rect 41524 571976 42675 571978
rect 41524 571920 42614 571976
rect 42670 571920 42675 571976
rect 41524 571918 42675 571920
rect 41524 571916 41530 571918
rect 42609 571915 42675 571918
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 669957 571570 670023 571573
rect 676262 571570 676322 571676
rect 669957 571568 676322 571570
rect 669957 571512 669962 571568
rect 670018 571512 676322 571568
rect 669957 571510 676322 571512
rect 669957 571507 670023 571510
rect 671470 571100 671476 571164
rect 671540 571162 671546 571164
rect 676262 571162 676322 571268
rect 671540 571102 676322 571162
rect 671540 571100 671546 571102
rect 41638 570964 41644 571028
rect 41708 571026 41714 571028
rect 42057 571026 42123 571029
rect 41708 571024 42123 571026
rect 41708 570968 42062 571024
rect 42118 570968 42123 571024
rect 41708 570966 42123 570968
rect 41708 570964 41714 570966
rect 42057 570963 42123 570966
rect 676262 570754 676322 570860
rect 683113 570754 683179 570757
rect 674790 570694 676322 570754
rect 683070 570752 683179 570754
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 669405 570346 669471 570349
rect 674790 570346 674850 570694
rect 669405 570344 674850 570346
rect 669405 570288 669410 570344
rect 669466 570288 674850 570344
rect 669405 570286 674850 570288
rect 683070 570691 683179 570696
rect 669405 570283 669471 570286
rect 683070 570044 683130 570691
rect 670785 569530 670851 569533
rect 676262 569530 676322 569636
rect 670785 569528 676322 569530
rect 670785 569472 670790 569528
rect 670846 569472 676322 569528
rect 670785 569470 676322 569472
rect 670785 569467 670851 569470
rect 42333 569258 42399 569261
rect 62113 569258 62179 569261
rect 42333 569256 62179 569258
rect 42333 569200 42338 569256
rect 42394 569200 62118 569256
rect 62174 569200 62179 569256
rect 42333 569198 62179 569200
rect 42333 569195 42399 569198
rect 62113 569195 62179 569198
rect 668209 564498 668275 564501
rect 675201 564498 675267 564501
rect 668209 564496 675267 564498
rect 668209 564440 668214 564496
rect 668270 564440 675206 564496
rect 675262 564440 675267 564496
rect 668209 564438 675267 564440
rect 668209 564435 668275 564438
rect 675201 564435 675267 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675385 563140 675451 563141
rect 675334 563138 675340 563140
rect 675294 563078 675340 563138
rect 675404 563136 675451 563140
rect 675446 563080 675451 563136
rect 675334 563076 675340 563078
rect 675404 563076 675451 563080
rect 675385 563075 675451 563076
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 672901 559466 672967 559469
rect 675293 559466 675359 559469
rect 672901 559464 675359 559466
rect 672901 559408 672906 559464
rect 672962 559408 675298 559464
rect 675354 559408 675359 559464
rect 672901 559406 675359 559408
rect 672901 559403 672967 559406
rect 675293 559403 675359 559406
rect 669037 559058 669103 559061
rect 675293 559058 675359 559061
rect 669037 559056 675359 559058
rect 669037 559000 669042 559056
rect 669098 559000 675298 559056
rect 675354 559000 675359 559056
rect 669037 558998 675359 559000
rect 669037 558995 669103 558998
rect 675293 558995 675359 558998
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 42057 558514 42123 558517
rect 41492 558512 42123 558514
rect 41492 558456 42062 558512
rect 42118 558456 42123 558512
rect 41492 558454 42123 558456
rect 42057 558451 42123 558454
rect 674649 558378 674715 558381
rect 675385 558378 675451 558381
rect 674649 558376 675451 558378
rect 674649 558320 674654 558376
rect 674710 558320 675390 558376
rect 675446 558320 675451 558376
rect 674649 558318 675451 558320
rect 674649 558315 674715 558318
rect 675385 558315 675451 558318
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 48957 557834 49023 557837
rect 41830 557832 49023 557834
rect 41830 557776 48962 557832
rect 49018 557776 49023 557832
rect 41830 557774 49023 557776
rect 41830 557698 41890 557774
rect 48957 557771 49023 557774
rect 41492 557638 41890 557698
rect 42057 557562 42123 557565
rect 51717 557562 51783 557565
rect 42057 557560 51783 557562
rect 42057 557504 42062 557560
rect 42118 557504 51722 557560
rect 51778 557504 51783 557560
rect 42057 557502 51783 557504
rect 42057 557499 42123 557502
rect 51717 557499 51783 557502
rect 675293 557562 675359 557565
rect 676806 557562 676812 557564
rect 675293 557560 676812 557562
rect 675293 557504 675298 557560
rect 675354 557504 676812 557560
rect 675293 557502 676812 557504
rect 675293 557499 675359 557502
rect 676806 557500 676812 557502
rect 676876 557500 676882 557564
rect 44909 557290 44975 557293
rect 41492 557288 44975 557290
rect 41492 557232 44914 557288
rect 44970 557232 44975 557288
rect 41492 557230 44975 557232
rect 44909 557227 44975 557230
rect 45553 556882 45619 556885
rect 41492 556880 45619 556882
rect 41492 556824 45558 556880
rect 45614 556824 45619 556880
rect 41492 556822 45619 556824
rect 45553 556819 45619 556822
rect 44725 556474 44791 556477
rect 41492 556472 44791 556474
rect 41492 556416 44730 556472
rect 44786 556416 44791 556472
rect 41492 556414 44791 556416
rect 44725 556411 44791 556414
rect 669773 556202 669839 556205
rect 674833 556202 674899 556205
rect 669773 556200 674899 556202
rect 669773 556144 669778 556200
rect 669834 556144 674838 556200
rect 674894 556144 674899 556200
rect 669773 556142 674899 556144
rect 669773 556139 669839 556142
rect 674833 556139 674899 556142
rect 44633 556066 44699 556069
rect 41492 556064 44699 556066
rect 41492 556008 44638 556064
rect 44694 556008 44699 556064
rect 41492 556006 44699 556008
rect 44633 556003 44699 556006
rect 45093 555658 45159 555661
rect 41492 555656 45159 555658
rect 41492 555600 45098 555656
rect 45154 555600 45159 555656
rect 41492 555598 45159 555600
rect 45093 555595 45159 555598
rect 44817 555250 44883 555253
rect 41492 555248 44883 555250
rect 41492 555192 44822 555248
rect 44878 555192 44883 555248
rect 41492 555190 44883 555192
rect 44817 555187 44883 555190
rect 671705 555250 671771 555253
rect 675385 555250 675451 555253
rect 671705 555248 675451 555250
rect 671705 555192 671710 555248
rect 671766 555192 675390 555248
rect 675446 555192 675451 555248
rect 671705 555190 675451 555192
rect 671705 555187 671771 555190
rect 675385 555187 675451 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 674833 554842 674899 554845
rect 675293 554842 675359 554845
rect 674833 554840 675359 554842
rect 674833 554784 674838 554840
rect 674894 554784 675298 554840
rect 675354 554784 675359 554840
rect 674833 554782 675359 554784
rect 674833 554779 674899 554782
rect 675293 554779 675359 554782
rect 44357 554434 44423 554437
rect 41492 554432 44423 554434
rect 41492 554376 44362 554432
rect 44418 554376 44423 554432
rect 41492 554374 44423 554376
rect 44357 554371 44423 554374
rect 35617 554026 35683 554029
rect 35604 554024 35683 554026
rect 35604 553968 35622 554024
rect 35678 553968 35683 554024
rect 35604 553966 35683 553968
rect 35617 553963 35683 553966
rect 658917 554026 658983 554029
rect 675293 554026 675359 554029
rect 658917 554024 675359 554026
rect 658917 553968 658922 554024
rect 658978 553968 675298 554024
rect 675354 553968 675359 554024
rect 658917 553966 675359 553968
rect 658917 553963 658983 553966
rect 675293 553963 675359 553966
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 669589 553482 669655 553485
rect 675385 553482 675451 553485
rect 669589 553480 675451 553482
rect 669589 553424 669594 553480
rect 669650 553424 675390 553480
rect 675446 553424 675451 553480
rect 669589 553422 675451 553424
rect 669589 553419 669655 553422
rect 675385 553419 675451 553422
rect 40953 553410 41019 553413
rect 40910 553408 41019 553410
rect 40910 553352 40958 553408
rect 41014 553352 41019 553408
rect 40910 553347 41019 553352
rect 40910 553180 40970 553347
rect 41689 553074 41755 553077
rect 42006 553074 42012 553076
rect 41689 553072 42012 553074
rect 41689 553016 41694 553072
rect 41750 553016 42012 553072
rect 41689 553014 42012 553016
rect 41689 553011 41755 553014
rect 42006 553012 42012 553014
rect 42076 553012 42082 553076
rect 41137 552802 41203 552805
rect 41124 552800 41203 552802
rect 41124 552744 41142 552800
rect 41198 552744 41203 552800
rect 41124 552742 41203 552744
rect 41137 552739 41203 552742
rect 41321 552394 41387 552397
rect 41308 552392 41387 552394
rect 41308 552336 41326 552392
rect 41382 552336 41387 552392
rect 41308 552334 41387 552336
rect 41321 552331 41387 552334
rect 41781 552122 41847 552125
rect 42977 552122 43043 552125
rect 41781 552120 43043 552122
rect 41781 552064 41786 552120
rect 41842 552064 42982 552120
rect 43038 552064 43043 552120
rect 41781 552062 43043 552064
rect 41781 552059 41847 552062
rect 42977 552059 43043 552062
rect 674189 552122 674255 552125
rect 675385 552122 675451 552125
rect 674189 552120 675451 552122
rect 674189 552064 674194 552120
rect 674250 552064 675390 552120
rect 675446 552064 675451 552120
rect 674189 552062 675451 552064
rect 674189 552059 674255 552062
rect 675385 552059 675451 552062
rect 33777 551986 33843 551989
rect 33764 551984 33843 551986
rect 33764 551928 33782 551984
rect 33838 551928 33843 551984
rect 33764 551926 33843 551928
rect 33777 551923 33843 551926
rect 41689 551850 41755 551853
rect 42190 551850 42196 551852
rect 41689 551848 42196 551850
rect 41689 551792 41694 551848
rect 41750 551792 42196 551848
rect 41689 551790 42196 551792
rect 41689 551787 41755 551790
rect 42190 551788 42196 551790
rect 42260 551788 42266 551852
rect 45001 551578 45067 551581
rect 41492 551576 45067 551578
rect 41492 551520 45006 551576
rect 45062 551520 45067 551576
rect 41492 551518 45067 551520
rect 45001 551515 45067 551518
rect 41321 551170 41387 551173
rect 41308 551168 41387 551170
rect 41308 551112 41326 551168
rect 41382 551112 41387 551168
rect 41308 551110 41387 551112
rect 41321 551107 41387 551110
rect 45369 550898 45435 550901
rect 651465 550898 651531 550901
rect 41830 550896 45435 550898
rect 41830 550840 45374 550896
rect 45430 550840 45435 550896
rect 41830 550838 45435 550840
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 41830 550796 41890 550838
rect 45369 550835 45435 550838
rect 651465 550835 651531 550838
rect 41462 550736 41890 550796
rect 675753 550762 675819 550765
rect 677174 550762 677180 550764
rect 675753 550760 677180 550762
rect 41462 550732 41522 550736
rect 675753 550704 675758 550760
rect 675814 550704 677180 550760
rect 675753 550702 677180 550704
rect 675753 550699 675819 550702
rect 677174 550700 677180 550702
rect 677244 550700 677250 550764
rect 41781 550626 41847 550629
rect 42793 550626 42859 550629
rect 41781 550624 42859 550626
rect 41781 550568 41786 550624
rect 41842 550568 42798 550624
rect 42854 550568 42859 550624
rect 41781 550566 42859 550568
rect 41781 550563 41847 550566
rect 42793 550563 42859 550566
rect 41492 550294 41936 550354
rect 41876 550218 41936 550294
rect 42057 550218 42123 550221
rect 41876 550216 42123 550218
rect 41876 550160 42062 550216
rect 42118 550160 42123 550216
rect 41876 550158 42123 550160
rect 42057 550155 42123 550158
rect 41781 549946 41847 549949
rect 41492 549944 41847 549946
rect 41492 549888 41786 549944
rect 41842 549888 41847 549944
rect 41492 549886 41847 549888
rect 41781 549883 41847 549886
rect 675109 549674 675175 549677
rect 675477 549674 675543 549677
rect 675109 549672 675543 549674
rect 675109 549616 675114 549672
rect 675170 549616 675482 549672
rect 675538 549616 675543 549672
rect 675109 549614 675543 549616
rect 675109 549611 675175 549614
rect 675477 549611 675543 549614
rect 43161 549538 43227 549541
rect 41492 549536 43227 549538
rect 41492 549480 43166 549536
rect 43222 549480 43227 549536
rect 41492 549478 43227 549480
rect 43161 549475 43227 549478
rect 44173 549130 44239 549133
rect 41492 549128 44239 549130
rect 41492 549072 44178 549128
rect 44234 549072 44239 549128
rect 41492 549070 44239 549072
rect 44173 549067 44239 549070
rect 45185 548722 45251 548725
rect 41492 548720 45251 548722
rect 41492 548664 45190 548720
rect 45246 548664 45251 548720
rect 41492 548662 45251 548664
rect 45185 548659 45251 548662
rect 672809 548450 672875 548453
rect 675477 548450 675543 548453
rect 672809 548448 675543 548450
rect 672809 548392 672814 548448
rect 672870 548392 675482 548448
rect 675538 548392 675543 548448
rect 672809 548390 675543 548392
rect 672809 548387 672875 548390
rect 675477 548387 675543 548390
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 28766 547498 28826 547890
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 674833 547634 674899 547637
rect 675845 547634 675911 547637
rect 674833 547632 675911 547634
rect 674833 547576 674838 547632
rect 674894 547576 675850 547632
rect 675906 547576 675911 547632
rect 674833 547574 675911 547576
rect 674833 547571 674899 547574
rect 675845 547571 675911 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 43805 547090 43871 547093
rect 41492 547088 43871 547090
rect 41492 547032 43810 547088
rect 43866 547032 43871 547088
rect 41492 547030 43871 547032
rect 43805 547027 43871 547030
rect 674373 547090 674439 547093
rect 683205 547090 683271 547093
rect 674373 547088 683271 547090
rect 674373 547032 674378 547088
rect 674434 547032 683210 547088
rect 683266 547032 683271 547088
rect 674373 547030 683271 547032
rect 674373 547027 674439 547030
rect 683205 547027 683271 547030
rect 675293 546546 675359 546549
rect 675518 546546 675524 546548
rect 675293 546544 675524 546546
rect 675293 546488 675298 546544
rect 675354 546488 675524 546544
rect 675293 546486 675524 546488
rect 675293 546483 675359 546486
rect 675518 546484 675524 546486
rect 675588 546484 675594 546548
rect 676070 546484 676076 546548
rect 676140 546546 676146 546548
rect 679617 546546 679683 546549
rect 676140 546544 679683 546546
rect 676140 546488 679622 546544
rect 679678 546488 679683 546544
rect 676140 546486 679683 546488
rect 676140 546484 676146 546486
rect 679617 546483 679683 546486
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 672625 546274 672691 546277
rect 676397 546274 676463 546277
rect 672625 546272 676463 546274
rect 672625 546216 672630 546272
rect 672686 546216 676402 546272
rect 676458 546216 676463 546272
rect 672625 546214 676463 546216
rect 672625 546211 672691 546214
rect 676397 546211 676463 546214
rect 674833 546002 674899 546005
rect 675334 546002 675340 546004
rect 674833 546000 675340 546002
rect 674833 545944 674838 546000
rect 674894 545944 675340 546000
rect 674833 545942 675340 545944
rect 674833 545939 674899 545942
rect 675334 545940 675340 545942
rect 675404 545940 675410 546004
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40534 545668 40540 545732
rect 40604 545730 40610 545732
rect 42057 545730 42123 545733
rect 40604 545728 42123 545730
rect 40604 545672 42062 545728
rect 42118 545672 42123 545728
rect 40604 545670 42123 545672
rect 40604 545668 40610 545670
rect 42057 545667 42123 545670
rect 674005 545730 674071 545733
rect 683389 545730 683455 545733
rect 674005 545728 683455 545730
rect 674005 545672 674010 545728
rect 674066 545672 683394 545728
rect 683450 545672 683455 545728
rect 674005 545670 683455 545672
rect 674005 545667 674071 545670
rect 683389 545667 683455 545670
rect 40718 545396 40724 545460
rect 40788 545458 40794 545460
rect 41505 545458 41571 545461
rect 40788 545456 41571 545458
rect 40788 545400 41510 545456
rect 41566 545400 41571 545456
rect 40788 545398 41571 545400
rect 40788 545396 40794 545398
rect 41505 545395 41571 545398
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 670141 537842 670207 537845
rect 676029 537842 676095 537845
rect 670141 537840 676095 537842
rect 670141 537784 670146 537840
rect 670202 537784 676034 537840
rect 676090 537784 676095 537840
rect 670141 537782 676095 537784
rect 670141 537779 670207 537782
rect 676029 537779 676095 537782
rect 42517 537570 42583 537573
rect 44173 537570 44239 537573
rect 651465 537570 651531 537573
rect 42517 537568 44239 537570
rect 42517 537512 42522 537568
rect 42578 537512 44178 537568
rect 44234 537512 44239 537568
rect 42517 537510 44239 537512
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 42517 537507 42583 537510
rect 44173 537507 44239 537510
rect 651465 537507 651531 537510
rect 40534 536964 40540 537028
rect 40604 537026 40610 537028
rect 41781 537026 41847 537029
rect 40604 537024 41847 537026
rect 40604 536968 41786 537024
rect 41842 536968 41847 537024
rect 40604 536966 41847 536968
rect 40604 536964 40610 536966
rect 41781 536963 41847 536966
rect 42149 537026 42215 537029
rect 45185 537026 45251 537029
rect 42149 537024 45251 537026
rect 42149 536968 42154 537024
rect 42210 536968 45190 537024
rect 45246 536968 45251 537024
rect 42149 536966 45251 536968
rect 42149 536963 42215 536966
rect 45185 536963 45251 536966
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 668577 535875 668643 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 674005 535394 674071 535397
rect 674005 535392 676322 535394
rect 674005 535336 674010 535392
rect 674066 535336 676322 535392
rect 674005 535334 676322 535336
rect 674005 535331 674071 535334
rect 676262 535296 676322 535334
rect 40718 535196 40724 535260
rect 40788 535258 40794 535260
rect 41781 535258 41847 535261
rect 40788 535256 41847 535258
rect 40788 535200 41786 535256
rect 41842 535200 41847 535256
rect 40788 535198 41847 535200
rect 40788 535196 40794 535198
rect 41781 535195 41847 535198
rect 670969 535122 671035 535125
rect 674465 535122 674531 535125
rect 670969 535120 674531 535122
rect 670969 535064 670974 535120
rect 671030 535064 674470 535120
rect 674526 535064 674531 535120
rect 670969 535062 674531 535064
rect 670969 535059 671035 535062
rect 674465 535059 674531 535062
rect 671429 534714 671495 534717
rect 676262 534714 676322 534888
rect 671429 534712 676322 534714
rect 671429 534656 671434 534712
rect 671490 534656 676322 534712
rect 671429 534654 676322 534656
rect 671429 534651 671495 534654
rect 671521 534442 671587 534445
rect 676262 534442 676322 534480
rect 671521 534440 676322 534442
rect 671521 534384 671526 534440
rect 671582 534384 676322 534440
rect 671521 534382 676322 534384
rect 671521 534379 671587 534382
rect 667197 534170 667263 534173
rect 674005 534170 674071 534173
rect 667197 534168 674071 534170
rect 667197 534112 667202 534168
rect 667258 534112 674010 534168
rect 674066 534112 674071 534168
rect 667197 534110 674071 534112
rect 667197 534107 667263 534110
rect 674005 534107 674071 534110
rect 674465 534170 674531 534173
rect 674465 534168 676322 534170
rect 674465 534112 674470 534168
rect 674526 534112 676322 534168
rect 674465 534110 676322 534112
rect 674465 534107 674531 534110
rect 676262 534072 676322 534110
rect 42149 533898 42215 533901
rect 42977 533898 43043 533901
rect 42149 533896 43043 533898
rect 42149 533840 42154 533896
rect 42210 533840 42982 533896
rect 43038 533840 43043 533896
rect 42149 533838 43043 533840
rect 42149 533835 42215 533838
rect 42977 533835 43043 533838
rect 672625 533898 672691 533901
rect 672625 533896 676322 533898
rect 672625 533840 672630 533896
rect 672686 533840 676322 533896
rect 672625 533838 676322 533840
rect 672625 533835 672691 533838
rect 676262 533664 676322 533838
rect 671061 533490 671127 533493
rect 671061 533488 676322 533490
rect 671061 533432 671066 533488
rect 671122 533432 676322 533488
rect 671061 533430 676322 533432
rect 671061 533427 671127 533430
rect 676262 533256 676322 533430
rect 42241 533218 42307 533221
rect 43161 533218 43227 533221
rect 42241 533216 43227 533218
rect 42241 533160 42246 533216
rect 42302 533160 43166 533216
rect 43222 533160 43227 533216
rect 42241 533158 43227 533160
rect 42241 533155 42307 533158
rect 43161 533155 43227 533158
rect 671061 532946 671127 532949
rect 671061 532944 676322 532946
rect 671061 532888 671066 532944
rect 671122 532888 676322 532944
rect 671061 532886 676322 532888
rect 671061 532883 671127 532886
rect 676262 532848 676322 532886
rect 42517 532810 42583 532813
rect 45369 532810 45435 532813
rect 42517 532808 45435 532810
rect 42517 532752 42522 532808
rect 42578 532752 45374 532808
rect 45430 532752 45435 532808
rect 42517 532750 45435 532752
rect 42517 532747 42583 532750
rect 45369 532747 45435 532750
rect 62113 532810 62179 532813
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 62113 532747 62179 532750
rect 672257 532674 672323 532677
rect 672257 532672 676322 532674
rect 672257 532616 672262 532672
rect 672318 532616 676322 532672
rect 672257 532614 676322 532616
rect 672257 532611 672323 532614
rect 676262 532440 676322 532614
rect 673821 532266 673887 532269
rect 683573 532266 683639 532269
rect 673821 532264 683639 532266
rect 673821 532208 673826 532264
rect 673882 532208 683578 532264
rect 683634 532208 683639 532264
rect 673821 532206 683639 532208
rect 673821 532203 673887 532206
rect 683573 532203 683639 532206
rect 673821 531858 673887 531861
rect 676262 531858 676322 532032
rect 673821 531856 676322 531858
rect 673821 531800 673826 531856
rect 673882 531800 676322 531856
rect 673821 531798 676322 531800
rect 683205 531858 683271 531861
rect 683205 531856 683314 531858
rect 683205 531800 683210 531856
rect 683266 531800 683314 531856
rect 673821 531795 673887 531798
rect 683205 531795 683314 531800
rect 683254 531624 683314 531795
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 679617 531042 679683 531045
rect 679574 531040 679683 531042
rect 679574 530984 679622 531040
rect 679678 530984 679683 531040
rect 679574 530979 679683 530984
rect 679574 530808 679634 530979
rect 41454 530572 41460 530636
rect 41524 530634 41530 530636
rect 42517 530634 42583 530637
rect 41524 530632 42583 530634
rect 41524 530576 42522 530632
rect 42578 530576 42583 530632
rect 41524 530574 42583 530576
rect 41524 530572 41530 530574
rect 42517 530571 42583 530574
rect 673177 530634 673243 530637
rect 673177 530632 676322 530634
rect 673177 530576 673182 530632
rect 673238 530576 676322 530632
rect 673177 530574 676322 530576
rect 673177 530571 673243 530574
rect 676262 530400 676322 530574
rect 42149 530090 42215 530093
rect 42701 530090 42767 530093
rect 42149 530088 42767 530090
rect 42149 530032 42154 530088
rect 42210 530032 42706 530088
rect 42762 530032 42767 530088
rect 42149 530030 42767 530032
rect 42149 530027 42215 530030
rect 42701 530027 42767 530030
rect 666461 529954 666527 529957
rect 676262 529954 676322 529992
rect 666461 529952 676322 529954
rect 666461 529896 666466 529952
rect 666522 529896 676322 529952
rect 666461 529894 676322 529896
rect 666461 529891 666527 529894
rect 42609 529682 42675 529685
rect 45001 529682 45067 529685
rect 42609 529680 45067 529682
rect 42609 529624 42614 529680
rect 42670 529624 45006 529680
rect 45062 529624 45067 529680
rect 42609 529622 45067 529624
rect 42609 529619 42675 529622
rect 45001 529619 45067 529622
rect 670601 529682 670667 529685
rect 675753 529682 675819 529685
rect 670601 529680 675819 529682
rect 670601 529624 670606 529680
rect 670662 529624 675758 529680
rect 675814 529624 675819 529680
rect 670601 529622 675819 529624
rect 670601 529619 670667 529622
rect 675753 529619 675819 529622
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 676262 529410 676322 529584
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 669270 529350 676322 529410
rect 41638 529076 41644 529140
rect 41708 529138 41714 529140
rect 42885 529138 42951 529141
rect 41708 529136 42951 529138
rect 41708 529080 42890 529136
rect 42946 529080 42951 529136
rect 41708 529078 42951 529080
rect 41708 529076 41714 529078
rect 42885 529075 42951 529078
rect 668853 528594 668919 528597
rect 669270 528594 669330 529350
rect 675753 529206 675819 529209
rect 675753 529204 676292 529206
rect 675753 529148 675758 529204
rect 675814 529148 676292 529204
rect 675753 529146 676292 529148
rect 675753 529143 675819 529146
rect 672441 529002 672507 529005
rect 672441 529000 676322 529002
rect 672441 528944 672446 529000
rect 672502 528944 676322 529000
rect 672441 528942 676322 528944
rect 672441 528939 672507 528942
rect 676262 528768 676322 528942
rect 668853 528592 669330 528594
rect 668853 528536 668858 528592
rect 668914 528536 669330 528592
rect 668853 528534 669330 528536
rect 668853 528531 668919 528534
rect 673637 528458 673703 528461
rect 673637 528456 676322 528458
rect 673637 528400 673642 528456
rect 673698 528400 676322 528456
rect 673637 528398 676322 528400
rect 673637 528395 673703 528398
rect 676262 528360 676322 528398
rect 670325 528186 670391 528189
rect 670325 528184 676322 528186
rect 670325 528128 670330 528184
rect 670386 528128 676322 528184
rect 670325 528126 676322 528128
rect 670325 528123 670391 528126
rect 676262 527952 676322 528126
rect 683389 527778 683455 527781
rect 683389 527776 683498 527778
rect 683389 527720 683394 527776
rect 683450 527720 683498 527776
rect 683389 527715 683498 527720
rect 683438 527544 683498 527715
rect 674414 527036 674420 527100
rect 674484 527098 674490 527100
rect 676262 527098 676322 527136
rect 674484 527038 676322 527098
rect 674484 527036 674490 527038
rect 668393 526554 668459 526557
rect 676262 526554 676322 526728
rect 668393 526552 676322 526554
rect 668393 526496 668398 526552
rect 668454 526496 676322 526552
rect 668393 526494 676322 526496
rect 683573 526554 683639 526557
rect 683573 526552 683682 526554
rect 683573 526496 683578 526552
rect 683634 526496 683682 526552
rect 668393 526491 668459 526494
rect 683573 526491 683682 526496
rect 683622 526320 683682 526491
rect 676814 525741 676874 525912
rect 671245 525738 671311 525741
rect 671245 525736 676322 525738
rect 671245 525680 671250 525736
rect 671306 525680 676322 525736
rect 671245 525678 676322 525680
rect 676814 525736 676923 525741
rect 676814 525680 676862 525736
rect 676918 525680 676923 525736
rect 676814 525678 676923 525680
rect 671245 525675 671311 525678
rect 676262 525096 676322 525678
rect 676857 525675 676923 525678
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 674925 503842 674991 503845
rect 675845 503842 675911 503845
rect 674925 503840 675911 503842
rect 674925 503784 674930 503840
rect 674986 503784 675850 503840
rect 675906 503784 675911 503840
rect 674925 503782 675911 503784
rect 674925 503779 674991 503782
rect 675845 503779 675911 503782
rect 676806 503644 676812 503708
rect 676876 503706 676882 503708
rect 683205 503706 683271 503709
rect 676876 503704 683271 503706
rect 676876 503648 683210 503704
rect 683266 503648 683271 503704
rect 676876 503646 683271 503648
rect 676876 503644 676882 503646
rect 683205 503643 683271 503646
rect 675017 503570 675083 503573
rect 676029 503570 676095 503573
rect 675017 503568 676095 503570
rect 675017 503512 675022 503568
rect 675078 503512 676034 503568
rect 676090 503512 676095 503568
rect 675017 503510 676095 503512
rect 675017 503507 675083 503510
rect 676029 503507 676095 503510
rect 675017 503298 675083 503301
rect 676029 503298 676095 503301
rect 675017 503296 676095 503298
rect 675017 503240 675022 503296
rect 675078 503240 676034 503296
rect 676090 503240 676095 503296
rect 675017 503238 676095 503240
rect 675017 503235 675083 503238
rect 676029 503235 676095 503238
rect 669405 500986 669471 500989
rect 674925 500986 674991 500989
rect 669405 500984 674991 500986
rect 669405 500928 669410 500984
rect 669466 500928 674930 500984
rect 674986 500928 674991 500984
rect 669405 500926 674991 500928
rect 669405 500923 669471 500926
rect 674925 500923 674991 500926
rect 652569 497722 652635 497725
rect 650164 497720 652635 497722
rect 650164 497664 652574 497720
rect 652630 497664 652635 497720
rect 650164 497662 652635 497664
rect 652569 497659 652635 497662
rect 666001 494730 666067 494733
rect 683573 494730 683639 494733
rect 666001 494728 683639 494730
rect 666001 494672 666006 494728
rect 666062 494672 683578 494728
rect 683634 494672 683639 494728
rect 666001 494670 683639 494672
rect 666001 494667 666067 494670
rect 683573 494667 683639 494670
rect 664621 494050 664687 494053
rect 676029 494050 676095 494053
rect 664621 494048 676095 494050
rect 664621 493992 664626 494048
rect 664682 493992 676034 494048
rect 676090 493992 676095 494048
rect 664621 493990 676095 493992
rect 664621 493987 664687 493990
rect 676029 493987 676095 493990
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 677317 492420 677383 492421
rect 677317 492416 677364 492420
rect 677428 492418 677434 492420
rect 677317 492360 677322 492416
rect 677317 492356 677364 492360
rect 677428 492358 677474 492418
rect 677428 492356 677434 492358
rect 677317 492355 677383 492356
rect 663750 492086 676292 492146
rect 662045 492010 662111 492013
rect 663750 492010 663810 492086
rect 662045 492008 663810 492010
rect 662045 491952 662050 492008
rect 662106 491952 663810 492008
rect 662045 491950 663810 491952
rect 662045 491947 662111 491950
rect 683389 491738 683455 491741
rect 683389 491736 683468 491738
rect 683389 491680 683394 491736
rect 683450 491680 683468 491736
rect 683389 491678 683468 491680
rect 683389 491675 683455 491678
rect 683573 491330 683639 491333
rect 683573 491328 683652 491330
rect 683573 491272 683578 491328
rect 683634 491272 683652 491328
rect 683573 491270 683652 491272
rect 683573 491267 683639 491270
rect 671521 490922 671587 490925
rect 671521 490920 676292 490922
rect 671521 490864 671526 490920
rect 671582 490864 676292 490920
rect 671521 490862 676292 490864
rect 671521 490859 671587 490862
rect 675886 490452 675892 490516
rect 675956 490514 675962 490516
rect 675956 490454 676292 490514
rect 675956 490452 675962 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 672441 489698 672507 489701
rect 672441 489696 676292 489698
rect 672441 489640 672446 489696
rect 672502 489640 676292 489696
rect 672441 489638 676292 489640
rect 672441 489635 672507 489638
rect 671061 489290 671127 489293
rect 671061 489288 676292 489290
rect 671061 489232 671066 489288
rect 671122 489232 676292 489288
rect 671061 489230 676292 489232
rect 671061 489227 671127 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 673361 488474 673427 488477
rect 673361 488472 676292 488474
rect 673361 488416 673366 488472
rect 673422 488416 676292 488472
rect 673361 488414 676292 488416
rect 673361 488411 673427 488414
rect 672625 488066 672691 488069
rect 672625 488064 676292 488066
rect 672625 488008 672630 488064
rect 672686 488008 676292 488064
rect 672625 488006 676292 488008
rect 672625 488003 672691 488006
rect 680997 487658 681063 487661
rect 680997 487656 681076 487658
rect 680997 487600 681002 487656
rect 681058 487600 681076 487656
rect 680997 487598 681076 487600
rect 680997 487595 681063 487598
rect 677317 487250 677383 487253
rect 677317 487248 677396 487250
rect 677317 487192 677322 487248
rect 677378 487192 677396 487248
rect 677317 487190 677396 487192
rect 677317 487187 677383 487190
rect 679617 486842 679683 486845
rect 679604 486840 679683 486842
rect 679604 486784 679622 486840
rect 679678 486784 679683 486840
rect 679604 486782 679683 486784
rect 679617 486779 679683 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 671705 486026 671771 486029
rect 671705 486024 676292 486026
rect 671705 485968 671710 486024
rect 671766 485968 676292 486024
rect 671705 485966 676292 485968
rect 671705 485963 671771 485966
rect 672901 485618 672967 485621
rect 672901 485616 676292 485618
rect 672901 485560 672906 485616
rect 672962 485560 676292 485616
rect 672901 485558 676292 485560
rect 672901 485555 672967 485558
rect 668209 485210 668275 485213
rect 668209 485208 676292 485210
rect 668209 485152 668214 485208
rect 668270 485152 676292 485208
rect 668209 485150 676292 485152
rect 668209 485147 668275 485150
rect 673085 484802 673151 484805
rect 673085 484800 676292 484802
rect 673085 484744 673090 484800
rect 673146 484744 676292 484800
rect 673085 484742 676292 484744
rect 673085 484739 673151 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 674189 483986 674255 483989
rect 674189 483984 676292 483986
rect 674189 483928 674194 483984
rect 674250 483928 676292 483984
rect 674189 483926 676292 483928
rect 674189 483923 674255 483926
rect 669773 483578 669839 483581
rect 669773 483576 676292 483578
rect 669773 483520 669778 483576
rect 669834 483520 676292 483576
rect 669773 483518 676292 483520
rect 669773 483515 669839 483518
rect 669037 483170 669103 483173
rect 669037 483168 676292 483170
rect 669037 483112 669042 483168
rect 669098 483112 676292 483168
rect 669037 483110 676292 483112
rect 669037 483107 669103 483110
rect 683205 482762 683271 482765
rect 683205 482760 683284 482762
rect 683205 482704 683210 482760
rect 683266 482704 683284 482760
rect 683205 482702 683284 482704
rect 683205 482699 683271 482702
rect 669589 482354 669655 482357
rect 669589 482352 676292 482354
rect 669589 482296 669594 482352
rect 669650 482296 676292 482352
rect 669589 482294 676292 482296
rect 669589 482291 669655 482294
rect 675845 481946 675911 481949
rect 675845 481944 676292 481946
rect 675845 481888 675850 481944
rect 675906 481888 676292 481944
rect 675845 481886 676292 481888
rect 675845 481883 675911 481886
rect 682377 481538 682443 481541
rect 682364 481536 682443 481538
rect 682364 481508 682382 481536
rect 682334 481480 682382 481508
rect 682438 481480 682443 481536
rect 682334 481475 682443 481480
rect 682334 481100 682394 481475
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 673678 475356 673684 475420
rect 673748 475418 673754 475420
rect 674046 475418 674052 475420
rect 673748 475358 674052 475418
rect 673748 475356 673754 475358
rect 674046 475356 674052 475358
rect 674116 475356 674122 475420
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 673678 464748 673684 464812
rect 673748 464810 673754 464812
rect 674741 464810 674807 464813
rect 673748 464808 674807 464810
rect 673748 464752 674746 464808
rect 674802 464752 674807 464808
rect 673748 464750 674807 464752
rect 673748 464748 673754 464750
rect 674741 464747 674807 464750
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 673821 456922 673887 456925
rect 674741 456922 674807 456925
rect 673821 456920 674807 456922
rect 673821 456864 673826 456920
rect 673882 456864 674746 456920
rect 674802 456864 674807 456920
rect 673821 456862 674807 456864
rect 673821 456859 673887 456862
rect 674741 456859 674807 456862
rect 669221 456242 669287 456245
rect 673941 456242 674007 456245
rect 669221 456240 674007 456242
rect 669221 456184 669226 456240
rect 669282 456184 673946 456240
rect 674002 456184 674007 456240
rect 669221 456182 674007 456184
rect 669221 456179 669287 456182
rect 673941 456179 674007 456182
rect 673591 455698 673657 455701
rect 676765 455698 676831 455701
rect 673591 455696 676831 455698
rect 673591 455640 673596 455696
rect 673652 455640 676770 455696
rect 676826 455640 676831 455696
rect 673591 455638 676831 455640
rect 673591 455635 673657 455638
rect 676765 455635 676831 455638
rect 671981 455426 672047 455429
rect 673499 455426 673565 455429
rect 671981 455424 673565 455426
rect 671981 455368 671986 455424
rect 672042 455368 673504 455424
rect 673560 455368 673565 455424
rect 671981 455366 673565 455368
rect 671981 455363 672047 455366
rect 673499 455363 673565 455366
rect 670877 455154 670943 455157
rect 671981 455154 672047 455157
rect 670877 455152 672047 455154
rect 670877 455096 670882 455152
rect 670938 455096 671986 455152
rect 672042 455096 672047 455152
rect 670877 455094 672047 455096
rect 670877 455091 670943 455094
rect 671981 455091 672047 455094
rect 673381 455154 673447 455157
rect 673862 455154 673868 455156
rect 673381 455152 673868 455154
rect 673381 455096 673386 455152
rect 673442 455096 673868 455152
rect 673381 455094 673868 455096
rect 673381 455091 673447 455094
rect 673862 455092 673868 455094
rect 673932 455092 673938 455156
rect 673157 454882 673223 454885
rect 674925 454882 674991 454885
rect 673157 454880 674991 454882
rect 673157 454824 673162 454880
rect 673218 454824 674930 454880
rect 674986 454824 674991 454880
rect 673157 454822 674991 454824
rect 673157 454819 673223 454822
rect 674925 454819 674991 454822
rect 62113 454610 62179 454613
rect 673039 454610 673105 454613
rect 675477 454610 675543 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 673039 454608 675543 454610
rect 673039 454552 673044 454608
rect 673100 454552 675482 454608
rect 675538 454552 675543 454608
rect 673039 454550 675543 454552
rect 62113 454547 62179 454550
rect 673039 454547 673105 454550
rect 675477 454547 675543 454550
rect 672947 454338 673013 454341
rect 675661 454338 675727 454341
rect 672947 454336 675727 454338
rect 672947 454280 672952 454336
rect 673008 454280 675666 454336
rect 675722 454280 675727 454336
rect 672947 454278 675727 454280
rect 672947 454275 673013 454278
rect 675661 454275 675727 454278
rect 672809 454066 672875 454069
rect 676029 454066 676095 454069
rect 672809 454064 676095 454066
rect 672809 454008 672814 454064
rect 672870 454008 676034 454064
rect 676090 454008 676095 454064
rect 672809 454006 676095 454008
rect 672809 454003 672875 454006
rect 676029 454003 676095 454006
rect 672257 453794 672323 453797
rect 675845 453794 675911 453797
rect 672257 453792 675911 453794
rect 672257 453736 672262 453792
rect 672318 453736 675850 453792
rect 675906 453736 675911 453792
rect 672257 453734 675911 453736
rect 672257 453731 672323 453734
rect 675845 453731 675911 453734
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45553 429722 45619 429725
rect 41492 429720 45619 429722
rect 41492 429664 45558 429720
rect 45614 429664 45619 429720
rect 41492 429662 45619 429664
rect 45553 429659 45619 429662
rect 45001 429314 45067 429317
rect 41492 429312 45067 429314
rect 41492 429256 45006 429312
rect 45062 429256 45067 429312
rect 41492 429254 45067 429256
rect 45001 429251 45067 429254
rect 44633 428906 44699 428909
rect 41492 428904 44699 428906
rect 41492 428848 44638 428904
rect 44694 428848 44699 428904
rect 41492 428846 44699 428848
rect 44633 428843 44699 428846
rect 44173 428498 44239 428501
rect 41492 428496 44239 428498
rect 41492 428440 44178 428496
rect 44234 428440 44239 428496
rect 41492 428438 44239 428440
rect 44173 428435 44239 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44817 428090 44883 428093
rect 41492 428088 44883 428090
rect 41492 428032 44822 428088
rect 44878 428032 44883 428088
rect 41492 428030 44883 428032
rect 44817 428027 44883 428030
rect 45185 427682 45251 427685
rect 41492 427680 45251 427682
rect 41492 427624 45190 427680
rect 45246 427624 45251 427680
rect 41492 427622 45251 427624
rect 45185 427619 45251 427622
rect 44357 427274 44423 427277
rect 41492 427272 44423 427274
rect 41492 427216 44362 427272
rect 44418 427216 44423 427272
rect 41492 427214 44423 427216
rect 44357 427211 44423 427214
rect 44449 426866 44515 426869
rect 41492 426864 44515 426866
rect 41492 426808 44454 426864
rect 44510 426808 44515 426864
rect 41492 426806 44515 426808
rect 44449 426803 44515 426806
rect 46933 426458 46999 426461
rect 41492 426456 46999 426458
rect 41492 426400 46938 426456
rect 46994 426400 46999 426456
rect 41492 426398 46999 426400
rect 46933 426395 46999 426398
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 40953 425642 41019 425645
rect 40940 425640 41019 425642
rect 40940 425584 40958 425640
rect 41014 425584 41019 425640
rect 40940 425582 41019 425584
rect 40953 425579 41019 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 36537 424418 36603 424421
rect 36524 424416 36603 424418
rect 36524 424360 36542 424416
rect 36598 424360 36603 424416
rect 36524 424358 36603 424360
rect 36537 424355 36603 424358
rect 41321 424010 41387 424013
rect 41308 424008 41387 424010
rect 41308 423952 41326 424008
rect 41382 423952 41387 424008
rect 41308 423950 41387 423952
rect 41321 423947 41387 423950
rect 47117 423602 47183 423605
rect 41492 423600 47183 423602
rect 41492 423544 47122 423600
rect 47178 423544 47183 423600
rect 41492 423542 47183 423544
rect 47117 423539 47183 423542
rect 43069 423194 43135 423197
rect 41492 423192 43135 423194
rect 41492 423136 43074 423192
rect 43130 423136 43135 423192
rect 41492 423134 43135 423136
rect 43069 423131 43135 423134
rect 41965 422786 42031 422789
rect 41492 422784 42031 422786
rect 41492 422728 41970 422784
rect 42026 422728 42031 422784
rect 41492 422726 42031 422728
rect 41965 422723 42031 422726
rect 45369 422378 45435 422381
rect 41492 422376 45435 422378
rect 41492 422320 45374 422376
rect 45430 422320 45435 422376
rect 41492 422318 45435 422320
rect 45369 422315 45435 422318
rect 41781 421970 41847 421973
rect 41492 421968 41847 421970
rect 41492 421912 41786 421968
rect 41842 421912 41847 421968
rect 41492 421910 41847 421912
rect 41781 421907 41847 421910
rect 44633 421562 44699 421565
rect 41492 421560 44699 421562
rect 41492 421504 44638 421560
rect 44694 421504 44699 421560
rect 41492 421502 44699 421504
rect 44633 421499 44699 421502
rect 43253 421154 43319 421157
rect 41492 421152 43319 421154
rect 41492 421096 43258 421152
rect 43314 421096 43319 421152
rect 41492 421094 43319 421096
rect 43253 421091 43319 421094
rect 44817 420746 44883 420749
rect 41492 420744 44883 420746
rect 41492 420688 44822 420744
rect 44878 420688 44883 420744
rect 41492 420686 44883 420688
rect 44817 420683 44883 420686
rect 41462 419930 41522 420308
rect 42425 419930 42491 419933
rect 41462 419928 42491 419930
rect 41462 419900 42430 419928
rect 41492 419872 42430 419900
rect 42486 419872 42491 419928
rect 41492 419870 42491 419872
rect 42425 419867 42491 419870
rect 43989 419522 44055 419525
rect 41492 419520 44055 419522
rect 41492 419464 43994 419520
rect 44050 419464 44055 419520
rect 41492 419462 44055 419464
rect 43989 419459 44055 419462
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 40718 418508 40724 418572
rect 40788 418570 40794 418572
rect 41965 418570 42031 418573
rect 40788 418568 42031 418570
rect 40788 418512 41970 418568
rect 42026 418512 42031 418568
rect 40788 418510 42031 418512
rect 40788 418508 40794 418510
rect 41965 418507 42031 418510
rect 40534 418236 40540 418300
rect 40604 418298 40610 418300
rect 41781 418298 41847 418301
rect 40604 418296 41847 418298
rect 40604 418240 41786 418296
rect 41842 418240 41847 418296
rect 40604 418238 41847 418240
rect 40604 418236 40610 418238
rect 41781 418235 41847 418238
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 43253 407826 43319 407829
rect 42425 407824 43319 407826
rect 42425 407768 42430 407824
rect 42486 407768 43258 407824
rect 43314 407768 43319 407824
rect 42425 407766 43319 407768
rect 42425 407763 42491 407766
rect 43253 407763 43319 407766
rect 42425 407010 42491 407013
rect 44633 407010 44699 407013
rect 42425 407008 44699 407010
rect 42425 406952 42430 407008
rect 42486 406952 44638 407008
rect 44694 406952 44699 407008
rect 42425 406950 44699 406952
rect 42425 406947 42491 406950
rect 44633 406947 44699 406950
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 42609 405650 42675 405653
rect 45369 405650 45435 405653
rect 42609 405648 45435 405650
rect 42609 405592 42614 405648
rect 42670 405592 45374 405648
rect 45430 405592 45435 405648
rect 42609 405590 45435 405592
rect 42609 405587 42675 405590
rect 45369 405587 45435 405590
rect 660297 405650 660363 405653
rect 676029 405650 676095 405653
rect 660297 405648 676095 405650
rect 660297 405592 660302 405648
rect 660358 405592 676034 405648
rect 676090 405592 676095 405648
rect 660297 405590 676095 405592
rect 660297 405587 660363 405590
rect 676029 405587 676095 405590
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669957 403746 670023 403749
rect 676262 403746 676322 403852
rect 669957 403744 676322 403746
rect 669957 403688 669962 403744
rect 670018 403688 676322 403744
rect 669957 403686 676322 403688
rect 669957 403683 670023 403686
rect 676029 403474 676095 403477
rect 676029 403472 676292 403474
rect 676029 403416 676034 403472
rect 676090 403416 676292 403472
rect 676029 403414 676292 403416
rect 676029 403411 676095 403414
rect 683113 403338 683179 403341
rect 683070 403336 683179 403338
rect 683070 403280 683118 403336
rect 683174 403280 683179 403336
rect 683070 403275 683179 403280
rect 683070 403036 683130 403275
rect 42333 402930 42399 402933
rect 43069 402930 43135 402933
rect 42333 402928 43135 402930
rect 42333 402872 42338 402928
rect 42394 402872 43074 402928
rect 43130 402872 43135 402928
rect 42333 402870 43135 402872
rect 42333 402867 42399 402870
rect 43069 402867 43135 402870
rect 676990 402868 676996 402932
rect 677060 402868 677066 402932
rect 676998 402628 677058 402868
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674649 402250 674715 402253
rect 674649 402248 676292 402250
rect 674649 402192 674654 402248
rect 674710 402192 676292 402248
rect 674649 402190 676292 402192
rect 674649 402187 674715 402190
rect 41781 401844 41847 401845
rect 41781 401840 41828 401844
rect 41892 401842 41898 401844
rect 41781 401784 41786 401840
rect 41781 401780 41828 401784
rect 41892 401782 41938 401842
rect 41892 401780 41898 401782
rect 41781 401779 41847 401780
rect 672441 401706 672507 401709
rect 676262 401706 676322 401812
rect 672441 401704 676322 401706
rect 672441 401648 672446 401704
rect 672502 401648 676322 401704
rect 672441 401646 676322 401648
rect 672441 401643 672507 401646
rect 674189 401434 674255 401437
rect 674189 401432 676292 401434
rect 674189 401376 674194 401432
rect 674250 401376 676292 401432
rect 674189 401374 676292 401376
rect 674189 401371 674255 401374
rect 676806 401236 676812 401300
rect 676876 401236 676882 401300
rect 676814 400996 676874 401236
rect 672441 400482 672507 400485
rect 676262 400482 676322 400588
rect 672441 400480 676322 400482
rect 672441 400424 672446 400480
rect 672502 400424 676322 400480
rect 672441 400422 676322 400424
rect 672441 400419 672507 400422
rect 42425 400210 42491 400213
rect 47117 400210 47183 400213
rect 42425 400208 47183 400210
rect 42425 400152 42430 400208
rect 42486 400152 47122 400208
rect 47178 400152 47183 400208
rect 42425 400150 47183 400152
rect 42425 400147 42491 400150
rect 47117 400147 47183 400150
rect 672625 400074 672691 400077
rect 676262 400074 676322 400180
rect 672625 400072 676322 400074
rect 672625 400016 672630 400072
rect 672686 400016 676322 400072
rect 672625 400014 676322 400016
rect 672625 400011 672691 400014
rect 42425 399802 42491 399805
rect 46933 399802 46999 399805
rect 42425 399800 46999 399802
rect 42425 399744 42430 399800
rect 42486 399744 46938 399800
rect 46994 399744 46999 399800
rect 42425 399742 46999 399744
rect 42425 399739 42491 399742
rect 46933 399739 46999 399742
rect 676262 399666 676322 399772
rect 674790 399606 676322 399666
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 673177 398850 673243 398853
rect 674790 398850 674850 399606
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 673177 398848 674850 398850
rect 673177 398792 673182 398848
rect 673238 398792 674850 398848
rect 673177 398790 674850 398792
rect 673177 398787 673243 398790
rect 675886 398788 675892 398852
rect 675956 398850 675962 398852
rect 676262 398850 676322 398956
rect 675956 398790 676322 398850
rect 675956 398788 675962 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 672993 397218 673059 397221
rect 676262 397218 676322 397324
rect 672993 397216 676322 397218
rect 672993 397160 672998 397216
rect 673054 397160 676322 397216
rect 672993 397158 676322 397160
rect 672993 397155 673059 397158
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 673361 396402 673427 396405
rect 676262 396402 676322 396508
rect 673361 396400 676322 396402
rect 673361 396344 673366 396400
rect 673422 396344 676322 396400
rect 673361 396342 676322 396344
rect 673361 396339 673427 396342
rect 673821 396130 673887 396133
rect 673821 396128 676292 396130
rect 673821 396072 673826 396128
rect 673882 396072 676292 396128
rect 673821 396070 676292 396072
rect 673821 396067 673887 396070
rect 674005 395722 674071 395725
rect 674005 395720 676292 395722
rect 674005 395664 674010 395720
rect 674066 395664 676292 395720
rect 674005 395662 676292 395664
rect 674005 395659 674071 395662
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 674465 394498 674531 394501
rect 674465 394496 676292 394498
rect 674465 394440 674470 394496
rect 674526 394440 676292 394496
rect 674465 394438 676292 394440
rect 674465 394435 674531 394438
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 670601 393546 670667 393549
rect 676262 393546 676322 393652
rect 670601 393544 676322 393546
rect 670601 393488 670606 393544
rect 670662 393488 676322 393544
rect 670601 393486 676322 393488
rect 670601 393483 670667 393486
rect 676070 393076 676076 393140
rect 676140 393138 676146 393140
rect 676262 393138 676322 393244
rect 676140 393078 676322 393138
rect 676140 393076 676146 393078
rect 676262 392836 676322 393078
rect 672809 392594 672875 392597
rect 672809 392592 676322 392594
rect 672809 392536 672814 392592
rect 672870 392536 676322 392592
rect 672809 392534 676322 392536
rect 672809 392531 672875 392534
rect 676262 392428 676322 392534
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 41492 387638 51090 387698
rect 41492 387230 49250 387290
rect 41137 387154 41203 387157
rect 41094 387152 41203 387154
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387091 41203 387096
rect 41094 386852 41154 387091
rect 41873 387018 41939 387021
rect 48957 387018 49023 387021
rect 41873 387016 49023 387018
rect 41873 386960 41878 387016
rect 41934 386960 48962 387016
rect 49018 386960 49023 387016
rect 41873 386958 49023 386960
rect 41873 386955 41939 386958
rect 48957 386955 49023 386958
rect 41321 386746 41387 386749
rect 41278 386744 41387 386746
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386683 41387 386688
rect 41505 386746 41571 386749
rect 45001 386746 45067 386749
rect 41505 386744 45067 386746
rect 41505 386688 41510 386744
rect 41566 386688 45006 386744
rect 45062 386688 45067 386744
rect 41505 386686 45067 386688
rect 41505 386683 41571 386686
rect 45001 386683 45067 386686
rect 41278 386444 41338 386683
rect 49190 386474 49250 387230
rect 51030 386746 51090 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 51717 386746 51783 386749
rect 51030 386744 51783 386746
rect 51030 386688 51722 386744
rect 51778 386688 51783 386744
rect 51030 386686 51783 386688
rect 51717 386683 51783 386686
rect 51901 386474 51967 386477
rect 49190 386472 51967 386474
rect 49190 386416 51906 386472
rect 51962 386416 51967 386472
rect 49190 386414 51967 386416
rect 51901 386411 51967 386414
rect 45369 386066 45435 386069
rect 41492 386064 45435 386066
rect 41492 386008 45374 386064
rect 45430 386008 45435 386064
rect 41492 386006 45435 386008
rect 45369 386003 45435 386006
rect 44173 385658 44239 385661
rect 41492 385656 44239 385658
rect 41492 385600 44178 385656
rect 44234 385600 44239 385656
rect 41492 385598 44239 385600
rect 44173 385595 44239 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 675753 384978 675819 384981
rect 676254 384978 676260 384980
rect 675753 384976 676260 384978
rect 675753 384920 675758 384976
rect 675814 384920 676260 384976
rect 675753 384918 676260 384920
rect 675753 384915 675819 384918
rect 676254 384916 676260 384918
rect 676324 384916 676330 384980
rect 45185 384842 45251 384845
rect 41492 384840 45251 384842
rect 41492 384784 45190 384840
rect 45246 384784 45251 384840
rect 41492 384782 45251 384784
rect 45185 384779 45251 384782
rect 45001 384434 45067 384437
rect 41492 384432 45067 384434
rect 41492 384376 45006 384432
rect 45062 384376 45067 384432
rect 41492 384374 45067 384376
rect 45001 384371 45067 384374
rect 44449 384026 44515 384029
rect 41492 384024 44515 384026
rect 41492 383968 44454 384024
rect 44510 383968 44515 384024
rect 41492 383966 44515 383968
rect 44449 383963 44515 383966
rect 45185 383618 45251 383621
rect 41492 383616 45251 383618
rect 41492 383560 45190 383616
rect 45246 383560 45251 383616
rect 41492 383558 45251 383560
rect 45185 383555 45251 383558
rect 45553 383210 45619 383213
rect 41492 383208 45619 383210
rect 41492 383152 45558 383208
rect 45614 383152 45619 383208
rect 41492 383150 45619 383152
rect 45553 383147 45619 383150
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 673361 382258 673427 382261
rect 675385 382258 675451 382261
rect 673361 382256 675451 382258
rect 673361 382200 673366 382256
rect 673422 382200 675390 382256
rect 675446 382200 675451 382256
rect 673361 382198 675451 382200
rect 673361 382195 673427 382198
rect 675385 382195 675451 382198
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 37966 381445 38026 381548
rect 37917 381440 38026 381445
rect 37917 381384 37922 381440
rect 37978 381384 38026 381440
rect 37917 381382 38026 381384
rect 673821 381442 673887 381445
rect 675109 381442 675175 381445
rect 673821 381440 675175 381442
rect 673821 381384 673826 381440
rect 673882 381384 675114 381440
rect 675170 381384 675175 381440
rect 673821 381382 675175 381384
rect 37917 381379 37983 381382
rect 673821 381379 673887 381382
rect 675109 381379 675175 381382
rect 40174 381037 40234 381140
rect 40174 381032 40283 381037
rect 40174 380976 40222 381032
rect 40278 380976 40283 381032
rect 40174 380974 40283 380976
rect 40217 380971 40283 380974
rect 46933 380762 46999 380765
rect 41492 380760 46999 380762
rect 41492 380704 46938 380760
rect 46994 380704 46999 380760
rect 41492 380702 46999 380704
rect 46933 380699 46999 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 33734 380221 33794 380324
rect 33734 380216 33843 380221
rect 33734 380160 33782 380216
rect 33838 380160 33843 380216
rect 33734 380158 33843 380160
rect 33777 380155 33843 380158
rect 47117 379946 47183 379949
rect 41492 379944 47183 379946
rect 41492 379888 47122 379944
rect 47178 379888 47183 379944
rect 41492 379886 47183 379888
rect 47117 379883 47183 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 45737 379130 45803 379133
rect 41492 379128 45803 379130
rect 41492 379072 45742 379128
rect 45798 379072 45803 379128
rect 41492 379070 45803 379072
rect 45737 379067 45803 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 652017 378178 652083 378181
rect 650164 378176 652083 378178
rect 650164 378120 652022 378176
rect 652078 378120 652083 378176
rect 650164 378118 652083 378120
rect 652017 378115 652083 378118
rect 672993 378042 673059 378045
rect 674782 378042 674788 378044
rect 672993 378040 674788 378042
rect 672993 377984 672998 378040
rect 673054 377984 674788 378040
rect 672993 377982 674788 377984
rect 672993 377979 673059 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 44449 377906 44515 377909
rect 41492 377904 44515 377906
rect 41492 377848 44454 377904
rect 44510 377848 44515 377904
rect 41492 377846 44515 377848
rect 44449 377843 44515 377846
rect 674465 377770 674531 377773
rect 675109 377770 675175 377773
rect 674465 377768 675175 377770
rect 674465 377712 674470 377768
rect 674526 377712 675114 377768
rect 675170 377712 675175 377768
rect 674465 377710 675175 377712
rect 674465 377707 674531 377710
rect 675109 377707 675175 377710
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675201 377498 675267 377501
rect 675886 377498 675892 377500
rect 675201 377496 675892 377498
rect 675201 377440 675206 377496
rect 675262 377440 675892 377496
rect 675201 377438 675892 377440
rect 675201 377435 675267 377438
rect 675886 377436 675892 377438
rect 675956 377436 675962 377500
rect 675753 377226 675819 377229
rect 676622 377226 676628 377228
rect 675753 377224 676628 377226
rect 675753 377168 675758 377224
rect 675814 377168 676628 377224
rect 675753 377166 676628 377168
rect 675753 377163 675819 377166
rect 676622 377164 676628 377166
rect 676692 377164 676698 377228
rect 27662 376546 27722 377060
rect 40033 376954 40099 376957
rect 41638 376954 41644 376956
rect 40033 376952 41644 376954
rect 40033 376896 40038 376952
rect 40094 376896 41644 376952
rect 40033 376894 41644 376896
rect 40033 376891 40099 376894
rect 41638 376892 41644 376894
rect 41708 376892 41714 376956
rect 28533 376546 28599 376549
rect 27662 376544 28599 376546
rect 27662 376488 28538 376544
rect 28594 376488 28599 376544
rect 27662 376486 28599 376488
rect 28533 376483 28599 376486
rect 62113 376274 62179 376277
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 62113 376272 64492 376274
rect 35758 376141 35818 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 62113 376211 62179 376214
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 35758 376136 35867 376141
rect 35758 376080 35806 376136
rect 35862 376080 35867 376136
rect 35758 376078 35867 376080
rect 35801 376075 35867 376078
rect 41689 375458 41755 375461
rect 43345 375458 43411 375461
rect 41689 375456 43411 375458
rect 41689 375400 41694 375456
rect 41750 375400 43350 375456
rect 43406 375400 43411 375456
rect 41689 375398 43411 375400
rect 41689 375395 41755 375398
rect 43345 375395 43411 375398
rect 674005 375458 674071 375461
rect 675385 375458 675451 375461
rect 674005 375456 675451 375458
rect 674005 375400 674010 375456
rect 674066 375400 675390 375456
rect 675446 375400 675451 375456
rect 674005 375398 675451 375400
rect 674005 375395 674071 375398
rect 675385 375395 675451 375398
rect 28533 373282 28599 373285
rect 41270 373282 41276 373284
rect 28533 373280 41276 373282
rect 28533 373224 28538 373280
rect 28594 373224 41276 373280
rect 28533 373222 41276 373224
rect 28533 373219 28599 373222
rect 41270 373220 41276 373222
rect 41340 373220 41346 373284
rect 41689 373282 41755 373285
rect 42609 373282 42675 373285
rect 41689 373280 42675 373282
rect 41689 373224 41694 373280
rect 41750 373224 42614 373280
rect 42670 373224 42675 373280
rect 41689 373222 42675 373224
rect 41689 373219 41755 373222
rect 42609 373219 42675 373222
rect 675753 373010 675819 373013
rect 676070 373010 676076 373012
rect 675753 373008 676076 373010
rect 675753 372952 675758 373008
rect 675814 372952 676076 373008
rect 675753 372950 676076 372952
rect 675753 372947 675819 372950
rect 676070 372948 676076 372950
rect 676140 372948 676146 373012
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 33777 371922 33843 371925
rect 41822 371922 41828 371924
rect 33777 371920 41828 371922
rect 33777 371864 33782 371920
rect 33838 371864 41828 371920
rect 33777 371862 41828 371864
rect 33777 371859 33843 371862
rect 41822 371860 41828 371862
rect 41892 371860 41898 371924
rect 41270 368460 41276 368524
rect 41340 368522 41346 368524
rect 41781 368522 41847 368525
rect 41340 368520 41847 368522
rect 41340 368464 41786 368520
rect 41842 368464 41847 368520
rect 41340 368462 41847 368464
rect 41340 368460 41346 368462
rect 41781 368459 41847 368462
rect 42425 367026 42491 367029
rect 46197 367026 46263 367029
rect 42425 367024 46263 367026
rect 42425 366968 42430 367024
rect 42486 366968 46202 367024
rect 46258 366968 46263 367024
rect 42425 366966 46263 366968
rect 42425 366963 42491 366966
rect 46197 366963 46263 366966
rect 42333 365802 42399 365805
rect 42793 365802 42859 365805
rect 42333 365800 42859 365802
rect 42333 365744 42338 365800
rect 42394 365744 42798 365800
rect 42854 365744 42859 365800
rect 42333 365742 42859 365744
rect 42333 365739 42399 365742
rect 42793 365739 42859 365742
rect 42149 364986 42215 364989
rect 44449 364986 44515 364989
rect 42149 364984 44515 364986
rect 42149 364928 42154 364984
rect 42210 364928 44454 364984
rect 44510 364928 44515 364984
rect 42149 364926 44515 364928
rect 42149 364923 42215 364926
rect 44449 364923 44515 364926
rect 651649 364850 651715 364853
rect 650164 364848 651715 364850
rect 650164 364792 651654 364848
rect 651710 364792 651715 364848
rect 650164 364790 651715 364792
rect 651649 364787 651715 364790
rect 42425 364306 42491 364309
rect 45737 364306 45803 364309
rect 42425 364304 45803 364306
rect 42425 364248 42430 364304
rect 42486 364248 45742 364304
rect 45798 364248 45803 364304
rect 42425 364246 45803 364248
rect 42425 364243 42491 364246
rect 45737 364243 45803 364246
rect 40718 363564 40724 363628
rect 40788 363626 40794 363628
rect 41781 363626 41847 363629
rect 40788 363624 41847 363626
rect 40788 363568 41786 363624
rect 41842 363568 41847 363624
rect 40788 363566 41847 363568
rect 40788 363564 40794 363566
rect 41781 363563 41847 363566
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 668761 360906 668827 360909
rect 675845 360906 675911 360909
rect 668761 360904 675911 360906
rect 668761 360848 668766 360904
rect 668822 360848 675850 360904
rect 675906 360848 675911 360904
rect 668761 360846 675911 360848
rect 668761 360843 668827 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 41781 359412 41847 359413
rect 41781 359408 41828 359412
rect 41892 359410 41898 359412
rect 41781 359352 41786 359408
rect 41781 359348 41828 359352
rect 41892 359350 41938 359410
rect 41892 359348 41898 359350
rect 41781 359347 41847 359348
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 665817 358730 665883 358733
rect 665817 358728 676292 358730
rect 665817 358672 665822 358728
rect 665878 358672 676292 358728
rect 665817 358670 676292 358672
rect 665817 358667 665883 358670
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 674649 357506 674715 357509
rect 674649 357504 676292 357506
rect 674649 357448 674654 357504
rect 674710 357448 676292 357504
rect 674649 357446 676292 357448
rect 674649 357443 674715 357446
rect 42425 357370 42491 357373
rect 47117 357370 47183 357373
rect 42425 357368 47183 357370
rect 42425 357312 42430 357368
rect 42486 357312 47122 357368
rect 47178 357312 47183 357368
rect 42425 357310 47183 357312
rect 42425 357307 42491 357310
rect 47117 357307 47183 357310
rect 674649 357098 674715 357101
rect 674649 357096 676292 357098
rect 674649 357040 674654 357096
rect 674710 357040 676292 357096
rect 674649 357038 676292 357040
rect 674649 357035 674715 357038
rect 42057 356962 42123 356965
rect 45553 356962 45619 356965
rect 42057 356960 45619 356962
rect 42057 356904 42062 356960
rect 42118 356904 45558 356960
rect 45614 356904 45619 356960
rect 42057 356902 45619 356904
rect 42057 356899 42123 356902
rect 45553 356899 45619 356902
rect 44265 356690 44331 356693
rect 45645 356690 45711 356693
rect 44265 356688 45711 356690
rect 44265 356632 44270 356688
rect 44326 356632 45650 356688
rect 45706 356632 45711 356688
rect 44265 356630 45711 356632
rect 44265 356627 44331 356630
rect 45645 356627 45711 356630
rect 674189 356690 674255 356693
rect 674189 356688 676292 356690
rect 674189 356632 674194 356688
rect 674250 356632 676292 356688
rect 674189 356630 676292 356632
rect 674189 356627 674255 356630
rect 674097 356282 674163 356285
rect 674097 356280 676292 356282
rect 674097 356224 674102 356280
rect 674158 356224 676292 356280
rect 674097 356222 676292 356224
rect 674097 356219 674163 356222
rect 42425 356146 42491 356149
rect 46933 356146 46999 356149
rect 42425 356144 46999 356146
rect 42425 356088 42430 356144
rect 42486 356088 46938 356144
rect 46994 356088 46999 356144
rect 42425 356086 46999 356088
rect 42425 356083 42491 356086
rect 46933 356083 46999 356086
rect 43345 355874 43411 355877
rect 45921 355874 45987 355877
rect 43345 355872 45987 355874
rect 43345 355816 43350 355872
rect 43406 355816 45926 355872
rect 45982 355816 45987 355872
rect 43345 355814 45987 355816
rect 43345 355811 43411 355814
rect 45921 355811 45987 355814
rect 672441 355874 672507 355877
rect 672441 355872 676292 355874
rect 672441 355816 672446 355872
rect 672502 355816 676292 355872
rect 672441 355814 676292 355816
rect 672441 355811 672507 355814
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 672441 355466 672507 355469
rect 672441 355464 676292 355466
rect 672441 355408 672446 355464
rect 672502 355408 676292 355464
rect 672441 355406 676292 355408
rect 672441 355403 672507 355406
rect 673177 355058 673243 355061
rect 673177 355056 676292 355058
rect 673177 355000 673182 355056
rect 673238 355000 676292 355056
rect 673177 354998 676292 355000
rect 673177 354995 673243 354998
rect 672993 354650 673059 354653
rect 672993 354648 676292 354650
rect 672993 354592 672998 354648
rect 673054 354592 676292 354648
rect 672993 354590 676292 354592
rect 672993 354587 673059 354590
rect 43897 354244 43963 354245
rect 43846 354180 43852 354244
rect 43916 354242 43963 354244
rect 43916 354240 44008 354242
rect 43958 354184 44008 354240
rect 43916 354182 44008 354184
rect 43916 354180 43963 354182
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 43897 354179 43963 354180
rect 44214 353772 44220 353836
rect 44284 353834 44290 353836
rect 44725 353834 44791 353837
rect 44284 353832 44791 353834
rect 44284 353776 44730 353832
rect 44786 353776 44791 353832
rect 44284 353774 44791 353776
rect 44284 353772 44290 353774
rect 44725 353771 44791 353774
rect 676029 353834 676095 353837
rect 676029 353832 676292 353834
rect 676029 353776 676034 353832
rect 676090 353776 676292 353832
rect 676029 353774 676292 353776
rect 676029 353771 676095 353774
rect 673177 353426 673243 353429
rect 673177 353424 676292 353426
rect 673177 353368 673182 353424
rect 673238 353368 676292 353424
rect 673177 353366 676292 353368
rect 673177 353363 673243 353366
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 673913 352610 673979 352613
rect 673913 352608 676292 352610
rect 673913 352552 673918 352608
rect 673974 352552 676292 352608
rect 673913 352550 676292 352552
rect 673913 352547 673979 352550
rect 673545 352202 673611 352205
rect 673545 352200 676292 352202
rect 673545 352144 673550 352200
rect 673606 352144 676292 352200
rect 673545 352142 676292 352144
rect 673545 352139 673611 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 651465 351658 651531 351661
rect 650164 351656 651531 351658
rect 650164 351600 651470 351656
rect 651526 351600 651531 351656
rect 650164 351598 651531 351600
rect 651465 351595 651531 351598
rect 672257 351386 672323 351389
rect 672257 351384 676292 351386
rect 672257 351328 672262 351384
rect 672318 351328 676292 351384
rect 672257 351326 676292 351328
rect 672257 351323 672323 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 673729 350570 673795 350573
rect 673729 350568 676292 350570
rect 673729 350512 673734 350568
rect 673790 350512 676292 350568
rect 673729 350510 676292 350512
rect 673729 350507 673795 350510
rect 62757 350298 62823 350301
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 62757 350235 62823 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 673361 349754 673427 349757
rect 673361 349752 676292 349754
rect 673361 349696 673366 349752
rect 673422 349696 676292 349752
rect 673361 349694 676292 349696
rect 673361 349691 673427 349694
rect 674465 349482 674531 349485
rect 674465 349480 676230 349482
rect 674465 349424 674470 349480
rect 674526 349424 676230 349480
rect 674465 349422 676230 349424
rect 674465 349419 674531 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 675937 349212 676003 349213
rect 675886 349210 675892 349212
rect 675846 349150 675892 349210
rect 675956 349208 676003 349212
rect 675998 349152 676003 349208
rect 675886 349148 675892 349150
rect 675956 349148 676003 349152
rect 675937 349147 676003 349148
rect 671981 348938 672047 348941
rect 671981 348936 676292 348938
rect 671981 348880 671986 348936
rect 672042 348880 676292 348936
rect 671981 348878 676292 348880
rect 671981 348875 672047 348878
rect 672625 348530 672691 348533
rect 672625 348528 676292 348530
rect 672625 348472 672630 348528
rect 672686 348472 676292 348528
rect 672625 348470 676292 348472
rect 672625 348467 672691 348470
rect 674281 347714 674347 347717
rect 683070 347714 683130 348092
rect 674281 347712 683130 347714
rect 674281 347656 674286 347712
rect 674342 347684 683130 347712
rect 674342 347656 683100 347684
rect 674281 347654 683100 347656
rect 674281 347651 674347 347654
rect 669957 347306 670023 347309
rect 669957 347304 676292 347306
rect 669957 347248 669962 347304
rect 670018 347248 676292 347304
rect 669957 347246 676292 347248
rect 669957 347243 670023 347246
rect 38285 346354 38351 346357
rect 49141 346354 49207 346357
rect 38285 346352 49207 346354
rect 38285 346296 38290 346352
rect 38346 346296 49146 346352
rect 49202 346296 49207 346352
rect 38285 346294 49207 346296
rect 38285 346291 38351 346294
rect 49141 346291 49207 346294
rect 28901 344314 28967 344317
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 28901 344312 29010 344314
rect 28901 344256 28906 344312
rect 28962 344256 29010 344312
rect 28901 344251 29010 344256
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 28950 344148 29010 344251
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 28582 343740 28642 343843
rect 45369 343362 45435 343365
rect 41492 343360 45435 343362
rect 41492 343304 45374 343360
rect 45430 343304 45435 343360
rect 41492 343302 45435 343304
rect 45369 343299 45435 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 44214 342546 44220 342548
rect 41492 342486 44220 342546
rect 44214 342484 44220 342486
rect 44284 342484 44290 342548
rect 44582 342138 44588 342140
rect 41492 342078 44588 342138
rect 44582 342076 44588 342078
rect 44652 342076 44658 342140
rect 45001 341730 45067 341733
rect 41492 341728 45067 341730
rect 41492 341672 45006 341728
rect 45062 341672 45067 341728
rect 41492 341670 45067 341672
rect 45001 341667 45067 341670
rect 44398 341322 44404 341324
rect 41492 341262 44404 341322
rect 44398 341260 44404 341262
rect 44468 341260 44474 341324
rect 45185 340914 45251 340917
rect 41492 340912 45251 340914
rect 41492 340856 45190 340912
rect 45246 340856 45251 340912
rect 41492 340854 45251 340856
rect 45185 340851 45251 340854
rect 673177 340778 673243 340781
rect 675109 340778 675175 340781
rect 673177 340776 675175 340778
rect 673177 340720 673182 340776
rect 673238 340720 675114 340776
rect 675170 340720 675175 340776
rect 673177 340718 675175 340720
rect 673177 340715 673243 340718
rect 675109 340715 675175 340718
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340370 675819 340373
rect 676622 340370 676628 340372
rect 675753 340368 676628 340370
rect 675753 340312 675758 340368
rect 675814 340312 676628 340368
rect 675753 340310 676628 340312
rect 675753 340307 675819 340310
rect 676622 340308 676628 340310
rect 676692 340308 676698 340372
rect 46933 340098 46999 340101
rect 41492 340096 46999 340098
rect 41492 340040 46938 340096
rect 46994 340040 46999 340096
rect 41492 340038 46999 340040
rect 46933 340035 46999 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 35758 339013 35818 339252
rect 35758 339008 35867 339013
rect 675385 339012 675451 339013
rect 675334 339010 675340 339012
rect 35758 338952 35806 339008
rect 35862 338952 35867 339008
rect 35758 338950 35867 338952
rect 675294 338950 675340 339010
rect 675404 339008 675451 339012
rect 675446 338952 675451 339008
rect 35801 338947 35867 338950
rect 675334 338948 675340 338950
rect 675404 338948 675451 338952
rect 675385 338947 675451 338948
rect 30974 338605 31034 338844
rect 30974 338600 31083 338605
rect 30974 338544 31022 338600
rect 31078 338544 31083 338600
rect 30974 338542 31083 338544
rect 31017 338539 31083 338542
rect 45645 338466 45711 338469
rect 41492 338464 45711 338466
rect 41492 338408 45650 338464
rect 45706 338408 45711 338464
rect 41492 338406 45711 338408
rect 45645 338403 45711 338406
rect 651465 338330 651531 338333
rect 650164 338328 651531 338330
rect 650164 338272 651470 338328
rect 651526 338272 651531 338328
rect 650164 338270 651531 338272
rect 651465 338267 651531 338270
rect 40726 337788 40786 338028
rect 675569 337788 675635 337789
rect 40718 337724 40724 337788
rect 40788 337724 40794 337788
rect 675518 337786 675524 337788
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 42742 337650 42748 337652
rect 41492 337590 42748 337650
rect 42742 337588 42748 337590
rect 42812 337588 42818 337652
rect 45461 337242 45527 337245
rect 41492 337240 45527 337242
rect 41492 337184 45466 337240
rect 45522 337184 45527 337240
rect 41492 337182 45527 337184
rect 45461 337179 45527 337182
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 42926 336834 42932 336836
rect 41492 336774 42932 336834
rect 42926 336772 42932 336774
rect 42996 336772 43002 336836
rect 673913 336698 673979 336701
rect 675109 336698 675175 336701
rect 673913 336696 675175 336698
rect 673913 336640 673918 336696
rect 673974 336640 675114 336696
rect 675170 336640 675175 336696
rect 673913 336638 675175 336640
rect 673913 336635 673979 336638
rect 675109 336635 675175 336638
rect 675753 336698 675819 336701
rect 676438 336698 676444 336700
rect 675753 336696 676444 336698
rect 675753 336640 675758 336696
rect 675814 336640 676444 336696
rect 675753 336638 676444 336640
rect 675753 336635 675819 336638
rect 676438 336636 676444 336638
rect 676508 336636 676514 336700
rect 41462 336154 41522 336396
rect 43110 336154 43116 336156
rect 41462 336094 43116 336154
rect 43110 336092 43116 336094
rect 43180 336092 43186 336156
rect 40542 335748 40602 335988
rect 673361 335882 673427 335885
rect 675477 335882 675543 335885
rect 673361 335880 675543 335882
rect 673361 335824 673366 335880
rect 673422 335824 675482 335880
rect 675538 335824 675543 335880
rect 673361 335822 675543 335824
rect 673361 335819 673427 335822
rect 675477 335819 675543 335822
rect 40534 335684 40540 335748
rect 40604 335684 40610 335748
rect 41462 335474 41522 335580
rect 42558 335474 42564 335476
rect 41462 335414 42564 335474
rect 42558 335412 42564 335414
rect 42628 335412 42634 335476
rect 37917 335338 37983 335341
rect 41270 335338 41276 335340
rect 37917 335336 41276 335338
rect 37917 335280 37922 335336
rect 37978 335280 41276 335336
rect 37917 335278 41276 335280
rect 37917 335275 37983 335278
rect 41270 335276 41276 335278
rect 41340 335276 41346 335340
rect 672257 335338 672323 335341
rect 675293 335338 675359 335341
rect 672257 335336 675359 335338
rect 672257 335280 672262 335336
rect 672318 335280 675298 335336
rect 675354 335280 675359 335336
rect 672257 335278 675359 335280
rect 672257 335275 672323 335278
rect 675293 335275 675359 335278
rect 41462 334930 41522 335172
rect 41462 334870 43546 334930
rect 41462 334658 41522 334764
rect 41462 334598 42258 334658
rect 42198 334386 42258 334598
rect 42558 334596 42564 334660
rect 42628 334658 42634 334660
rect 42793 334658 42859 334661
rect 43161 334660 43227 334661
rect 43110 334658 43116 334660
rect 42628 334656 42859 334658
rect 42628 334600 42798 334656
rect 42854 334600 42859 334656
rect 42628 334598 42859 334600
rect 43070 334598 43116 334658
rect 43180 334656 43227 334660
rect 43222 334600 43227 334656
rect 42628 334596 42634 334598
rect 42793 334595 42859 334598
rect 43110 334596 43116 334598
rect 43180 334596 43227 334600
rect 43486 334658 43546 334870
rect 44265 334658 44331 334661
rect 43486 334656 44331 334658
rect 43486 334600 44270 334656
rect 44326 334600 44331 334656
rect 43486 334598 44331 334600
rect 43161 334595 43227 334596
rect 44265 334595 44331 334598
rect 42977 334386 43043 334389
rect 42198 334384 43043 334386
rect 41462 334114 41522 334356
rect 42198 334328 42982 334384
rect 43038 334328 43043 334384
rect 42198 334326 43043 334328
rect 42977 334323 43043 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 674465 332890 674531 332893
rect 675385 332890 675451 332893
rect 674465 332888 675451 332890
rect 674465 332832 674470 332888
rect 674526 332832 675390 332888
rect 675446 332832 675451 332888
rect 674465 332830 675451 332832
rect 674465 332827 674531 332830
rect 675385 332827 675451 332830
rect 671981 332346 672047 332349
rect 675109 332346 675175 332349
rect 671981 332344 675175 332346
rect 671981 332288 671986 332344
rect 672042 332288 675114 332344
rect 675170 332288 675175 332344
rect 671981 332286 675175 332288
rect 671981 332283 672047 332286
rect 675109 332283 675175 332286
rect 675753 332210 675819 332213
rect 676254 332210 676260 332212
rect 675753 332208 676260 332210
rect 675753 332152 675758 332208
rect 675814 332152 676260 332208
rect 675753 332150 676260 332152
rect 675753 332147 675819 332150
rect 676254 332148 676260 332150
rect 676324 332148 676330 332212
rect 673729 331122 673795 331125
rect 675109 331122 675175 331125
rect 673729 331120 675175 331122
rect 673729 331064 673734 331120
rect 673790 331064 675114 331120
rect 675170 331064 675175 331120
rect 673729 331062 675175 331064
rect 673729 331059 673795 331062
rect 675109 331059 675175 331062
rect 31017 329082 31083 329085
rect 41638 329082 41644 329084
rect 31017 329080 41644 329082
rect 31017 329024 31022 329080
rect 31078 329024 41644 329080
rect 31017 329022 41644 329024
rect 31017 329019 31083 329022
rect 41638 329020 41644 329022
rect 41708 329020 41714 329084
rect 36537 328402 36603 328405
rect 42006 328402 42012 328404
rect 36537 328400 42012 328402
rect 36537 328344 36542 328400
rect 36598 328344 42012 328400
rect 36537 328342 42012 328344
rect 36537 328339 36603 328342
rect 42006 328340 42012 328342
rect 42076 328340 42082 328404
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 674281 327586 674347 327589
rect 675109 327586 675175 327589
rect 674281 327584 675175 327586
rect 674281 327528 674286 327584
rect 674342 327528 675114 327584
rect 675170 327528 675175 327584
rect 674281 327526 675175 327528
rect 674281 327523 674347 327526
rect 675109 327523 675175 327526
rect 40718 326708 40724 326772
rect 40788 326770 40794 326772
rect 41781 326770 41847 326773
rect 40788 326768 41847 326770
rect 40788 326712 41786 326768
rect 41842 326712 41847 326768
rect 40788 326710 41847 326712
rect 40788 326708 40794 326710
rect 41781 326707 41847 326710
rect 673545 325682 673611 325685
rect 675109 325682 675175 325685
rect 673545 325680 675175 325682
rect 673545 325624 673550 325680
rect 673606 325624 675114 325680
rect 675170 325624 675175 325680
rect 673545 325622 675175 325624
rect 673545 325619 673611 325622
rect 675109 325619 675175 325622
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41454 324668 41460 324732
rect 41524 324730 41530 324732
rect 41781 324730 41847 324733
rect 41524 324728 41847 324730
rect 41524 324672 41786 324728
rect 41842 324672 41847 324728
rect 41524 324670 41847 324672
rect 41524 324668 41530 324670
rect 41781 324667 41847 324670
rect 42241 323642 42307 323645
rect 42977 323642 43043 323645
rect 42241 323640 43043 323642
rect 42241 323584 42246 323640
rect 42302 323584 42982 323640
rect 43038 323584 43043 323640
rect 42241 323582 43043 323584
rect 42241 323579 42307 323582
rect 42977 323579 43043 323582
rect 43437 322962 43503 322965
rect 64462 322962 64522 324156
rect 43437 322960 64522 322962
rect 43437 322904 43442 322960
rect 43498 322904 64522 322960
rect 43437 322902 64522 322904
rect 43437 322899 43503 322902
rect 42057 322826 42123 322829
rect 43161 322826 43227 322829
rect 42057 322824 43227 322826
rect 42057 322768 42062 322824
rect 42118 322768 43166 322824
rect 43222 322768 43227 322824
rect 42057 322766 43227 322768
rect 42057 322763 42123 322766
rect 43161 322763 43227 322766
rect 42425 321466 42491 321469
rect 53097 321466 53163 321469
rect 42425 321464 53163 321466
rect 42425 321408 42430 321464
rect 42486 321408 53102 321464
rect 53158 321408 53163 321464
rect 42425 321406 53163 321408
rect 42425 321403 42491 321406
rect 53097 321403 53163 321406
rect 40534 321132 40540 321196
rect 40604 321194 40610 321196
rect 41781 321194 41847 321197
rect 40604 321192 41847 321194
rect 40604 321136 41786 321192
rect 41842 321136 41847 321192
rect 40604 321134 41847 321136
rect 40604 321132 40610 321134
rect 41781 321131 41847 321134
rect 42425 320106 42491 320109
rect 44265 320106 44331 320109
rect 42425 320104 44331 320106
rect 42425 320048 42430 320104
rect 42486 320048 44270 320104
rect 44326 320048 44331 320104
rect 42425 320046 44331 320048
rect 42425 320043 42491 320046
rect 44265 320043 44331 320046
rect 42425 318882 42491 318885
rect 45645 318882 45711 318885
rect 42425 318880 45711 318882
rect 42425 318824 42430 318880
rect 42486 318824 45650 318880
rect 45706 318824 45711 318880
rect 42425 318822 45711 318824
rect 42425 318819 42491 318822
rect 45645 318819 45711 318822
rect 42425 316434 42491 316437
rect 43110 316434 43116 316436
rect 42425 316432 43116 316434
rect 42425 316376 42430 316432
rect 42486 316376 43116 316432
rect 42425 316374 43116 316376
rect 42425 316371 42491 316374
rect 43110 316372 43116 316374
rect 43180 316372 43186 316436
rect 42149 316026 42215 316029
rect 45461 316026 45527 316029
rect 42149 316024 45527 316026
rect 42149 315968 42154 316024
rect 42210 315968 45466 316024
rect 45522 315968 45527 316024
rect 42149 315966 45527 315968
rect 42149 315963 42215 315966
rect 45461 315963 45527 315966
rect 41873 315620 41939 315621
rect 41822 315618 41828 315620
rect 41782 315558 41828 315618
rect 41892 315616 41939 315620
rect 41934 315560 41939 315616
rect 41822 315556 41828 315558
rect 41892 315556 41939 315560
rect 41873 315555 41939 315556
rect 663057 315482 663123 315485
rect 676029 315482 676095 315485
rect 663057 315480 676095 315482
rect 663057 315424 663062 315480
rect 663118 315424 676034 315480
rect 676090 315424 676095 315480
rect 663057 315422 676095 315424
rect 663057 315419 663123 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 46933 313714 46999 313717
rect 42149 313712 46999 313714
rect 42149 313656 42154 313712
rect 42210 313656 46938 313712
rect 46994 313656 46999 313712
rect 42149 313654 46999 313656
rect 42149 313651 42215 313654
rect 46933 313651 46999 313654
rect 667197 313714 667263 313717
rect 667197 313712 676292 313714
rect 667197 313656 667202 313712
rect 667258 313656 676292 313712
rect 667197 313654 676292 313656
rect 667197 313651 667263 313654
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 668577 312898 668643 312901
rect 668577 312896 676292 312898
rect 668577 312840 668582 312896
rect 668638 312840 676292 312896
rect 668577 312838 676292 312840
rect 668577 312835 668643 312838
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 42057 312628 42123 312629
rect 42006 312626 42012 312628
rect 41966 312566 42012 312626
rect 42076 312624 42123 312628
rect 42118 312568 42123 312624
rect 42006 312564 42012 312566
rect 42076 312564 42123 312568
rect 42057 312563 42123 312564
rect 674649 312490 674715 312493
rect 674649 312488 676292 312490
rect 674649 312432 674654 312488
rect 674710 312432 676292 312488
rect 674649 312430 676292 312432
rect 674649 312427 674715 312430
rect 673913 312082 673979 312085
rect 673913 312080 676292 312082
rect 673913 312024 673918 312080
rect 673974 312024 676292 312080
rect 673913 312022 676292 312024
rect 673913 312019 673979 312022
rect 651465 311810 651531 311813
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 651465 311747 651531 311750
rect 674097 311674 674163 311677
rect 674097 311672 676292 311674
rect 674097 311616 674102 311672
rect 674158 311616 676292 311672
rect 674097 311614 676292 311616
rect 674097 311611 674163 311614
rect 44214 311476 44220 311540
rect 44284 311538 44290 311540
rect 44725 311538 44791 311541
rect 44284 311536 44791 311538
rect 44284 311480 44730 311536
rect 44786 311480 44791 311536
rect 44284 311478 44791 311480
rect 44284 311476 44290 311478
rect 44725 311475 44791 311478
rect 44357 311268 44423 311269
rect 44357 311266 44404 311268
rect 44312 311264 44404 311266
rect 44312 311208 44362 311264
rect 44312 311206 44404 311208
rect 44357 311204 44404 311206
rect 44468 311204 44474 311268
rect 673177 311266 673243 311269
rect 673177 311264 676292 311266
rect 673177 311208 673182 311264
rect 673238 311208 676292 311264
rect 673177 311206 676292 311208
rect 44357 311203 44423 311204
rect 673177 311203 673243 311206
rect 44541 311132 44607 311133
rect 44541 311128 44588 311132
rect 44652 311130 44658 311132
rect 62113 311130 62179 311133
rect 44541 311072 44546 311128
rect 44541 311068 44588 311072
rect 44652 311070 44698 311130
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 44652 311068 44658 311070
rect 44541 311067 44607 311068
rect 62113 311067 62179 311070
rect 672441 310858 672507 310861
rect 672441 310856 676292 310858
rect 672441 310800 672446 310856
rect 672502 310800 676292 310856
rect 672441 310798 676292 310800
rect 672441 310795 672507 310798
rect 674465 310450 674531 310453
rect 674465 310448 676292 310450
rect 674465 310392 674470 310448
rect 674526 310392 676292 310448
rect 674465 310390 676292 310392
rect 674465 310387 674531 310390
rect 672993 310042 673059 310045
rect 672993 310040 676292 310042
rect 672993 309984 672998 310040
rect 673054 309984 676292 310040
rect 672993 309982 676292 309984
rect 672993 309979 673059 309982
rect 674189 309634 674255 309637
rect 674189 309632 676292 309634
rect 674189 309576 674194 309632
rect 674250 309576 676292 309632
rect 674189 309574 676292 309576
rect 674189 309571 674255 309574
rect 674833 309226 674899 309229
rect 674833 309224 676292 309226
rect 674833 309168 674838 309224
rect 674894 309168 676292 309224
rect 674833 309166 676292 309168
rect 674833 309163 674899 309166
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675017 308002 675083 308005
rect 675017 308000 676292 308002
rect 675017 307944 675022 308000
rect 675078 307944 676292 308000
rect 675017 307942 676292 307944
rect 675017 307939 675083 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 675886 306716 675892 306780
rect 675956 306778 675962 306780
rect 675956 306718 676292 306778
rect 675956 306716 675962 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 676397 305962 676463 305965
rect 676397 305960 676476 305962
rect 676397 305904 676402 305960
rect 676458 305904 676476 305960
rect 676397 305902 676476 305904
rect 676397 305899 676463 305902
rect 673729 305554 673795 305557
rect 673729 305552 676292 305554
rect 673729 305496 673734 305552
rect 673790 305496 676292 305552
rect 673729 305494 676292 305496
rect 673729 305491 673795 305494
rect 676673 305146 676739 305149
rect 676660 305144 676739 305146
rect 676660 305088 676678 305144
rect 676734 305088 676739 305144
rect 676660 305086 676739 305088
rect 676673 305083 676739 305086
rect 673361 304738 673427 304741
rect 673361 304736 676292 304738
rect 673361 304680 673366 304736
rect 673422 304680 676292 304736
rect 673361 304678 676292 304680
rect 673361 304675 673427 304678
rect 672993 304330 673059 304333
rect 672993 304328 676292 304330
rect 672993 304272 672998 304328
rect 673054 304272 676292 304328
rect 672993 304270 676292 304272
rect 672993 304267 673059 304270
rect 674649 303922 674715 303925
rect 674649 303920 676292 303922
rect 674649 303864 674654 303920
rect 674710 303864 676292 303920
rect 674649 303862 676292 303864
rect 674649 303859 674715 303862
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 41781 303106 41847 303109
rect 46381 303106 46447 303109
rect 41781 303104 46447 303106
rect 41781 303048 41786 303104
rect 41842 303048 46386 303104
rect 46442 303048 46447 303104
rect 41781 303046 46447 303048
rect 41781 303043 41847 303046
rect 46381 303043 46447 303046
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 668301 302290 668367 302293
rect 668301 302288 676292 302290
rect 668301 302232 668306 302288
rect 668362 302232 676292 302288
rect 668301 302230 676292 302232
rect 668301 302227 668367 302230
rect 671981 302018 672047 302021
rect 676029 302018 676095 302021
rect 671981 302016 676095 302018
rect 671981 301960 671986 302016
rect 672042 301960 676034 302016
rect 676090 301960 676095 302016
rect 671981 301958 676095 301960
rect 671981 301955 672047 301958
rect 676029 301955 676095 301958
rect 676397 301612 676463 301613
rect 676397 301608 676444 301612
rect 676508 301610 676514 301612
rect 676397 301552 676402 301608
rect 676397 301548 676444 301552
rect 676508 301550 676554 301610
rect 676508 301548 676514 301550
rect 676397 301547 676463 301548
rect 676673 301476 676739 301477
rect 676622 301412 676628 301476
rect 676692 301474 676739 301476
rect 676692 301472 676784 301474
rect 676734 301416 676784 301472
rect 676692 301414 676784 301416
rect 676692 301412 676739 301414
rect 676673 301411 676739 301412
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44725 300114 44791 300117
rect 41492 300112 44791 300114
rect 41492 300056 44730 300112
rect 44786 300056 44791 300112
rect 41492 300054 44791 300056
rect 44725 300051 44791 300054
rect 42885 299706 42951 299709
rect 41492 299704 42951 299706
rect 41492 299648 42890 299704
rect 42946 299648 42951 299704
rect 41492 299646 42951 299648
rect 42885 299643 42951 299646
rect 44541 299298 44607 299301
rect 41492 299296 44607 299298
rect 41492 299240 44546 299296
rect 44602 299240 44607 299296
rect 41492 299238 44607 299240
rect 44541 299235 44607 299238
rect 43253 298890 43319 298893
rect 41492 298888 43319 298890
rect 41492 298832 43258 298888
rect 43314 298832 43319 298888
rect 41492 298830 43319 298832
rect 43253 298827 43319 298830
rect 44357 298482 44423 298485
rect 652201 298482 652267 298485
rect 41492 298480 44423 298482
rect 41492 298424 44362 298480
rect 44418 298424 44423 298480
rect 41492 298422 44423 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 44357 298419 44423 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 44173 298074 44239 298077
rect 41492 298072 44239 298074
rect 41492 298016 44178 298072
rect 44234 298016 44239 298072
rect 41492 298014 44239 298016
rect 44173 298011 44239 298014
rect 674833 298074 674899 298077
rect 675293 298074 675359 298077
rect 674833 298072 675359 298074
rect 674833 298016 674838 298072
rect 674894 298016 675298 298072
rect 675354 298016 675359 298072
rect 674833 298014 675359 298016
rect 674833 298011 674899 298014
rect 675293 298011 675359 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 678237 297394 678303 297397
rect 675772 297392 678303 297394
rect 675772 297336 678242 297392
rect 678298 297336 678303 297392
rect 675772 297334 678303 297336
rect 675772 297332 675778 297334
rect 678237 297331 678303 297334
rect 44633 297258 44699 297261
rect 41492 297256 44699 297258
rect 41492 297200 44638 297256
rect 44694 297200 44699 297256
rect 41492 297198 44699 297200
rect 44633 297195 44699 297198
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 674833 296850 674899 296853
rect 676121 296850 676187 296853
rect 674833 296848 676187 296850
rect 674833 296792 674838 296848
rect 674894 296792 676126 296848
rect 676182 296792 676187 296848
rect 674833 296790 676187 296792
rect 674833 296787 674899 296790
rect 676121 296787 676187 296790
rect 675017 296578 675083 296581
rect 675937 296578 676003 296581
rect 675017 296576 676003 296578
rect 675017 296520 675022 296576
rect 675078 296520 675942 296576
rect 675998 296520 676003 296576
rect 675017 296518 676003 296520
rect 675017 296515 675083 296518
rect 675937 296515 676003 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 675753 296304 675819 296309
rect 675753 296248 675758 296304
rect 675814 296248 675819 296304
rect 675753 296243 675819 296248
rect 41321 296034 41387 296037
rect 41308 296032 41387 296034
rect 41308 295976 41326 296032
rect 41382 295976 41387 296032
rect 41308 295974 41387 295976
rect 41321 295971 41387 295974
rect 675756 295901 675816 296243
rect 675753 295896 675819 295901
rect 675753 295840 675758 295896
rect 675814 295840 675819 295896
rect 675753 295835 675819 295840
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 43069 295218 43135 295221
rect 41492 295216 43135 295218
rect 41492 295160 43074 295216
rect 43130 295160 43135 295216
rect 41492 295158 43135 295160
rect 43069 295155 43135 295158
rect 675753 295218 675819 295221
rect 676254 295218 676260 295220
rect 675753 295216 676260 295218
rect 675753 295160 675758 295216
rect 675814 295160 676260 295216
rect 675753 295158 676260 295160
rect 675753 295155 675819 295158
rect 676254 295156 676260 295158
rect 676324 295156 676330 295220
rect 32397 294810 32463 294813
rect 32397 294808 32476 294810
rect 32397 294752 32402 294808
rect 32458 294752 32476 294808
rect 32397 294750 32476 294752
rect 32397 294747 32463 294750
rect 44357 294402 44423 294405
rect 41492 294400 44423 294402
rect 41492 294344 44362 294400
rect 44418 294344 44423 294400
rect 41492 294342 44423 294344
rect 44357 294339 44423 294342
rect 43621 293994 43687 293997
rect 41492 293992 43687 293994
rect 41492 293936 43626 293992
rect 43682 293936 43687 293992
rect 41492 293934 43687 293936
rect 43621 293931 43687 293934
rect 45001 293586 45067 293589
rect 41492 293584 45067 293586
rect 41492 293528 45006 293584
rect 45062 293528 45067 293584
rect 41492 293526 45067 293528
rect 45001 293523 45067 293526
rect 43805 293178 43871 293181
rect 41492 293176 43871 293178
rect 41492 293120 43810 293176
rect 43866 293120 43871 293176
rect 41492 293118 43871 293120
rect 43805 293115 43871 293118
rect 40910 292592 40970 292740
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40542 292332 40602 292528
rect 41781 292500 41847 292501
rect 41781 292496 41828 292500
rect 41892 292498 41898 292500
rect 41781 292440 41786 292496
rect 41781 292436 41828 292440
rect 41892 292438 41938 292498
rect 41892 292436 41898 292438
rect 41781 292435 41847 292436
rect 43989 291954 44055 291957
rect 41492 291952 44055 291954
rect 41492 291896 43994 291952
rect 44050 291896 44055 291952
rect 41492 291894 44055 291896
rect 43989 291891 44055 291894
rect 45185 291682 45251 291685
rect 41830 291680 45251 291682
rect 41830 291624 45190 291680
rect 45246 291624 45251 291680
rect 41830 291622 45251 291624
rect 41830 291546 41890 291622
rect 45185 291619 45251 291622
rect 41492 291486 41890 291546
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 41492 291078 51090 291138
rect 46197 290730 46263 290733
rect 41492 290728 46263 290730
rect 41492 290672 46202 290728
rect 46258 290672 46263 290728
rect 41492 290670 46263 290672
rect 46197 290667 46263 290670
rect 41781 290460 41847 290461
rect 41781 290456 41828 290460
rect 41892 290458 41898 290460
rect 41781 290400 41786 290456
rect 41781 290396 41828 290400
rect 41892 290398 41938 290458
rect 41892 290396 41898 290398
rect 41781 290395 41847 290396
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 49141 289914 49207 289917
rect 41492 289912 49207 289914
rect 41492 289856 49146 289912
rect 49202 289856 49207 289912
rect 41492 289854 49207 289856
rect 51030 289914 51090 291078
rect 673361 290050 673427 290053
rect 675109 290050 675175 290053
rect 673361 290048 675175 290050
rect 673361 289992 673366 290048
rect 673422 289992 675114 290048
rect 675170 289992 675175 290048
rect 673361 289990 675175 289992
rect 673361 289987 673427 289990
rect 675109 289987 675175 289990
rect 51717 289914 51783 289917
rect 51030 289912 51783 289914
rect 51030 289856 51722 289912
rect 51778 289856 51783 289912
rect 51030 289854 51783 289856
rect 49141 289851 49207 289854
rect 51717 289851 51783 289854
rect 672993 287874 673059 287877
rect 675109 287874 675175 287877
rect 672993 287872 675175 287874
rect 672993 287816 672998 287872
rect 673054 287816 675114 287872
rect 675170 287816 675175 287872
rect 672993 287814 675175 287816
rect 672993 287811 673059 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676622 287058 676628 287060
rect 675753 287056 676628 287058
rect 675753 287000 675758 287056
rect 675814 287000 676628 287056
rect 675753 286998 676628 287000
rect 675753 286995 675819 286998
rect 676622 286996 676628 286998
rect 676692 286996 676698 287060
rect 673729 285562 673795 285565
rect 675109 285562 675175 285565
rect 673729 285560 675175 285562
rect 673729 285504 673734 285560
rect 673790 285504 675114 285560
rect 675170 285504 675175 285560
rect 673729 285502 675175 285504
rect 673729 285499 673795 285502
rect 675109 285499 675175 285502
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62941 285154 63007 285157
rect 62941 285152 64492 285154
rect 62941 285096 62946 285152
rect 63002 285096 64492 285152
rect 62941 285094 64492 285096
rect 62941 285091 63007 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 42149 279850 42215 279853
rect 43805 279850 43871 279853
rect 42149 279848 43871 279850
rect 42149 279792 42154 279848
rect 42210 279792 43810 279848
rect 43866 279792 43871 279848
rect 42149 279790 43871 279792
rect 42149 279787 42215 279790
rect 43805 279787 43871 279790
rect 42425 278762 42491 278765
rect 55857 278762 55923 278765
rect 42425 278760 55923 278762
rect 42425 278704 42430 278760
rect 42486 278704 55862 278760
rect 55918 278704 55923 278760
rect 42425 278702 55923 278704
rect 42425 278699 42491 278702
rect 55857 278699 55923 278702
rect 40718 278428 40724 278492
rect 40788 278490 40794 278492
rect 42333 278490 42399 278493
rect 40788 278488 42399 278490
rect 40788 278432 42338 278488
rect 42394 278432 42399 278488
rect 40788 278430 42399 278432
rect 40788 278428 40794 278430
rect 42333 278427 42399 278430
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 41781 277946 41847 277949
rect 40972 277944 41847 277946
rect 40972 277888 41786 277944
rect 41842 277888 41847 277944
rect 40972 277886 41847 277888
rect 40972 277884 40978 277886
rect 41781 277883 41847 277886
rect 42149 277946 42215 277949
rect 45185 277946 45251 277949
rect 42149 277944 45251 277946
rect 42149 277888 42154 277944
rect 42210 277888 45190 277944
rect 45246 277888 45251 277944
rect 42149 277886 45251 277888
rect 42149 277883 42215 277886
rect 45185 277883 45251 277886
rect 42057 277130 42123 277133
rect 43989 277130 44055 277133
rect 42057 277128 44055 277130
rect 42057 277072 42062 277128
rect 42118 277072 43994 277128
rect 44050 277072 44055 277128
rect 42057 277070 44055 277072
rect 42057 277067 42123 277070
rect 43989 277067 44055 277070
rect 42057 276586 42123 276589
rect 43069 276586 43135 276589
rect 42057 276584 43135 276586
rect 42057 276528 42062 276584
rect 42118 276528 43074 276584
rect 43130 276528 43135 276584
rect 42057 276526 43135 276528
rect 42057 276523 42123 276526
rect 43069 276523 43135 276526
rect 525793 275770 525859 275773
rect 527357 275770 527423 275773
rect 525793 275768 527423 275770
rect 525793 275712 525798 275768
rect 525854 275712 527362 275768
rect 527418 275712 527423 275768
rect 525793 275710 527423 275712
rect 525793 275707 525859 275710
rect 527357 275707 527423 275710
rect 534901 275770 534967 275773
rect 538029 275770 538095 275773
rect 534901 275768 538095 275770
rect 534901 275712 534906 275768
rect 534962 275712 538034 275768
rect 538090 275712 538095 275768
rect 534901 275710 538095 275712
rect 534901 275707 534967 275710
rect 538029 275707 538095 275710
rect 538213 275498 538279 275501
rect 539041 275498 539107 275501
rect 538213 275496 539107 275498
rect 538213 275440 538218 275496
rect 538274 275440 539046 275496
rect 539102 275440 539107 275496
rect 538213 275438 539107 275440
rect 538213 275435 538279 275438
rect 539041 275435 539107 275438
rect 535085 275090 535151 275093
rect 538397 275090 538463 275093
rect 535085 275088 538463 275090
rect 535085 275032 535090 275088
rect 535146 275032 538402 275088
rect 538458 275032 538463 275088
rect 535085 275030 538463 275032
rect 535085 275027 535151 275030
rect 538397 275027 538463 275030
rect 538673 275090 538739 275093
rect 541157 275090 541223 275093
rect 538673 275088 541223 275090
rect 538673 275032 538678 275088
rect 538734 275032 541162 275088
rect 541218 275032 541223 275088
rect 538673 275030 541223 275032
rect 538673 275027 538739 275030
rect 541157 275027 541223 275030
rect 538213 274818 538279 274821
rect 543181 274818 543247 274821
rect 538213 274816 543247 274818
rect 538213 274760 538218 274816
rect 538274 274760 543186 274816
rect 543242 274760 543247 274816
rect 538213 274758 543247 274760
rect 538213 274755 538279 274758
rect 543181 274755 543247 274758
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 533889 274274 533955 274277
rect 539041 274274 539107 274277
rect 533889 274272 539107 274274
rect 533889 274216 533894 274272
rect 533950 274216 539046 274272
rect 539102 274216 539107 274272
rect 533889 274214 539107 274216
rect 533889 274211 533955 274214
rect 539041 274211 539107 274214
rect 516593 274138 516659 274141
rect 517053 274138 517119 274141
rect 516593 274136 517119 274138
rect 516593 274080 516598 274136
rect 516654 274080 517058 274136
rect 517114 274080 517119 274136
rect 516593 274078 517119 274080
rect 516593 274075 516659 274078
rect 517053 274075 517119 274078
rect 528001 273866 528067 273869
rect 533889 273866 533955 273869
rect 528001 273864 533955 273866
rect 528001 273808 528006 273864
rect 528062 273808 533894 273864
rect 533950 273808 533955 273864
rect 528001 273806 533955 273808
rect 528001 273803 528067 273806
rect 533889 273803 533955 273806
rect 536741 273866 536807 273869
rect 635641 273866 635707 273869
rect 536741 273864 635707 273866
rect 536741 273808 536746 273864
rect 536802 273808 635646 273864
rect 635702 273808 635707 273864
rect 536741 273806 635707 273808
rect 536741 273803 536807 273806
rect 635641 273803 635707 273806
rect 521101 273730 521167 273733
rect 524229 273730 524295 273733
rect 521101 273728 524295 273730
rect 521101 273672 521106 273728
rect 521162 273672 524234 273728
rect 524290 273672 524295 273728
rect 521101 273670 524295 273672
rect 521101 273667 521167 273670
rect 524229 273667 524295 273670
rect 42057 273458 42123 273461
rect 45001 273458 45067 273461
rect 42057 273456 45067 273458
rect 42057 273400 42062 273456
rect 42118 273400 45006 273456
rect 45062 273400 45067 273456
rect 42057 273398 45067 273400
rect 42057 273395 42123 273398
rect 45001 273395 45067 273398
rect 42057 273050 42123 273053
rect 43621 273050 43687 273053
rect 42057 273048 43687 273050
rect 42057 272992 42062 273048
rect 42118 272992 43626 273048
rect 43682 272992 43687 273048
rect 42057 272990 43687 272992
rect 42057 272987 42123 272990
rect 43621 272987 43687 272990
rect 534073 272778 534139 272781
rect 544469 272778 544535 272781
rect 534073 272776 544535 272778
rect 534073 272720 534078 272776
rect 534134 272720 544474 272776
rect 544530 272720 544535 272776
rect 534073 272718 544535 272720
rect 534073 272715 534139 272718
rect 544469 272715 544535 272718
rect 521469 272642 521535 272645
rect 524873 272642 524939 272645
rect 521469 272640 524939 272642
rect 521469 272584 521474 272640
rect 521530 272584 524878 272640
rect 524934 272584 524939 272640
rect 521469 272582 524939 272584
rect 521469 272579 521535 272582
rect 524873 272579 524939 272582
rect 533705 272506 533771 272509
rect 534165 272506 534231 272509
rect 533705 272504 534231 272506
rect 533705 272448 533710 272504
rect 533766 272448 534170 272504
rect 534226 272448 534231 272504
rect 533705 272446 534231 272448
rect 533705 272443 533771 272446
rect 534165 272443 534231 272446
rect 542997 272506 543063 272509
rect 645117 272506 645183 272509
rect 542997 272504 645183 272506
rect 542997 272448 543002 272504
rect 543058 272448 645122 272504
rect 645178 272448 645183 272504
rect 542997 272446 645183 272448
rect 542997 272443 543063 272446
rect 645117 272443 645183 272446
rect 513189 272370 513255 272373
rect 518433 272370 518499 272373
rect 513189 272368 518499 272370
rect 513189 272312 513194 272368
rect 513250 272312 518438 272368
rect 518494 272312 518499 272368
rect 513189 272310 518499 272312
rect 513189 272307 513255 272310
rect 518433 272307 518499 272310
rect 524505 272370 524571 272373
rect 531589 272370 531655 272373
rect 524505 272368 531655 272370
rect 524505 272312 524510 272368
rect 524566 272312 531594 272368
rect 531650 272312 531655 272368
rect 524505 272310 531655 272312
rect 524505 272307 524571 272310
rect 531589 272307 531655 272310
rect 523953 271690 524019 271693
rect 524689 271690 524755 271693
rect 523953 271688 524755 271690
rect 523953 271632 523958 271688
rect 524014 271632 524694 271688
rect 524750 271632 524755 271688
rect 523953 271630 524755 271632
rect 523953 271627 524019 271630
rect 524689 271627 524755 271630
rect 543549 271554 543615 271557
rect 546217 271554 546283 271557
rect 543549 271552 546283 271554
rect 543549 271496 543554 271552
rect 543610 271496 546222 271552
rect 546278 271496 546283 271552
rect 543549 271494 546283 271496
rect 543549 271491 543615 271494
rect 546217 271491 546283 271494
rect 511717 271418 511783 271421
rect 515305 271418 515371 271421
rect 511717 271416 515371 271418
rect 511717 271360 511722 271416
rect 511778 271360 515310 271416
rect 515366 271360 515371 271416
rect 511717 271358 515371 271360
rect 511717 271355 511783 271358
rect 515305 271355 515371 271358
rect 529197 271282 529263 271285
rect 529197 271280 534090 271282
rect 529197 271224 529202 271280
rect 529258 271224 534090 271280
rect 529197 271222 534090 271224
rect 529197 271219 529263 271222
rect 534030 271146 534090 271222
rect 625061 271146 625127 271149
rect 534030 271144 625127 271146
rect 534030 271088 625066 271144
rect 625122 271088 625127 271144
rect 534030 271086 625127 271088
rect 625061 271083 625127 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 526253 271010 526319 271013
rect 529565 271010 529631 271013
rect 526253 271008 529631 271010
rect 526253 270952 526258 271008
rect 526314 270952 529570 271008
rect 529626 270952 529631 271008
rect 526253 270950 529631 270952
rect 526253 270947 526319 270950
rect 529565 270947 529631 270950
rect 522021 270874 522087 270877
rect 524781 270874 524847 270877
rect 522021 270872 524847 270874
rect 522021 270816 522026 270872
rect 522082 270816 524786 270872
rect 524842 270816 524847 270872
rect 522021 270814 524847 270816
rect 522021 270811 522087 270814
rect 524781 270811 524847 270814
rect 528645 270738 528711 270741
rect 533153 270738 533219 270741
rect 528645 270736 533219 270738
rect 528645 270680 528650 270736
rect 528706 270680 533158 270736
rect 533214 270680 533219 270736
rect 528645 270678 533219 270680
rect 528645 270675 528711 270678
rect 533153 270675 533219 270678
rect 552197 270738 552263 270741
rect 553393 270738 553459 270741
rect 552197 270736 553459 270738
rect 552197 270680 552202 270736
rect 552258 270680 553398 270736
rect 553454 270680 553459 270736
rect 552197 270678 553459 270680
rect 552197 270675 552263 270678
rect 553393 270675 553459 270678
rect 504173 270602 504239 270605
rect 507853 270602 507919 270605
rect 504173 270600 507919 270602
rect 504173 270544 504178 270600
rect 504234 270544 507858 270600
rect 507914 270544 507919 270600
rect 504173 270542 507919 270544
rect 504173 270539 504239 270542
rect 507853 270539 507919 270542
rect 538305 270602 538371 270605
rect 543549 270602 543615 270605
rect 538305 270600 543615 270602
rect 538305 270544 538310 270600
rect 538366 270544 543554 270600
rect 543610 270544 543615 270600
rect 538305 270542 543615 270544
rect 538305 270539 538371 270542
rect 543549 270539 543615 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 42425 270466 42491 270469
rect 44357 270466 44423 270469
rect 42425 270464 44423 270466
rect 42425 270408 42430 270464
rect 42486 270408 44362 270464
rect 44418 270408 44423 270464
rect 42425 270406 44423 270408
rect 42425 270403 42491 270406
rect 44357 270403 44423 270406
rect 574921 270330 574987 270333
rect 499530 270328 574987 270330
rect 499530 270272 574926 270328
rect 574982 270272 574987 270328
rect 499530 270270 574987 270272
rect 494145 270058 494211 270061
rect 499530 270058 499590 270270
rect 574921 270267 574987 270270
rect 494145 270056 499590 270058
rect 494145 270000 494150 270056
rect 494206 270000 499590 270056
rect 494145 269998 499590 270000
rect 531405 270058 531471 270061
rect 627913 270058 627979 270061
rect 531405 270056 627979 270058
rect 531405 270000 531410 270056
rect 531466 270000 627918 270056
rect 627974 270000 627979 270056
rect 531405 269998 627979 270000
rect 494145 269995 494211 269998
rect 531405 269995 531471 269998
rect 627913 269995 627979 269998
rect 136541 269786 136607 269789
rect 139945 269786 140011 269789
rect 136541 269784 140011 269786
rect 136541 269728 136546 269784
rect 136602 269728 139950 269784
rect 140006 269728 140011 269784
rect 136541 269726 140011 269728
rect 136541 269723 136607 269726
rect 139945 269723 140011 269726
rect 509877 269786 509943 269789
rect 523309 269786 523375 269789
rect 509877 269784 523375 269786
rect 509877 269728 509882 269784
rect 509938 269728 523314 269784
rect 523370 269728 523375 269784
rect 509877 269726 523375 269728
rect 509877 269723 509943 269726
rect 523309 269723 523375 269726
rect 533521 269786 533587 269789
rect 534349 269786 534415 269789
rect 533521 269784 534415 269786
rect 533521 269728 533526 269784
rect 533582 269728 534354 269784
rect 534410 269728 534415 269784
rect 533521 269726 534415 269728
rect 533521 269723 533587 269726
rect 534349 269723 534415 269726
rect 538029 269786 538095 269789
rect 637573 269786 637639 269789
rect 538029 269784 637639 269786
rect 538029 269728 538034 269784
rect 538090 269728 637578 269784
rect 637634 269728 637639 269784
rect 538029 269726 637639 269728
rect 538029 269723 538095 269726
rect 637573 269723 637639 269726
rect 671337 269786 671403 269789
rect 676029 269786 676095 269789
rect 671337 269784 676095 269786
rect 671337 269728 671342 269784
rect 671398 269728 676034 269784
rect 676090 269728 676095 269784
rect 671337 269726 676095 269728
rect 671337 269723 671403 269726
rect 676029 269723 676095 269726
rect 503069 269650 503135 269653
rect 504541 269650 504607 269653
rect 503069 269648 504607 269650
rect 503069 269592 503074 269648
rect 503130 269592 504546 269648
rect 504602 269592 504607 269648
rect 503069 269590 504607 269592
rect 503069 269587 503135 269590
rect 504541 269587 504607 269590
rect 521653 269514 521719 269517
rect 530945 269514 531011 269517
rect 521653 269512 531011 269514
rect 521653 269456 521658 269512
rect 521714 269456 530950 269512
rect 531006 269456 531011 269512
rect 521653 269454 531011 269456
rect 521653 269451 521719 269454
rect 530945 269451 531011 269454
rect 535913 269514 535979 269517
rect 541985 269514 542051 269517
rect 535913 269512 542051 269514
rect 535913 269456 535918 269512
rect 535974 269456 541990 269512
rect 542046 269456 542051 269512
rect 535913 269454 542051 269456
rect 535913 269451 535979 269454
rect 541985 269451 542051 269454
rect 537017 269242 537083 269245
rect 538673 269242 538739 269245
rect 537017 269240 538739 269242
rect 537017 269184 537022 269240
rect 537078 269184 538678 269240
rect 538734 269184 538739 269240
rect 537017 269182 538739 269184
rect 537017 269179 537083 269182
rect 538673 269179 538739 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 530945 269106 531011 269109
rect 533889 269106 533955 269109
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 530945 269104 533955 269106
rect 530945 269048 530950 269104
rect 531006 269048 533894 269104
rect 533950 269048 533955 269104
rect 530945 269046 533955 269048
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 530945 269043 531011 269046
rect 533889 269043 533955 269046
rect 525517 268698 525583 268701
rect 533889 268698 533955 268701
rect 525517 268696 533955 268698
rect 525517 268640 525522 268696
rect 525578 268640 533894 268696
rect 533950 268640 533955 268696
rect 525517 268638 533955 268640
rect 525517 268635 525583 268638
rect 533889 268635 533955 268638
rect 518433 268562 518499 268565
rect 518985 268562 519051 268565
rect 676262 268562 676322 268668
rect 518433 268560 519051 268562
rect 518433 268504 518438 268560
rect 518494 268504 518990 268560
rect 519046 268504 519051 268560
rect 518433 268502 519051 268504
rect 518433 268499 518499 268502
rect 518985 268499 519051 268502
rect 663750 268502 676322 268562
rect 519169 268426 519235 268429
rect 520457 268426 520523 268429
rect 519169 268424 520523 268426
rect 519169 268368 519174 268424
rect 519230 268368 520462 268424
rect 520518 268368 520523 268424
rect 519169 268366 520523 268368
rect 519169 268363 519235 268366
rect 520457 268363 520523 268366
rect 547505 268426 547571 268429
rect 549253 268426 549319 268429
rect 547505 268424 549319 268426
rect 547505 268368 547510 268424
rect 547566 268368 549258 268424
rect 549314 268368 549319 268424
rect 547505 268366 549319 268368
rect 547505 268363 547571 268366
rect 549253 268363 549319 268366
rect 539225 268154 539291 268157
rect 547689 268154 547755 268157
rect 539225 268152 547755 268154
rect 539225 268096 539230 268152
rect 539286 268096 547694 268152
rect 547750 268096 547755 268152
rect 539225 268094 547755 268096
rect 539225 268091 539291 268094
rect 547689 268091 547755 268094
rect 661677 268154 661743 268157
rect 663750 268154 663810 268502
rect 676029 268290 676095 268293
rect 676029 268288 676292 268290
rect 676029 268232 676034 268288
rect 676090 268232 676292 268288
rect 676029 268230 676292 268232
rect 676029 268227 676095 268230
rect 683113 268154 683179 268157
rect 661677 268152 663810 268154
rect 661677 268096 661682 268152
rect 661738 268096 663810 268152
rect 661677 268094 663810 268096
rect 682886 268152 683179 268154
rect 682886 268096 683118 268152
rect 683174 268096 683179 268152
rect 682886 268094 683179 268096
rect 661677 268091 661743 268094
rect 533889 268018 533955 268021
rect 535453 268018 535519 268021
rect 533889 268016 535519 268018
rect 533889 267960 533894 268016
rect 533950 267960 535458 268016
rect 535514 267960 535519 268016
rect 533889 267958 535519 267960
rect 533889 267955 533955 267958
rect 535453 267955 535519 267958
rect 492305 267882 492371 267885
rect 498193 267882 498259 267885
rect 492305 267880 498259 267882
rect 492305 267824 492310 267880
rect 492366 267824 498198 267880
rect 498254 267824 498259 267880
rect 682886 267852 682946 268094
rect 683113 268091 683179 268094
rect 492305 267822 498259 267824
rect 492305 267819 492371 267822
rect 498193 267819 498259 267822
rect 516961 267746 517027 267749
rect 518985 267746 519051 267749
rect 516961 267744 519051 267746
rect 516961 267688 516966 267744
rect 517022 267688 518990 267744
rect 519046 267688 519051 267744
rect 516961 267686 519051 267688
rect 516961 267683 517027 267686
rect 518985 267683 519051 267686
rect 533981 267746 534047 267749
rect 538305 267746 538371 267749
rect 533981 267744 538371 267746
rect 533981 267688 533986 267744
rect 534042 267688 538310 267744
rect 538366 267688 538371 267744
rect 533981 267686 538371 267688
rect 533981 267683 534047 267686
rect 538305 267683 538371 267686
rect 543549 267746 543615 267749
rect 546585 267746 546651 267749
rect 543549 267744 546651 267746
rect 543549 267688 543554 267744
rect 543610 267688 546590 267744
rect 546646 267688 546651 267744
rect 543549 267686 546651 267688
rect 543549 267683 543615 267686
rect 546585 267683 546651 267686
rect 485727 267474 485793 267477
rect 487245 267474 487311 267477
rect 485727 267472 487311 267474
rect 485727 267416 485732 267472
rect 485788 267416 487250 267472
rect 487306 267416 487311 267472
rect 485727 267414 487311 267416
rect 485727 267411 485793 267414
rect 487245 267411 487311 267414
rect 673913 267474 673979 267477
rect 673913 267472 676292 267474
rect 673913 267416 673918 267472
rect 673974 267416 676292 267472
rect 673913 267414 676292 267416
rect 673913 267411 673979 267414
rect 533889 267338 533955 267341
rect 534165 267338 534231 267341
rect 533889 267336 534231 267338
rect 533889 267280 533894 267336
rect 533950 267280 534170 267336
rect 534226 267280 534231 267336
rect 533889 267278 534231 267280
rect 533889 267275 533955 267278
rect 534165 267275 534231 267278
rect 542169 267338 542235 267341
rect 607857 267338 607923 267341
rect 542169 267336 607923 267338
rect 542169 267280 542174 267336
rect 542230 267280 607862 267336
rect 607918 267280 607923 267336
rect 542169 267278 607923 267280
rect 542169 267275 542235 267278
rect 607857 267275 607923 267278
rect 499573 267202 499639 267205
rect 501045 267202 501111 267205
rect 499573 267200 501111 267202
rect 499573 267144 499578 267200
rect 499634 267144 501050 267200
rect 501106 267144 501111 267200
rect 499573 267142 501111 267144
rect 499573 267139 499639 267142
rect 501045 267139 501111 267142
rect 519169 267202 519235 267205
rect 527173 267202 527239 267205
rect 519169 267200 527239 267202
rect 519169 267144 519174 267200
rect 519230 267144 527178 267200
rect 527234 267144 527239 267200
rect 519169 267142 527239 267144
rect 519169 267139 519235 267142
rect 527173 267139 527239 267142
rect 40677 267066 40743 267069
rect 62757 267066 62823 267069
rect 40677 267064 62823 267066
rect 40677 267008 40682 267064
rect 40738 267008 62762 267064
rect 62818 267008 62823 267064
rect 40677 267006 62823 267008
rect 40677 267003 40743 267006
rect 62757 267003 62823 267006
rect 532233 267066 532299 267069
rect 629293 267066 629359 267069
rect 532233 267064 629359 267066
rect 532233 267008 532238 267064
rect 532294 267008 629298 267064
rect 629354 267008 629359 267064
rect 532233 267006 629359 267008
rect 532233 267003 532299 267006
rect 629293 267003 629359 267006
rect 674649 267066 674715 267069
rect 674649 267064 676292 267066
rect 674649 267008 674654 267064
rect 674710 267008 676292 267064
rect 674649 267006 676292 267008
rect 674649 267003 674715 267006
rect 485681 266930 485747 266933
rect 486049 266930 486115 266933
rect 485681 266928 486115 266930
rect 485681 266872 485686 266928
rect 485742 266872 486054 266928
rect 486110 266872 486115 266928
rect 485681 266870 486115 266872
rect 485681 266867 485747 266870
rect 486049 266867 486115 266870
rect 538673 266658 538739 266661
rect 543549 266658 543615 266661
rect 538673 266656 543615 266658
rect 538673 266600 538678 266656
rect 538734 266600 543554 266656
rect 543610 266600 543615 266656
rect 538673 266598 543615 266600
rect 538673 266595 538739 266598
rect 543549 266595 543615 266598
rect 673177 266522 673243 266525
rect 676262 266522 676322 266628
rect 673177 266520 676322 266522
rect 673177 266464 673182 266520
rect 673238 266464 676322 266520
rect 673177 266462 676322 266464
rect 673177 266459 673243 266462
rect 674005 266250 674071 266253
rect 674005 266248 676292 266250
rect 674005 266192 674010 266248
rect 674066 266192 676292 266248
rect 674005 266190 676292 266192
rect 674005 266187 674071 266190
rect 674465 265842 674531 265845
rect 674465 265840 676292 265842
rect 674465 265784 674470 265840
rect 674526 265784 676292 265840
rect 674465 265782 676292 265784
rect 674465 265779 674531 265782
rect 674373 265434 674439 265437
rect 674373 265432 676292 265434
rect 674373 265376 674378 265432
rect 674434 265376 676292 265432
rect 674373 265374 676292 265376
rect 674373 265371 674439 265374
rect 674189 265026 674255 265029
rect 674189 265024 676292 265026
rect 674189 264968 674194 265024
rect 674250 264968 676292 265024
rect 674189 264966 676292 264968
rect 674189 264963 674255 264966
rect 674833 264482 674899 264485
rect 676262 264482 676322 264588
rect 674833 264480 676322 264482
rect 674833 264424 674838 264480
rect 674894 264424 676322 264480
rect 674833 264422 676322 264424
rect 674833 264419 674899 264422
rect 676446 264077 676506 264180
rect 671521 264074 671587 264077
rect 671521 264072 676322 264074
rect 671521 264016 671526 264072
rect 671582 264016 676322 264072
rect 671521 264014 676322 264016
rect 676446 264072 676555 264077
rect 676446 264016 676494 264072
rect 676550 264016 676555 264072
rect 676446 264014 676555 264016
rect 671521 264011 671587 264014
rect 673177 263802 673243 263805
rect 674833 263802 674899 263805
rect 673177 263800 674899 263802
rect 673177 263744 673182 263800
rect 673238 263744 674838 263800
rect 674894 263744 674899 263800
rect 676262 263772 676322 264014
rect 676489 264011 676555 264014
rect 673177 263742 674899 263744
rect 673177 263739 673243 263742
rect 674833 263739 674899 263742
rect 674966 263604 674972 263668
rect 675036 263666 675042 263668
rect 676489 263666 676555 263669
rect 675036 263664 676555 263666
rect 675036 263608 676494 263664
rect 676550 263608 676555 263664
rect 675036 263606 676555 263608
rect 675036 263604 675042 263606
rect 676489 263603 676555 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 676070 262380 676076 262444
rect 676140 262442 676146 262444
rect 676262 262442 676322 262548
rect 676140 262382 676322 262442
rect 676140 262380 676146 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671337 262170 671403 262173
rect 671337 262168 676292 262170
rect 671337 262112 671342 262168
rect 671398 262112 676292 262168
rect 671337 262110 676292 262112
rect 671337 262107 671403 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 678470 261221 678530 261324
rect 678421 261216 678530 261221
rect 678421 261160 678426 261216
rect 678482 261160 678530 261216
rect 678421 261158 678530 261160
rect 678421 261155 678487 261158
rect 674281 260946 674347 260949
rect 674281 260944 676292 260946
rect 674281 260888 674286 260944
rect 674342 260888 676292 260944
rect 674281 260886 676292 260888
rect 674281 260883 674347 260886
rect 676262 260402 676322 260508
rect 672996 260342 676322 260402
rect 672996 260133 673056 260342
rect 672993 260128 673059 260133
rect 672993 260072 672998 260128
rect 673054 260072 673059 260128
rect 672993 260067 673059 260072
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 673729 259722 673795 259725
rect 673729 259720 676292 259722
rect 673729 259664 673734 259720
rect 673790 259664 676292 259720
rect 673729 259662 676292 259664
rect 673729 259659 673795 259662
rect 673361 259314 673427 259317
rect 673361 259312 676292 259314
rect 673361 259256 673366 259312
rect 673422 259256 676292 259312
rect 673361 259254 676292 259256
rect 673361 259251 673427 259254
rect 671797 258906 671863 258909
rect 671797 258904 676292 258906
rect 671797 258848 671802 258904
rect 671858 258848 676292 258904
rect 671797 258846 676292 258848
rect 671797 258843 671863 258846
rect 673913 258498 673979 258501
rect 673913 258496 676292 258498
rect 673913 258440 673918 258496
rect 673974 258440 676292 258496
rect 673913 258438 676292 258440
rect 673913 258435 673979 258438
rect 41492 258030 42074 258090
rect 42014 257954 42074 258030
rect 42014 257894 45570 257954
rect 45510 257818 45570 257894
rect 50337 257818 50403 257821
rect 553945 257818 554011 257821
rect 45510 257816 50403 257818
rect 45510 257760 50342 257816
rect 50398 257760 50403 257816
rect 45510 257758 50403 257760
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 50337 257755 50403 257758
rect 553945 257755 554011 257758
rect 43437 257682 43503 257685
rect 41492 257680 43503 257682
rect 41492 257624 43442 257680
rect 43498 257624 43503 257680
rect 41492 257622 43503 257624
rect 43437 257619 43503 257622
rect 670417 257682 670483 257685
rect 676262 257682 676322 258060
rect 670417 257680 676322 257682
rect 670417 257624 670422 257680
rect 670478 257652 676322 257680
rect 670478 257624 676292 257652
rect 670417 257622 676292 257624
rect 670417 257619 670483 257622
rect 35758 257141 35818 257244
rect 672582 257214 676292 257274
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 672582 257005 672642 257214
rect 672582 257000 672691 257005
rect 672582 256944 672630 257000
rect 672686 256944 672691 257000
rect 672582 256942 672691 256944
rect 672625 256939 672691 256942
rect 42885 256866 42951 256869
rect 41492 256864 42951 256866
rect 41492 256808 42890 256864
rect 42946 256808 42951 256864
rect 41492 256806 42951 256808
rect 42885 256803 42951 256806
rect 43621 256458 43687 256461
rect 41492 256456 43687 256458
rect 41492 256400 43626 256456
rect 43682 256400 43687 256456
rect 41492 256398 43687 256400
rect 43621 256395 43687 256398
rect 43253 256050 43319 256053
rect 41492 256048 43319 256050
rect 41492 255992 43258 256048
rect 43314 255992 43319 256048
rect 41492 255990 43319 255992
rect 43253 255987 43319 255990
rect 42977 255642 43043 255645
rect 553669 255642 553735 255645
rect 41492 255640 43043 255642
rect 41492 255584 42982 255640
rect 43038 255584 43043 255640
rect 41492 255582 43043 255584
rect 552460 255640 553735 255642
rect 552460 255584 553674 255640
rect 553730 255584 553735 255640
rect 552460 255582 553735 255584
rect 42977 255579 43043 255582
rect 553669 255579 553735 255582
rect 44173 255234 44239 255237
rect 41492 255232 44239 255234
rect 41492 255176 44178 255232
rect 44234 255176 44239 255232
rect 41492 255174 44239 255176
rect 44173 255171 44239 255174
rect 42793 254826 42859 254829
rect 41492 254824 42859 254826
rect 41492 254768 42798 254824
rect 42854 254768 42859 254824
rect 41492 254766 42859 254768
rect 42793 254763 42859 254766
rect 44633 254418 44699 254421
rect 41492 254416 44699 254418
rect 41492 254360 44638 254416
rect 44694 254360 44699 254416
rect 41492 254358 44699 254360
rect 44633 254355 44699 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35390 253469 35450 253572
rect 35390 253464 35499 253469
rect 554497 253466 554563 253469
rect 35390 253408 35438 253464
rect 35494 253408 35499 253464
rect 35390 253406 35499 253408
rect 552460 253464 554563 253466
rect 552460 253408 554502 253464
rect 554558 253408 554563 253464
rect 552460 253406 554563 253408
rect 35433 253403 35499 253406
rect 554497 253403 554563 253406
rect 35574 253061 35634 253164
rect 35574 253056 35683 253061
rect 35574 253000 35622 253056
rect 35678 253000 35683 253056
rect 35574 252998 35683 253000
rect 35617 252995 35683 252998
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 41321 252242 41387 252245
rect 42609 252242 42675 252245
rect 41321 252240 42675 252242
rect 41321 252184 41326 252240
rect 41382 252184 42614 252240
rect 42670 252184 42675 252240
rect 41321 252182 42675 252184
rect 41321 252179 41387 252182
rect 42609 252179 42675 252182
rect 44541 251970 44607 251973
rect 41492 251968 44607 251970
rect 41492 251912 44546 251968
rect 44602 251912 44607 251968
rect 41492 251910 44607 251912
rect 44541 251907 44607 251910
rect 674925 251562 674991 251565
rect 675845 251562 675911 251565
rect 674925 251560 675911 251562
rect 40726 251428 40786 251532
rect 674925 251504 674930 251560
rect 674986 251504 675850 251560
rect 675906 251504 675911 251560
rect 674925 251502 675911 251504
rect 674925 251499 674991 251502
rect 675845 251499 675911 251502
rect 40718 251364 40724 251428
rect 40788 251364 40794 251428
rect 553485 251290 553551 251293
rect 552460 251288 553551 251290
rect 552460 251232 553490 251288
rect 553546 251232 553551 251288
rect 552460 251230 553551 251232
rect 553485 251227 553551 251230
rect 43437 251154 43503 251157
rect 41492 251152 43503 251154
rect 41492 251096 43442 251152
rect 43498 251096 43503 251152
rect 41492 251094 43503 251096
rect 43437 251091 43503 251094
rect 45553 250746 45619 250749
rect 41492 250744 45619 250746
rect 41492 250688 45558 250744
rect 45614 250688 45619 250744
rect 41492 250686 45619 250688
rect 45553 250683 45619 250686
rect 45829 250338 45895 250341
rect 41492 250336 45895 250338
rect 41492 250280 45834 250336
rect 45890 250280 45895 250336
rect 41492 250278 45895 250280
rect 45829 250275 45895 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675385 249658 675451 249661
rect 674852 249656 675451 249658
rect 674852 249600 675390 249656
rect 675446 249600 675451 249656
rect 674852 249598 675451 249600
rect 674852 249596 674858 249598
rect 675385 249595 675451 249598
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 674925 249386 674991 249389
rect 676078 249386 676138 249596
rect 674925 249384 676138 249386
rect 674925 249328 674930 249384
rect 674986 249328 676138 249384
rect 674925 249326 676138 249328
rect 674925 249323 674991 249326
rect 43713 249114 43779 249117
rect 553853 249114 553919 249117
rect 41492 249112 43779 249114
rect 41492 249056 43718 249112
rect 43774 249056 43779 249112
rect 41492 249054 43779 249056
rect 552460 249112 553919 249114
rect 552460 249056 553858 249112
rect 553914 249056 553919 249112
rect 552460 249054 553919 249056
rect 43713 249051 43779 249054
rect 553853 249051 553919 249054
rect 44357 248706 44423 248709
rect 41492 248704 44423 248706
rect 41492 248648 44362 248704
rect 44418 248648 44423 248704
rect 41492 248646 44423 248648
rect 44357 248643 44423 248646
rect 45001 248298 45067 248301
rect 41492 248296 45067 248298
rect 41492 248240 45006 248296
rect 45062 248240 45067 248296
rect 41492 248238 45067 248240
rect 45001 248235 45067 248238
rect 41462 247754 41522 247860
rect 50521 247754 50587 247757
rect 41462 247752 50587 247754
rect 41462 247696 50526 247752
rect 50582 247696 50587 247752
rect 41462 247694 50587 247696
rect 50521 247691 50587 247694
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46933 247074 46999 247077
rect 41492 247072 46999 247074
rect 41492 247016 46938 247072
rect 46994 247016 46999 247072
rect 41492 247014 46999 247016
rect 46933 247011 46999 247014
rect 554405 246938 554471 246941
rect 552460 246936 554471 246938
rect 552460 246880 554410 246936
rect 554466 246880 554471 246936
rect 552460 246878 554471 246880
rect 554405 246875 554471 246878
rect 674281 246938 674347 246941
rect 675109 246938 675175 246941
rect 674281 246936 675175 246938
rect 674281 246880 674286 246936
rect 674342 246880 675114 246936
rect 675170 246880 675175 246936
rect 674281 246878 675175 246880
rect 674281 246875 674347 246878
rect 675109 246875 675175 246878
rect 41462 246530 41522 246636
rect 50337 246530 50403 246533
rect 41462 246528 50403 246530
rect 41462 246472 50342 246528
rect 50398 246472 50403 246528
rect 41462 246470 50403 246472
rect 50337 246467 50403 246470
rect 673729 245578 673795 245581
rect 675109 245578 675175 245581
rect 673729 245576 675175 245578
rect 673729 245520 673734 245576
rect 673790 245520 675114 245576
rect 675170 245520 675175 245576
rect 673729 245518 675175 245520
rect 673729 245515 673795 245518
rect 675109 245515 675175 245518
rect 674833 245306 674899 245309
rect 676806 245306 676812 245308
rect 674833 245304 676812 245306
rect 674833 245248 674838 245304
rect 674894 245248 676812 245304
rect 674833 245246 676812 245248
rect 674833 245243 674899 245246
rect 676806 245244 676812 245246
rect 676876 245244 676882 245308
rect 672993 245034 673059 245037
rect 675150 245034 675156 245036
rect 672993 245032 675156 245034
rect 672993 244976 672998 245032
rect 673054 244976 675156 245032
rect 672993 244974 675156 244976
rect 672993 244971 673059 244974
rect 675150 244972 675156 244974
rect 675220 244972 675226 245036
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 671337 244762 671403 244765
rect 675334 244762 675340 244764
rect 671337 244760 675340 244762
rect 671337 244704 671342 244760
rect 671398 244704 675340 244760
rect 671337 244702 675340 244704
rect 671337 244699 671403 244702
rect 675334 244700 675340 244702
rect 675404 244700 675410 244764
rect 41689 242858 41755 242861
rect 42333 242858 42399 242861
rect 41689 242856 42399 242858
rect 41689 242800 41694 242856
rect 41750 242800 42338 242856
rect 42394 242800 42399 242856
rect 41689 242798 42399 242800
rect 41689 242795 41755 242798
rect 42333 242795 42399 242798
rect 673361 242858 673427 242861
rect 675109 242858 675175 242861
rect 673361 242856 675175 242858
rect 673361 242800 673366 242856
rect 673422 242800 675114 242856
rect 675170 242800 675175 242856
rect 673361 242798 675175 242800
rect 673361 242795 673427 242798
rect 675109 242795 675175 242798
rect 40677 242586 40743 242589
rect 43253 242586 43319 242589
rect 553945 242586 554011 242589
rect 40677 242584 43319 242586
rect 40677 242528 40682 242584
rect 40738 242528 43258 242584
rect 43314 242528 43319 242584
rect 40677 242526 43319 242528
rect 552460 242584 554011 242586
rect 552460 242528 553950 242584
rect 554006 242528 554011 242584
rect 552460 242526 554011 242528
rect 40677 242523 40743 242526
rect 43253 242523 43319 242526
rect 553945 242523 554011 242526
rect 671797 241498 671863 241501
rect 675109 241498 675175 241501
rect 671797 241496 675175 241498
rect 671797 241440 671802 241496
rect 671858 241440 675114 241496
rect 675170 241440 675175 241496
rect 671797 241438 675175 241440
rect 671797 241435 671863 241438
rect 675109 241435 675175 241438
rect 553853 240410 553919 240413
rect 552460 240408 553919 240410
rect 552460 240352 553858 240408
rect 553914 240352 553919 240408
rect 552460 240350 553919 240352
rect 553853 240347 553919 240350
rect 675201 240276 675267 240277
rect 675150 240274 675156 240276
rect 675110 240214 675156 240274
rect 675220 240272 675267 240276
rect 675262 240216 675267 240272
rect 675150 240212 675156 240214
rect 675220 240212 675267 240216
rect 675201 240211 675267 240212
rect 40718 240076 40724 240140
rect 40788 240138 40794 240140
rect 41781 240138 41847 240141
rect 40788 240136 41847 240138
rect 40788 240080 41786 240136
rect 41842 240080 41847 240136
rect 40788 240078 41847 240080
rect 40788 240076 40794 240078
rect 41781 240075 41847 240078
rect 42057 238506 42123 238509
rect 46933 238506 46999 238509
rect 42057 238504 46999 238506
rect 42057 238448 42062 238504
rect 42118 238448 46938 238504
rect 46994 238448 46999 238504
rect 42057 238446 46999 238448
rect 42057 238443 42123 238446
rect 46933 238443 46999 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 671521 238234 671587 238237
rect 675109 238234 675175 238237
rect 671521 238232 675175 238234
rect 671521 238176 671526 238232
rect 671582 238176 675114 238232
rect 675170 238176 675175 238232
rect 671521 238174 675175 238176
rect 671521 238171 671587 238174
rect 675109 238171 675175 238174
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42517 238098 42583 238101
rect 42076 238096 42583 238098
rect 42076 238040 42522 238096
rect 42578 238040 42583 238096
rect 42076 238038 42583 238040
rect 42076 238036 42082 238038
rect 42517 238035 42583 238038
rect 675385 236876 675451 236877
rect 675334 236874 675340 236876
rect 675294 236814 675340 236874
rect 675404 236872 675451 236876
rect 675446 236816 675451 236872
rect 675334 236812 675340 236814
rect 675404 236812 675451 236816
rect 675385 236811 675451 236812
rect 668945 236738 669011 236741
rect 673521 236738 673587 236741
rect 668945 236736 673587 236738
rect 668945 236680 668950 236736
rect 669006 236680 673526 236736
rect 673582 236680 673587 236736
rect 668945 236678 673587 236680
rect 668945 236675 669011 236678
rect 673521 236675 673587 236678
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 40534 235860 40540 235924
rect 40604 235922 40610 235924
rect 41781 235922 41847 235925
rect 40604 235920 41847 235922
rect 40604 235864 41786 235920
rect 41842 235864 41847 235920
rect 40604 235862 41847 235864
rect 40604 235860 40610 235862
rect 41781 235859 41847 235862
rect 670417 235922 670483 235925
rect 675109 235922 675175 235925
rect 670417 235920 675175 235922
rect 670417 235864 670422 235920
rect 670478 235864 675114 235920
rect 675170 235864 675175 235920
rect 670417 235862 675175 235864
rect 670417 235859 670483 235862
rect 675109 235859 675175 235862
rect 42149 235378 42215 235381
rect 45001 235378 45067 235381
rect 42149 235376 45067 235378
rect 42149 235320 42154 235376
rect 42210 235320 45006 235376
rect 45062 235320 45067 235376
rect 42149 235318 45067 235320
rect 42149 235315 42215 235318
rect 45001 235315 45067 235318
rect 674097 235242 674163 235245
rect 675661 235242 675727 235245
rect 674097 235240 675727 235242
rect 674097 235184 674102 235240
rect 674158 235184 675666 235240
rect 675722 235184 675727 235240
rect 674097 235182 675727 235184
rect 674097 235179 674163 235182
rect 675661 235179 675727 235182
rect 674465 234970 674531 234973
rect 675845 234970 675911 234973
rect 674465 234968 675911 234970
rect 674465 234912 674470 234968
rect 674526 234912 675850 234968
rect 675906 234912 675911 234968
rect 674465 234910 675911 234912
rect 674465 234907 674531 234910
rect 675845 234907 675911 234910
rect 668577 234562 668643 234565
rect 672165 234562 672231 234565
rect 668577 234560 672231 234562
rect 668577 234504 668582 234560
rect 668638 234504 672170 234560
rect 672226 234504 672231 234560
rect 668577 234502 672231 234504
rect 668577 234499 668643 234502
rect 672165 234499 672231 234502
rect 674649 234426 674715 234429
rect 675845 234426 675911 234429
rect 674649 234424 675911 234426
rect 674649 234368 674654 234424
rect 674710 234368 675850 234424
rect 675906 234368 675911 234424
rect 674649 234366 675911 234368
rect 674649 234363 674715 234366
rect 675845 234363 675911 234366
rect 42241 234154 42307 234157
rect 44357 234154 44423 234157
rect 42241 234152 44423 234154
rect 42241 234096 42246 234152
rect 42302 234096 44362 234152
rect 44418 234096 44423 234152
rect 42241 234094 44423 234096
rect 42241 234091 42307 234094
rect 44357 234091 44423 234094
rect 663241 234154 663307 234157
rect 683849 234154 683915 234157
rect 663241 234152 683915 234154
rect 663241 234096 663246 234152
rect 663302 234096 683854 234152
rect 683910 234096 683915 234152
rect 663241 234094 683915 234096
rect 663241 234091 663307 234094
rect 683849 234091 683915 234094
rect 42425 233882 42491 233885
rect 46013 233882 46079 233885
rect 554405 233882 554471 233885
rect 42425 233880 46079 233882
rect 42425 233824 42430 233880
rect 42486 233824 46018 233880
rect 46074 233824 46079 233880
rect 42425 233822 46079 233824
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 42425 233819 42491 233822
rect 46013 233819 46079 233822
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683297 233882 683363 233885
rect 658917 233880 683363 233882
rect 658917 233824 658922 233880
rect 658978 233824 683302 233880
rect 683358 233824 683363 233880
rect 658917 233822 683363 233824
rect 658917 233819 658983 233822
rect 683297 233819 683363 233822
rect 42333 233202 42399 233205
rect 44541 233202 44607 233205
rect 42333 233200 44607 233202
rect 42333 233144 42338 233200
rect 42394 233144 44546 233200
rect 44602 233144 44607 233200
rect 42333 233142 44607 233144
rect 42333 233139 42399 233142
rect 44541 233139 44607 233142
rect 673177 233202 673243 233205
rect 674230 233202 674236 233204
rect 673177 233200 674236 233202
rect 673177 233144 673182 233200
rect 673238 233144 674236 233200
rect 673177 233142 674236 233144
rect 673177 233139 673243 233142
rect 674230 233140 674236 233142
rect 674300 233140 674306 233204
rect 670141 232930 670207 232933
rect 673177 232930 673243 232933
rect 670141 232928 673243 232930
rect 670141 232872 670146 232928
rect 670202 232872 673182 232928
rect 673238 232872 673243 232928
rect 670141 232870 673243 232872
rect 670141 232867 670207 232870
rect 673177 232867 673243 232870
rect 42425 231842 42491 231845
rect 43713 231842 43779 231845
rect 42425 231840 43779 231842
rect 42425 231784 42430 231840
rect 42486 231784 43718 231840
rect 43774 231784 43779 231840
rect 42425 231782 43779 231784
rect 42425 231779 42491 231782
rect 43713 231779 43779 231782
rect 663057 231842 663123 231845
rect 675173 231842 675239 231845
rect 663057 231840 675239 231842
rect 663057 231784 663062 231840
rect 663118 231784 675178 231840
rect 675234 231784 675239 231840
rect 663057 231782 675239 231784
rect 663057 231779 663123 231782
rect 675173 231779 675239 231782
rect 640241 231434 640307 231437
rect 672165 231434 672231 231437
rect 640241 231432 672231 231434
rect 640241 231376 640246 231432
rect 640302 231376 672170 231432
rect 672226 231376 672231 231432
rect 640241 231374 672231 231376
rect 640241 231371 640307 231374
rect 672165 231371 672231 231374
rect 672993 231434 673059 231437
rect 673678 231434 673684 231436
rect 672993 231432 673684 231434
rect 672993 231376 672998 231432
rect 673054 231376 673684 231432
rect 672993 231374 673684 231376
rect 672993 231371 673059 231374
rect 673678 231372 673684 231374
rect 673748 231372 673754 231436
rect 674949 231298 675015 231301
rect 675845 231298 675911 231301
rect 674949 231296 675911 231298
rect 674949 231240 674954 231296
rect 675010 231240 675850 231296
rect 675906 231240 675911 231296
rect 674949 231238 675911 231240
rect 674949 231235 675015 231238
rect 675845 231235 675911 231238
rect 663241 231162 663307 231165
rect 674833 231162 674899 231165
rect 663241 231160 674899 231162
rect 663241 231104 663246 231160
rect 663302 231104 674838 231160
rect 674894 231104 674899 231160
rect 663241 231102 674899 231104
rect 663241 231099 663307 231102
rect 674833 231099 674899 231102
rect 665541 230890 665607 230893
rect 668117 230890 668183 230893
rect 665541 230888 668183 230890
rect 665541 230832 665546 230888
rect 665602 230832 668122 230888
rect 668178 230832 668183 230888
rect 665541 230830 668183 230832
rect 665541 230827 665607 230830
rect 668117 230827 668183 230830
rect 669405 230890 669471 230893
rect 674725 230890 674791 230893
rect 669405 230888 674791 230890
rect 669405 230832 669410 230888
rect 669466 230832 674730 230888
rect 674786 230832 674791 230888
rect 669405 230830 674791 230832
rect 669405 230827 669471 230830
rect 674725 230827 674791 230830
rect 664437 230618 664503 230621
rect 675017 230618 675083 230621
rect 664437 230616 675083 230618
rect 664437 230560 664442 230616
rect 664498 230560 675022 230616
rect 675078 230560 675083 230616
rect 664437 230558 675083 230560
rect 664437 230555 664503 230558
rect 675017 230555 675083 230558
rect 672597 230346 672663 230349
rect 673361 230348 673427 230349
rect 673126 230346 673132 230348
rect 672597 230344 673132 230346
rect 672597 230288 672602 230344
rect 672658 230288 673132 230344
rect 672597 230286 673132 230288
rect 672597 230283 672663 230286
rect 673126 230284 673132 230286
rect 673196 230284 673202 230348
rect 673310 230284 673316 230348
rect 673380 230346 673427 230348
rect 674511 230346 674577 230349
rect 676765 230346 676831 230349
rect 673380 230344 673472 230346
rect 673422 230288 673472 230344
rect 673380 230286 673472 230288
rect 674511 230344 676831 230346
rect 674511 230288 674516 230344
rect 674572 230288 676770 230344
rect 676826 230288 676831 230344
rect 674511 230286 676831 230288
rect 673380 230284 673427 230286
rect 673361 230283 673427 230284
rect 674511 230283 674577 230286
rect 676765 230283 676831 230286
rect 42149 230210 42215 230213
rect 45829 230210 45895 230213
rect 42149 230208 45895 230210
rect 42149 230152 42154 230208
rect 42210 230152 45834 230208
rect 45890 230152 45895 230208
rect 42149 230150 45895 230152
rect 42149 230147 42215 230150
rect 45829 230147 45895 230150
rect 639597 230074 639663 230077
rect 673453 230074 673519 230077
rect 639597 230072 673519 230074
rect 639597 230016 639602 230072
rect 639658 230016 673458 230072
rect 673514 230016 673519 230072
rect 639597 230014 673519 230016
rect 639597 230011 639663 230014
rect 673453 230011 673519 230014
rect 674051 230074 674117 230077
rect 675109 230074 675175 230077
rect 674051 230072 675175 230074
rect 674051 230016 674056 230072
rect 674112 230016 675114 230072
rect 675170 230016 675175 230072
rect 674051 230014 675175 230016
rect 674051 230011 674117 230014
rect 675109 230011 675175 230014
rect 103605 229802 103671 229805
rect 145649 229802 145715 229805
rect 667933 229804 667999 229805
rect 667933 229802 667980 229804
rect 103605 229800 145715 229802
rect 103605 229744 103610 229800
rect 103666 229744 145654 229800
rect 145710 229744 145715 229800
rect 103605 229742 145715 229744
rect 667888 229800 667980 229802
rect 667888 229744 667938 229800
rect 667888 229742 667980 229744
rect 103605 229739 103671 229742
rect 145649 229739 145715 229742
rect 667933 229740 667980 229742
rect 668044 229740 668050 229804
rect 668158 229740 668164 229804
rect 668228 229802 668234 229804
rect 673085 229802 673151 229805
rect 668228 229800 673151 229802
rect 668228 229744 673090 229800
rect 673146 229744 673151 229800
rect 668228 229742 673151 229744
rect 668228 229740 668234 229742
rect 667933 229739 667999 229740
rect 673085 229739 673151 229742
rect 661677 229530 661743 229533
rect 671797 229530 671863 229533
rect 661677 229528 671863 229530
rect 661677 229472 661682 229528
rect 661738 229472 671802 229528
rect 671858 229472 671863 229528
rect 661677 229470 671863 229472
rect 661677 229467 661743 229470
rect 671797 229467 671863 229470
rect 673085 229530 673151 229533
rect 675109 229530 675175 229533
rect 673085 229528 675175 229530
rect 673085 229472 673090 229528
rect 673146 229472 675114 229528
rect 675170 229472 675175 229528
rect 673085 229470 675175 229472
rect 673085 229467 673151 229470
rect 675109 229467 675175 229470
rect 42425 229394 42491 229397
rect 45553 229394 45619 229397
rect 42425 229392 45619 229394
rect 42425 229336 42430 229392
rect 42486 229336 45558 229392
rect 45614 229336 45619 229392
rect 42425 229334 45619 229336
rect 42425 229331 42491 229334
rect 45553 229331 45619 229334
rect 146293 229394 146359 229397
rect 147949 229394 148015 229397
rect 146293 229392 148015 229394
rect 146293 229336 146298 229392
rect 146354 229336 147954 229392
rect 148010 229336 148015 229392
rect 146293 229334 148015 229336
rect 146293 229331 146359 229334
rect 147949 229331 148015 229334
rect 157977 229394 158043 229397
rect 163865 229394 163931 229397
rect 157977 229392 163931 229394
rect 157977 229336 157982 229392
rect 158038 229336 163870 229392
rect 163926 229336 163931 229392
rect 157977 229334 163931 229336
rect 157977 229331 158043 229334
rect 163865 229331 163931 229334
rect 660941 229258 661007 229261
rect 668158 229258 668164 229260
rect 660941 229256 668164 229258
rect 660941 229200 660946 229256
rect 661002 229200 668164 229256
rect 660941 229198 668164 229200
rect 660941 229195 661007 229198
rect 668158 229196 668164 229198
rect 668228 229196 668234 229260
rect 673453 229122 673519 229125
rect 675109 229122 675175 229125
rect 673453 229120 675175 229122
rect 673453 229064 673458 229120
rect 673514 229064 675114 229120
rect 675170 229064 675175 229120
rect 673453 229062 675175 229064
rect 673453 229059 673519 229062
rect 675109 229059 675175 229062
rect 172421 228850 172487 228853
rect 174169 228850 174235 228853
rect 172421 228848 174235 228850
rect 172421 228792 172426 228848
rect 172482 228792 174174 228848
rect 174230 228792 174235 228848
rect 172421 228790 174235 228792
rect 172421 228787 172487 228790
rect 174169 228787 174235 228790
rect 174813 228850 174879 228853
rect 175733 228850 175799 228853
rect 174813 228848 175799 228850
rect 174813 228792 174818 228848
rect 174874 228792 175738 228848
rect 175794 228792 175799 228848
rect 174813 228790 175799 228792
rect 174813 228787 174879 228790
rect 175733 228787 175799 228790
rect 188337 228850 188403 228853
rect 190361 228850 190427 228853
rect 188337 228848 190427 228850
rect 188337 228792 188342 228848
rect 188398 228792 190366 228848
rect 190422 228792 190427 228848
rect 188337 228790 190427 228792
rect 188337 228787 188403 228790
rect 190361 228787 190427 228790
rect 673499 228850 673565 228853
rect 675109 228850 675175 228853
rect 673499 228848 675175 228850
rect 673499 228792 673504 228848
rect 673560 228792 675114 228848
rect 675170 228792 675175 228848
rect 673499 228790 675175 228792
rect 673499 228787 673565 228790
rect 675109 228787 675175 228790
rect 171133 228714 171199 228717
rect 172237 228714 172303 228717
rect 672901 228716 672967 228717
rect 672901 228714 672948 228716
rect 171133 228712 172303 228714
rect 171133 228656 171138 228712
rect 171194 228656 172242 228712
rect 172298 228656 172303 228712
rect 171133 228654 172303 228656
rect 672856 228712 672948 228714
rect 672856 228656 672906 228712
rect 672856 228654 672948 228656
rect 171133 228651 171199 228654
rect 172237 228651 172303 228654
rect 672901 228652 672948 228654
rect 673012 228652 673018 228716
rect 672901 228651 672967 228652
rect 147673 228578 147739 228581
rect 149789 228578 149855 228581
rect 147673 228576 149855 228578
rect 147673 228520 147678 228576
rect 147734 228520 149794 228576
rect 149850 228520 149855 228576
rect 147673 228518 149855 228520
rect 147673 228515 147739 228518
rect 149789 228515 149855 228518
rect 157425 228578 157491 228581
rect 158805 228578 158871 228581
rect 157425 228576 158871 228578
rect 157425 228520 157430 228576
rect 157486 228520 158810 228576
rect 158866 228520 158871 228576
rect 157425 228518 158871 228520
rect 157425 228515 157491 228518
rect 158805 228515 158871 228518
rect 673381 228578 673447 228581
rect 675150 228578 675156 228580
rect 673381 228576 675156 228578
rect 673381 228520 673386 228576
rect 673442 228520 675156 228576
rect 673381 228518 675156 228520
rect 673381 228515 673447 228518
rect 675150 228516 675156 228518
rect 675220 228516 675226 228580
rect 166625 228442 166691 228445
rect 171225 228442 171291 228445
rect 166625 228440 171291 228442
rect 166625 228384 166630 228440
rect 166686 228384 171230 228440
rect 171286 228384 171291 228440
rect 166625 228382 171291 228384
rect 166625 228379 166691 228382
rect 171225 228379 171291 228382
rect 79961 228306 80027 228309
rect 160461 228306 160527 228309
rect 79961 228304 160527 228306
rect 79961 228248 79966 228304
rect 80022 228248 160466 228304
rect 160522 228248 160527 228304
rect 79961 228246 160527 228248
rect 79961 228243 80027 228246
rect 160461 228243 160527 228246
rect 155861 228034 155927 228037
rect 157793 228034 157859 228037
rect 155861 228032 157859 228034
rect 155861 227976 155866 228032
rect 155922 227976 157798 228032
rect 157854 227976 157859 228032
rect 155861 227974 157859 227976
rect 155861 227971 155927 227974
rect 157793 227971 157859 227974
rect 133781 227898 133847 227901
rect 141325 227898 141391 227901
rect 133781 227896 141391 227898
rect 133781 227840 133786 227896
rect 133842 227840 141330 227896
rect 141386 227840 141391 227896
rect 133781 227838 141391 227840
rect 133781 227835 133847 227838
rect 141325 227835 141391 227838
rect 151905 227490 151971 227493
rect 152917 227490 152983 227493
rect 151905 227488 152983 227490
rect 151905 227432 151910 227488
rect 151966 227432 152922 227488
rect 152978 227432 152983 227488
rect 151905 227430 152983 227432
rect 151905 227427 151971 227430
rect 152917 227427 152983 227430
rect 159633 227490 159699 227493
rect 166441 227490 166507 227493
rect 159633 227488 166507 227490
rect 159633 227432 159638 227488
rect 159694 227432 166446 227488
rect 166502 227432 166507 227488
rect 159633 227430 166507 227432
rect 159633 227427 159699 227430
rect 166441 227427 166507 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 142153 227218 142219 227221
rect 143073 227218 143139 227221
rect 142153 227216 143139 227218
rect 142153 227160 142158 227216
rect 142214 227160 143078 227216
rect 143134 227160 143139 227216
rect 142153 227158 143139 227160
rect 142153 227155 142219 227158
rect 143073 227155 143139 227158
rect 150157 227218 150223 227221
rect 154573 227218 154639 227221
rect 150157 227216 154639 227218
rect 150157 227160 150162 227216
rect 150218 227160 154578 227216
rect 154634 227160 154639 227216
rect 150157 227158 154639 227160
rect 150157 227155 150223 227158
rect 154573 227155 154639 227158
rect 671061 227220 671127 227221
rect 671061 227216 671108 227220
rect 671172 227218 671178 227220
rect 671061 227160 671066 227216
rect 671061 227156 671108 227160
rect 671172 227158 671218 227218
rect 671172 227156 671178 227158
rect 671061 227155 671127 227156
rect 672257 227082 672323 227085
rect 675017 227082 675083 227085
rect 672257 227080 675083 227082
rect 672257 227024 672262 227080
rect 672318 227024 675022 227080
rect 675078 227024 675083 227080
rect 672257 227022 675083 227024
rect 672257 227019 672323 227022
rect 675017 227019 675083 227022
rect 73061 226946 73127 226949
rect 155309 226946 155375 226949
rect 73061 226944 155375 226946
rect 73061 226888 73066 226944
rect 73122 226888 155314 226944
rect 155370 226888 155375 226944
rect 73061 226886 155375 226888
rect 73061 226883 73127 226886
rect 155309 226883 155375 226886
rect 673177 226810 673243 226813
rect 675334 226810 675340 226812
rect 673177 226808 675340 226810
rect 673177 226752 673182 226808
rect 673238 226752 675340 226808
rect 673177 226750 675340 226752
rect 673177 226747 673243 226750
rect 675334 226748 675340 226750
rect 675404 226748 675410 226812
rect 42149 226674 42215 226677
rect 43345 226674 43411 226677
rect 42149 226672 43411 226674
rect 42149 226616 42154 226672
rect 42210 226616 43350 226672
rect 43406 226616 43411 226672
rect 42149 226614 43411 226616
rect 42149 226611 42215 226614
rect 43345 226611 43411 226614
rect 671061 226674 671127 226677
rect 672022 226674 672028 226676
rect 671061 226672 672028 226674
rect 671061 226616 671066 226672
rect 671122 226616 672028 226672
rect 671061 226614 672028 226616
rect 671061 226611 671127 226614
rect 672022 226612 672028 226614
rect 672092 226612 672098 226676
rect 139301 226538 139367 226541
rect 142245 226538 142311 226541
rect 139301 226536 142311 226538
rect 139301 226480 139306 226536
rect 139362 226480 142250 226536
rect 142306 226480 142311 226536
rect 139301 226478 142311 226480
rect 139301 226475 139367 226478
rect 142245 226475 142311 226478
rect 672257 226538 672323 226541
rect 673494 226538 673500 226540
rect 672257 226536 673500 226538
rect 672257 226480 672262 226536
rect 672318 226480 673500 226536
rect 672257 226478 673500 226480
rect 672257 226475 672323 226478
rect 673494 226476 673500 226478
rect 673564 226476 673570 226540
rect 652753 226402 652819 226405
rect 669405 226402 669471 226405
rect 652753 226400 669471 226402
rect 652753 226344 652758 226400
rect 652814 226344 669410 226400
rect 669466 226344 669471 226400
rect 652753 226342 669471 226344
rect 652753 226339 652819 226342
rect 669405 226339 669471 226342
rect 671654 226340 671660 226404
rect 671724 226402 671730 226404
rect 671981 226402 672047 226405
rect 671724 226400 672047 226402
rect 671724 226344 671986 226400
rect 672042 226344 672047 226400
rect 671724 226342 672047 226344
rect 671724 226340 671730 226342
rect 671981 226339 672047 226342
rect 153101 226130 153167 226133
rect 157609 226130 157675 226133
rect 153101 226128 157675 226130
rect 153101 226072 153106 226128
rect 153162 226072 157614 226128
rect 157670 226072 157675 226128
rect 153101 226070 157675 226072
rect 153101 226067 153167 226070
rect 157609 226067 157675 226070
rect 176653 226130 176719 226133
rect 180793 226130 180859 226133
rect 176653 226128 180859 226130
rect 176653 226072 176658 226128
rect 176714 226072 180798 226128
rect 180854 226072 180859 226128
rect 176653 226070 180859 226072
rect 176653 226067 176719 226070
rect 180793 226067 180859 226070
rect 181069 226130 181135 226133
rect 186037 226130 186103 226133
rect 181069 226128 186103 226130
rect 181069 226072 181074 226128
rect 181130 226072 186042 226128
rect 186098 226072 186103 226128
rect 181069 226070 186103 226072
rect 181069 226067 181135 226070
rect 186037 226067 186103 226070
rect 672022 226068 672028 226132
rect 672092 226130 672098 226132
rect 675201 226130 675267 226133
rect 672092 226128 675267 226130
rect 672092 226072 675206 226128
rect 675262 226072 675267 226128
rect 672092 226070 675267 226072
rect 672092 226068 672098 226070
rect 675201 226067 675267 226070
rect 186267 226026 186333 226031
rect 147029 225994 147095 225997
rect 152825 225994 152891 225997
rect 147029 225992 152891 225994
rect 147029 225936 147034 225992
rect 147090 225936 152830 225992
rect 152886 225936 152891 225992
rect 147029 225934 152891 225936
rect 147029 225931 147095 225934
rect 152825 225931 152891 225934
rect 170857 225994 170923 225997
rect 171225 225994 171291 225997
rect 170857 225992 171291 225994
rect 170857 225936 170862 225992
rect 170918 225936 171230 225992
rect 171286 225936 171291 225992
rect 186267 225970 186272 226026
rect 186328 225994 186333 226026
rect 187233 225994 187299 225997
rect 671797 225994 671863 225997
rect 186328 225992 187299 225994
rect 186328 225970 187238 225992
rect 186267 225965 187238 225970
rect 170857 225934 171291 225936
rect 186270 225936 187238 225965
rect 187294 225936 187299 225992
rect 186270 225934 187299 225936
rect 170857 225931 170923 225934
rect 171225 225931 171291 225934
rect 187233 225931 187299 225934
rect 659610 225992 671863 225994
rect 659610 225936 671802 225992
rect 671858 225936 671863 225992
rect 659610 225934 671863 225936
rect 166809 225858 166875 225861
rect 169845 225858 169911 225861
rect 166809 225856 169911 225858
rect 166809 225800 166814 225856
rect 166870 225800 169850 225856
rect 169906 225800 169911 225856
rect 166809 225798 169911 225800
rect 166809 225795 166875 225798
rect 169845 225795 169911 225798
rect 42425 225722 42491 225725
rect 43161 225722 43227 225725
rect 42425 225720 43227 225722
rect 42425 225664 42430 225720
rect 42486 225664 43166 225720
rect 43222 225664 43227 225720
rect 42425 225662 43227 225664
rect 42425 225659 42491 225662
rect 43161 225659 43227 225662
rect 171041 225722 171107 225725
rect 176929 225722 176995 225725
rect 171041 225720 176995 225722
rect 171041 225664 171046 225720
rect 171102 225664 176934 225720
rect 176990 225664 176995 225720
rect 171041 225662 176995 225664
rect 171041 225659 171107 225662
rect 176929 225659 176995 225662
rect 184841 225722 184907 225725
rect 186405 225722 186471 225725
rect 184841 225720 186471 225722
rect 184841 225664 184846 225720
rect 184902 225664 186410 225720
rect 186466 225664 186471 225720
rect 184841 225662 186471 225664
rect 184841 225659 184907 225662
rect 186405 225659 186471 225662
rect 143165 225586 143231 225589
rect 147397 225586 147463 225589
rect 143165 225584 147463 225586
rect 143165 225528 143170 225584
rect 143226 225528 147402 225584
rect 147458 225528 147463 225584
rect 143165 225526 147463 225528
rect 143165 225523 143231 225526
rect 147397 225523 147463 225526
rect 161565 225586 161631 225589
rect 166717 225586 166783 225589
rect 161565 225584 166783 225586
rect 161565 225528 161570 225584
rect 161626 225528 166722 225584
rect 166778 225528 166783 225584
rect 161565 225526 166783 225528
rect 161565 225523 161631 225526
rect 166717 225523 166783 225526
rect 654777 225586 654843 225589
rect 659610 225586 659670 225934
rect 671797 225931 671863 225934
rect 669405 225722 669471 225725
rect 654777 225584 659670 225586
rect 654777 225528 654782 225584
rect 654838 225528 659670 225584
rect 654777 225526 659670 225528
rect 664486 225720 669471 225722
rect 664486 225664 669410 225720
rect 669466 225664 669471 225720
rect 664486 225662 669471 225664
rect 654777 225523 654843 225526
rect 185669 225450 185735 225453
rect 186589 225450 186655 225453
rect 185669 225448 186655 225450
rect 185669 225392 185674 225448
rect 185730 225392 186594 225448
rect 186650 225392 186655 225448
rect 185669 225390 186655 225392
rect 185669 225387 185735 225390
rect 186589 225387 186655 225390
rect 186865 225450 186931 225453
rect 194869 225450 194935 225453
rect 186865 225448 194935 225450
rect 186865 225392 186870 225448
rect 186926 225392 194874 225448
rect 194930 225392 194935 225448
rect 186865 225390 194935 225392
rect 186865 225387 186931 225390
rect 194869 225387 194935 225390
rect 136541 225314 136607 225317
rect 142245 225314 142311 225317
rect 136541 225312 142311 225314
rect 136541 225256 136546 225312
rect 136602 225256 142250 225312
rect 142306 225256 142311 225312
rect 136541 225254 142311 225256
rect 136541 225251 136607 225254
rect 142245 225251 142311 225254
rect 145925 225314 145991 225317
rect 153285 225314 153351 225317
rect 145925 225312 153351 225314
rect 145925 225256 145930 225312
rect 145986 225256 153290 225312
rect 153346 225256 153351 225312
rect 145925 225254 153351 225256
rect 145925 225251 145991 225254
rect 153285 225251 153351 225254
rect 176469 225314 176535 225317
rect 176745 225314 176811 225317
rect 176469 225312 176811 225314
rect 176469 225256 176474 225312
rect 176530 225256 176750 225312
rect 176806 225256 176811 225312
rect 176469 225254 176811 225256
rect 176469 225251 176535 225254
rect 176745 225251 176811 225254
rect 655881 225314 655947 225317
rect 664486 225314 664546 225662
rect 669405 225659 669471 225662
rect 671061 225722 671127 225725
rect 674281 225722 674347 225725
rect 671061 225720 674347 225722
rect 671061 225664 671066 225720
rect 671122 225664 674286 225720
rect 674342 225664 674347 225720
rect 671061 225662 674347 225664
rect 671061 225659 671127 225662
rect 674281 225659 674347 225662
rect 671061 225450 671127 225453
rect 673499 225450 673565 225453
rect 671061 225448 673565 225450
rect 671061 225392 671066 225448
rect 671122 225392 673504 225448
rect 673560 225392 673565 225448
rect 671061 225390 673565 225392
rect 671061 225387 671127 225390
rect 673499 225387 673565 225390
rect 655881 225312 664546 225314
rect 655881 225256 655886 225312
rect 655942 225256 664546 225312
rect 655881 225254 664546 225256
rect 655881 225251 655947 225254
rect 186313 225178 186379 225181
rect 195513 225178 195579 225181
rect 186313 225176 195579 225178
rect 186313 225120 186318 225176
rect 186374 225120 195518 225176
rect 195574 225120 195579 225176
rect 186313 225118 195579 225120
rect 186313 225115 186379 225118
rect 195513 225115 195579 225118
rect 202689 225178 202755 225181
rect 205081 225178 205147 225181
rect 202689 225176 205147 225178
rect 202689 225120 202694 225176
rect 202750 225120 205086 225176
rect 205142 225120 205147 225176
rect 202689 225118 205147 225120
rect 202689 225115 202755 225118
rect 205081 225115 205147 225118
rect 673177 225178 673243 225181
rect 673678 225178 673684 225180
rect 673177 225176 673684 225178
rect 673177 225120 673182 225176
rect 673238 225120 673684 225176
rect 673177 225118 673684 225120
rect 673177 225115 673243 225118
rect 673678 225116 673684 225118
rect 673748 225116 673754 225180
rect 166533 225042 166599 225045
rect 171041 225042 171107 225045
rect 166533 225040 171107 225042
rect 166533 224984 166538 225040
rect 166594 224984 171046 225040
rect 171102 224984 171107 225040
rect 166533 224982 171107 224984
rect 166533 224979 166599 224982
rect 171041 224979 171107 224982
rect 660205 225042 660271 225045
rect 668393 225042 668459 225045
rect 660205 225040 668459 225042
rect 660205 224984 660210 225040
rect 660266 224984 668398 225040
rect 668454 224984 668459 225040
rect 660205 224982 668459 224984
rect 660205 224979 660271 224982
rect 668393 224979 668459 224982
rect 671654 224980 671660 225044
rect 671724 225042 671730 225044
rect 671981 225042 672047 225045
rect 671724 225040 672047 225042
rect 671724 224984 671986 225040
rect 672042 224984 672047 225040
rect 671724 224982 672047 224984
rect 671724 224980 671730 224982
rect 671981 224979 672047 224982
rect 672257 225040 672323 225045
rect 672257 224984 672262 225040
rect 672318 224984 672323 225040
rect 672257 224979 672323 224984
rect 672260 224773 672320 224979
rect 673494 224844 673500 224908
rect 673564 224906 673570 224908
rect 675385 224906 675451 224909
rect 673564 224904 675451 224906
rect 673564 224848 675390 224904
rect 675446 224848 675451 224904
rect 673564 224846 675451 224848
rect 673564 224844 673570 224846
rect 675385 224843 675451 224846
rect 672257 224768 672323 224773
rect 672257 224712 672262 224768
rect 672318 224712 672323 224768
rect 672257 224707 672323 224712
rect 672901 224634 672967 224637
rect 675845 224634 675911 224637
rect 672901 224632 675911 224634
rect 672901 224576 672906 224632
rect 672962 224576 675850 224632
rect 675906 224576 675911 224632
rect 672901 224574 675911 224576
rect 672901 224571 672967 224574
rect 675845 224571 675911 224574
rect 658181 224498 658247 224501
rect 670923 224498 670989 224501
rect 658181 224496 670989 224498
rect 658181 224440 658186 224496
rect 658242 224440 670928 224496
rect 670984 224440 670989 224496
rect 658181 224438 670989 224440
rect 658181 224435 658247 224438
rect 670923 224435 670989 224438
rect 152457 224362 152523 224365
rect 137970 224360 152523 224362
rect 137970 224304 152462 224360
rect 152518 224304 152523 224360
rect 137970 224302 152523 224304
rect 68921 224226 68987 224229
rect 137970 224226 138030 224302
rect 152457 224299 152523 224302
rect 157057 224362 157123 224365
rect 162945 224362 163011 224365
rect 157057 224360 163011 224362
rect 157057 224304 157062 224360
rect 157118 224304 162950 224360
rect 163006 224304 163011 224360
rect 157057 224302 163011 224304
rect 157057 224299 157123 224302
rect 162945 224299 163011 224302
rect 672717 224362 672783 224365
rect 673126 224362 673132 224364
rect 672717 224360 673132 224362
rect 672717 224304 672722 224360
rect 672778 224304 673132 224360
rect 672717 224302 673132 224304
rect 672717 224299 672783 224302
rect 673126 224300 673132 224302
rect 673196 224300 673202 224364
rect 68921 224224 138030 224226
rect 68921 224168 68926 224224
rect 68982 224168 138030 224224
rect 68921 224166 138030 224168
rect 170949 224226 171015 224229
rect 171409 224226 171475 224229
rect 170949 224224 171475 224226
rect 170949 224168 170954 224224
rect 171010 224168 171414 224224
rect 171470 224168 171475 224224
rect 170949 224166 171475 224168
rect 68921 224163 68987 224166
rect 170949 224163 171015 224166
rect 171409 224163 171475 224166
rect 145649 224090 145715 224093
rect 147765 224090 147831 224093
rect 145649 224088 147831 224090
rect 145649 224032 145654 224088
rect 145710 224032 147770 224088
rect 147826 224032 147831 224088
rect 145649 224030 147831 224032
rect 145649 224027 145715 224030
rect 147765 224027 147831 224030
rect 156689 224090 156755 224093
rect 157425 224090 157491 224093
rect 156689 224088 157491 224090
rect 156689 224032 156694 224088
rect 156750 224032 157430 224088
rect 157486 224032 157491 224088
rect 156689 224030 157491 224032
rect 156689 224027 156755 224030
rect 157425 224027 157491 224030
rect 670877 224090 670943 224093
rect 671102 224090 671108 224092
rect 670877 224088 671108 224090
rect 670877 224032 670882 224088
rect 670938 224032 671108 224088
rect 670877 224030 671108 224032
rect 670877 224027 670943 224030
rect 671102 224028 671108 224030
rect 671172 224028 671178 224092
rect 672257 224090 672323 224093
rect 673310 224090 673316 224092
rect 672257 224088 673316 224090
rect 672257 224032 672262 224088
rect 672318 224032 673316 224088
rect 672257 224030 673316 224032
rect 672257 224027 672323 224030
rect 673310 224028 673316 224030
rect 673380 224028 673386 224092
rect 140957 223954 141023 223957
rect 145373 223954 145439 223957
rect 140957 223952 145439 223954
rect 140957 223896 140962 223952
rect 141018 223896 145378 223952
rect 145434 223896 145439 223952
rect 140957 223894 145439 223896
rect 140957 223891 141023 223894
rect 145373 223891 145439 223894
rect 163957 223954 164023 223957
rect 170949 223954 171015 223957
rect 163957 223952 171015 223954
rect 163957 223896 163962 223952
rect 164018 223896 170954 223952
rect 171010 223896 171015 223952
rect 163957 223894 171015 223896
rect 163957 223891 164023 223894
rect 170949 223891 171015 223894
rect 659561 223954 659627 223957
rect 670693 223954 670759 223957
rect 659561 223952 670759 223954
rect 659561 223896 659566 223952
rect 659622 223896 670698 223952
rect 670754 223896 670759 223952
rect 659561 223894 670759 223896
rect 659561 223891 659627 223894
rect 670693 223891 670759 223894
rect 151721 223818 151787 223821
rect 157241 223818 157307 223821
rect 679249 223818 679315 223821
rect 151721 223816 157307 223818
rect 151721 223760 151726 223816
rect 151782 223760 157246 223816
rect 157302 223760 157307 223816
rect 151721 223758 157307 223760
rect 151721 223755 151787 223758
rect 157241 223755 157307 223758
rect 679206 223816 679315 223818
rect 679206 223760 679254 223816
rect 679310 223760 679315 223816
rect 679206 223755 679315 223760
rect 656617 223682 656683 223685
rect 668393 223682 668459 223685
rect 656617 223680 668459 223682
rect 656617 223624 656622 223680
rect 656678 223624 668398 223680
rect 668454 223624 668459 223680
rect 656617 223622 668459 223624
rect 656617 223619 656683 223622
rect 668393 223619 668459 223622
rect 673494 223620 673500 223684
rect 673564 223682 673570 223684
rect 673821 223682 673887 223685
rect 673564 223680 673887 223682
rect 673564 223624 673826 223680
rect 673882 223624 673887 223680
rect 673564 223622 673887 223624
rect 673564 223620 673570 223622
rect 673821 223619 673887 223622
rect 679206 223516 679266 223755
rect 157241 223410 157307 223413
rect 157425 223410 157491 223413
rect 157241 223408 157491 223410
rect 157241 223352 157246 223408
rect 157302 223352 157430 223408
rect 157486 223352 157491 223408
rect 157241 223350 157491 223352
rect 157241 223347 157307 223350
rect 157425 223347 157491 223350
rect 658917 223410 658983 223413
rect 667013 223410 667079 223413
rect 658917 223408 667079 223410
rect 658917 223352 658922 223408
rect 658978 223352 667018 223408
rect 667074 223352 667079 223408
rect 658917 223350 667079 223352
rect 658917 223347 658983 223350
rect 667013 223347 667079 223350
rect 166809 223274 166875 223277
rect 170397 223274 170463 223277
rect 166809 223272 170463 223274
rect 166809 223216 166814 223272
rect 166870 223216 170402 223272
rect 170458 223216 170463 223272
rect 166809 223214 170463 223216
rect 166809 223211 166875 223214
rect 170397 223211 170463 223214
rect 155033 223138 155099 223141
rect 157057 223138 157123 223141
rect 155033 223136 157123 223138
rect 155033 223080 155038 223136
rect 155094 223080 157062 223136
rect 157118 223080 157123 223136
rect 155033 223078 157123 223080
rect 155033 223075 155099 223078
rect 157057 223075 157123 223078
rect 158345 223138 158411 223141
rect 165797 223138 165863 223141
rect 158345 223136 165863 223138
rect 158345 223080 158350 223136
rect 158406 223080 165802 223136
rect 165858 223080 165863 223136
rect 158345 223078 165863 223080
rect 158345 223075 158411 223078
rect 165797 223075 165863 223078
rect 650637 223138 650703 223141
rect 666829 223138 666895 223141
rect 683297 223138 683363 223141
rect 650637 223136 666895 223138
rect 650637 223080 650642 223136
rect 650698 223080 666834 223136
rect 666890 223080 666895 223136
rect 650637 223078 666895 223080
rect 683284 223136 683363 223138
rect 683284 223080 683302 223136
rect 683358 223080 683363 223136
rect 683284 223078 683363 223080
rect 650637 223075 650703 223078
rect 666829 223075 666895 223078
rect 683297 223075 683363 223078
rect 40677 222866 40743 222869
rect 62941 222866 63007 222869
rect 40677 222864 63007 222866
rect 40677 222808 40682 222864
rect 40738 222808 62946 222864
rect 63002 222808 63007 222864
rect 40677 222806 63007 222808
rect 40677 222803 40743 222806
rect 62941 222803 63007 222806
rect 123385 222866 123451 222869
rect 165613 222866 165679 222869
rect 123385 222864 165679 222866
rect 123385 222808 123390 222864
rect 123446 222808 165618 222864
rect 165674 222808 165679 222864
rect 123385 222806 165679 222808
rect 123385 222803 123451 222806
rect 165613 222803 165679 222806
rect 651833 222866 651899 222869
rect 673913 222866 673979 222869
rect 651833 222864 673979 222866
rect 651833 222808 651838 222864
rect 651894 222808 673918 222864
rect 673974 222808 673979 222864
rect 651833 222806 673979 222808
rect 651833 222803 651899 222806
rect 673913 222803 673979 222806
rect 683849 222730 683915 222733
rect 683836 222728 683915 222730
rect 683836 222672 683854 222728
rect 683910 222672 683915 222728
rect 683836 222670 683915 222672
rect 683849 222667 683915 222670
rect 160829 222594 160895 222597
rect 162301 222594 162367 222597
rect 565721 222596 565787 222597
rect 160829 222592 162367 222594
rect 160829 222536 160834 222592
rect 160890 222536 162306 222592
rect 162362 222536 162367 222592
rect 160829 222534 162367 222536
rect 160829 222531 160895 222534
rect 162301 222531 162367 222534
rect 565670 222532 565676 222596
rect 565740 222594 565787 222596
rect 567377 222594 567443 222597
rect 572621 222594 572687 222597
rect 565740 222592 565832 222594
rect 565782 222536 565832 222592
rect 565740 222534 565832 222536
rect 567377 222592 572687 222594
rect 567377 222536 567382 222592
rect 567438 222536 572626 222592
rect 572682 222536 572687 222592
rect 567377 222534 572687 222536
rect 565740 222532 565787 222534
rect 565721 222531 565787 222532
rect 567377 222531 567443 222534
rect 572621 222531 572687 222534
rect 171225 222322 171291 222325
rect 176653 222322 176719 222325
rect 171225 222320 176719 222322
rect 171225 222264 171230 222320
rect 171286 222264 176658 222320
rect 176714 222264 176719 222320
rect 171225 222262 176719 222264
rect 171225 222259 171291 222262
rect 176653 222259 176719 222262
rect 562225 222322 562291 222325
rect 571885 222322 571951 222325
rect 679985 222322 680051 222325
rect 562225 222320 571951 222322
rect 562225 222264 562230 222320
rect 562286 222264 571890 222320
rect 571946 222264 571951 222320
rect 562225 222262 571951 222264
rect 679972 222320 680051 222322
rect 679972 222264 679990 222320
rect 680046 222264 680051 222320
rect 679972 222262 680051 222264
rect 562225 222259 562291 222262
rect 571885 222259 571951 222262
rect 679985 222259 680051 222262
rect 572161 222210 572227 222213
rect 572161 222208 572684 222210
rect 147305 222186 147371 222189
rect 152089 222186 152155 222189
rect 147305 222184 152155 222186
rect 147305 222128 147310 222184
rect 147366 222128 152094 222184
rect 152150 222128 152155 222184
rect 572161 222152 572166 222208
rect 572222 222186 572684 222208
rect 575933 222186 575999 222189
rect 572222 222184 575999 222186
rect 572222 222152 575938 222184
rect 572161 222150 575938 222152
rect 572161 222147 572227 222150
rect 147305 222126 152155 222128
rect 572624 222128 575938 222150
rect 575994 222128 575999 222184
rect 572624 222126 575999 222128
rect 147305 222123 147371 222126
rect 152089 222123 152155 222126
rect 575933 222123 575999 222126
rect 667013 222186 667079 222189
rect 675385 222186 675451 222189
rect 667013 222184 675451 222186
rect 667013 222128 667018 222184
rect 667074 222128 675390 222184
rect 675446 222128 675451 222184
rect 667013 222126 675451 222128
rect 667013 222123 667079 222126
rect 675385 222123 675451 222126
rect 176101 222050 176167 222053
rect 176837 222050 176903 222053
rect 176101 222048 176903 222050
rect 176101 221992 176106 222048
rect 176162 221992 176842 222048
rect 176898 221992 176903 222048
rect 176101 221990 176903 221992
rect 176101 221987 176167 221990
rect 176837 221987 176903 221990
rect 555417 222050 555483 222053
rect 562593 222050 562659 222053
rect 555417 222048 562659 222050
rect 555417 221992 555422 222048
rect 555478 221992 562598 222048
rect 562654 221992 562659 222048
rect 555417 221990 562659 221992
rect 555417 221987 555483 221990
rect 562593 221987 562659 221990
rect 563145 222050 563211 222053
rect 572478 222050 572484 222052
rect 563145 222048 572484 222050
rect 563145 221992 563150 222048
rect 563206 221992 572484 222048
rect 563145 221990 572484 221992
rect 563145 221987 563211 221990
rect 572478 221988 572484 221990
rect 572548 221988 572554 222052
rect 597461 222050 597527 222053
rect 602245 222050 602311 222053
rect 597461 222048 602311 222050
rect 597461 221992 597466 222048
rect 597522 221992 602250 222048
rect 602306 221992 602311 222048
rect 597461 221990 602311 221992
rect 597461 221987 597527 221990
rect 602245 221987 602311 221990
rect 147489 221914 147555 221917
rect 149053 221914 149119 221917
rect 147489 221912 149119 221914
rect 147489 221856 147494 221912
rect 147550 221856 149058 221912
rect 149114 221856 149119 221912
rect 147489 221854 149119 221856
rect 147489 221851 147555 221854
rect 149053 221851 149119 221854
rect 171041 221914 171107 221917
rect 171501 221914 171567 221917
rect 171041 221912 171567 221914
rect 171041 221856 171046 221912
rect 171102 221856 171506 221912
rect 171562 221856 171567 221912
rect 171041 221854 171567 221856
rect 171041 221851 171107 221854
rect 171501 221851 171567 221854
rect 674557 221914 674623 221917
rect 674557 221912 676292 221914
rect 674557 221856 674562 221912
rect 674618 221856 676292 221912
rect 674557 221854 676292 221856
rect 674557 221851 674623 221854
rect 138289 221778 138355 221781
rect 146569 221778 146635 221781
rect 138289 221776 146635 221778
rect 138289 221720 138294 221776
rect 138350 221720 146574 221776
rect 146630 221720 146635 221776
rect 138289 221718 146635 221720
rect 138289 221715 138355 221718
rect 146569 221715 146635 221718
rect 177389 221778 177455 221781
rect 185025 221778 185091 221781
rect 177389 221776 185091 221778
rect 177389 221720 177394 221776
rect 177450 221720 185030 221776
rect 185086 221720 185091 221776
rect 177389 221718 185091 221720
rect 177389 221715 177455 221718
rect 185025 221715 185091 221718
rect 517697 221778 517763 221781
rect 616873 221778 616939 221781
rect 517697 221776 616939 221778
rect 517697 221720 517702 221776
rect 517758 221720 616878 221776
rect 616934 221720 616939 221776
rect 517697 221718 616939 221720
rect 517697 221715 517763 221718
rect 616873 221715 616939 221718
rect 657997 221778 658063 221781
rect 671797 221778 671863 221781
rect 657997 221776 671863 221778
rect 657997 221720 658002 221776
rect 658058 221720 671802 221776
rect 671858 221720 671863 221776
rect 657997 221718 671863 221720
rect 657997 221715 658063 221718
rect 671797 221715 671863 221718
rect 513373 221642 513439 221645
rect 513373 221640 514770 221642
rect 513373 221584 513378 221640
rect 513434 221584 514770 221640
rect 513373 221582 514770 221584
rect 513373 221579 513439 221582
rect 101857 221506 101923 221509
rect 178033 221506 178099 221509
rect 101857 221504 178099 221506
rect 101857 221448 101862 221504
rect 101918 221448 178038 221504
rect 178094 221448 178099 221504
rect 101857 221446 178099 221448
rect 101857 221443 101923 221446
rect 178033 221443 178099 221446
rect 181253 221506 181319 221509
rect 185853 221506 185919 221509
rect 181253 221504 185919 221506
rect 181253 221448 181258 221504
rect 181314 221448 185858 221504
rect 185914 221448 185919 221504
rect 181253 221446 185919 221448
rect 514710 221506 514770 221582
rect 599485 221506 599551 221509
rect 514710 221504 599551 221506
rect 514710 221448 599490 221504
rect 599546 221448 599551 221504
rect 514710 221446 599551 221448
rect 181253 221443 181319 221446
rect 185853 221443 185919 221446
rect 599485 221443 599551 221446
rect 651189 221506 651255 221509
rect 675017 221506 675083 221509
rect 679801 221506 679867 221509
rect 651189 221504 675083 221506
rect 651189 221448 651194 221504
rect 651250 221448 675022 221504
rect 675078 221448 675083 221504
rect 651189 221446 675083 221448
rect 679788 221504 679867 221506
rect 679788 221448 679806 221504
rect 679862 221448 679867 221504
rect 679788 221446 679867 221448
rect 651189 221443 651255 221446
rect 675017 221443 675083 221446
rect 679801 221443 679867 221446
rect 142429 221234 142495 221237
rect 144177 221234 144243 221237
rect 142429 221232 144243 221234
rect 142429 221176 142434 221232
rect 142490 221176 144182 221232
rect 144238 221176 144243 221232
rect 142429 221174 144243 221176
rect 142429 221171 142495 221174
rect 144177 221171 144243 221174
rect 515765 221234 515831 221237
rect 600773 221234 600839 221237
rect 515765 221232 600839 221234
rect 515765 221176 515770 221232
rect 515826 221176 600778 221232
rect 600834 221176 600839 221232
rect 515765 221174 600839 221176
rect 515765 221171 515831 221174
rect 600773 221171 600839 221174
rect 672022 221036 672028 221100
rect 672092 221098 672098 221100
rect 672092 221038 676292 221098
rect 672092 221036 672098 221038
rect 486601 220962 486667 220965
rect 611629 220962 611695 220965
rect 486601 220960 611695 220962
rect 486601 220904 486606 220960
rect 486662 220904 611634 220960
rect 611690 220904 611695 220960
rect 486601 220902 611695 220904
rect 486601 220899 486667 220902
rect 611629 220899 611695 220902
rect 670734 220900 670740 220964
rect 670804 220962 670810 220964
rect 671797 220962 671863 220965
rect 670804 220960 671863 220962
rect 670804 220904 671802 220960
rect 671858 220904 671863 220960
rect 670804 220902 671863 220904
rect 670804 220900 670810 220902
rect 671797 220899 671863 220902
rect 150065 220826 150131 220829
rect 156137 220826 156203 220829
rect 150065 220824 156203 220826
rect 150065 220768 150070 220824
rect 150126 220768 156142 220824
rect 156198 220768 156203 220824
rect 150065 220766 156203 220768
rect 150065 220763 150131 220766
rect 156137 220763 156203 220766
rect 555601 220690 555667 220693
rect 558545 220690 558611 220693
rect 555601 220688 558611 220690
rect 555601 220632 555606 220688
rect 555662 220632 558550 220688
rect 558606 220632 558611 220688
rect 555601 220630 558611 220632
rect 555601 220627 555667 220630
rect 558545 220627 558611 220630
rect 572478 220628 572484 220692
rect 572548 220690 572554 220692
rect 577589 220690 577655 220693
rect 572548 220688 577655 220690
rect 572548 220632 577594 220688
rect 577650 220632 577655 220688
rect 572548 220630 577655 220632
rect 572548 220628 572554 220630
rect 577589 220627 577655 220630
rect 653029 220690 653095 220693
rect 673729 220690 673795 220693
rect 679617 220690 679683 220693
rect 653029 220688 673795 220690
rect 653029 220632 653034 220688
rect 653090 220632 673734 220688
rect 673790 220632 673795 220688
rect 653029 220630 673795 220632
rect 679604 220688 679683 220690
rect 679604 220632 679622 220688
rect 679678 220632 679683 220688
rect 679604 220630 679683 220632
rect 653029 220627 653095 220630
rect 673729 220627 673795 220630
rect 679617 220627 679683 220630
rect 153653 220554 153719 220557
rect 137970 220552 153719 220554
rect 137970 220496 153658 220552
rect 153714 220496 153719 220552
rect 137970 220494 153719 220496
rect 72877 220418 72943 220421
rect 137970 220418 138030 220494
rect 153653 220491 153719 220494
rect 533705 220554 533771 220557
rect 540094 220554 540100 220556
rect 533705 220552 540100 220554
rect 533705 220496 533710 220552
rect 533766 220496 540100 220552
rect 533705 220494 540100 220496
rect 533705 220491 533771 220494
rect 540094 220492 540100 220494
rect 540164 220492 540170 220556
rect 541893 220554 541959 220557
rect 544653 220554 544719 220557
rect 541893 220552 544719 220554
rect 541893 220496 541898 220552
rect 541954 220496 544658 220552
rect 544714 220496 544719 220552
rect 541893 220494 544719 220496
rect 541893 220491 541959 220494
rect 544653 220491 544719 220494
rect 547413 220554 547479 220557
rect 549069 220554 549135 220557
rect 547413 220552 549135 220554
rect 547413 220496 547418 220552
rect 547474 220496 549074 220552
rect 549130 220496 549135 220552
rect 547413 220494 549135 220496
rect 547413 220491 547479 220494
rect 549069 220491 549135 220494
rect 553485 220554 553551 220557
rect 554957 220554 555023 220557
rect 559741 220554 559807 220557
rect 553485 220552 555023 220554
rect 553485 220496 553490 220552
rect 553546 220496 554962 220552
rect 555018 220496 555023 220552
rect 558686 220552 559807 220554
rect 558686 220520 559746 220552
rect 553485 220494 555023 220496
rect 553485 220491 553551 220494
rect 554957 220491 555023 220494
rect 557950 220496 559746 220520
rect 559802 220496 559807 220552
rect 557950 220494 559807 220496
rect 557950 220460 558746 220494
rect 559741 220491 559807 220494
rect 562041 220554 562107 220557
rect 563421 220554 563487 220557
rect 562041 220552 563487 220554
rect 562041 220496 562046 220552
rect 562102 220496 563426 220552
rect 563482 220496 563487 220552
rect 562041 220494 563487 220496
rect 562041 220491 562107 220494
rect 563421 220491 563487 220494
rect 563646 220492 563652 220556
rect 563716 220554 563722 220556
rect 572345 220554 572411 220557
rect 563716 220552 572411 220554
rect 563716 220496 572350 220552
rect 572406 220496 572411 220552
rect 563716 220494 572411 220496
rect 563716 220492 563722 220494
rect 572345 220491 572411 220494
rect 674925 220554 674991 220557
rect 675845 220554 675911 220557
rect 674925 220552 675911 220554
rect 674925 220496 674930 220552
rect 674986 220496 675850 220552
rect 675906 220496 675911 220552
rect 674925 220494 675911 220496
rect 674925 220491 674991 220494
rect 675845 220491 675911 220494
rect 72877 220416 138030 220418
rect 72877 220360 72882 220416
rect 72938 220360 138030 220416
rect 72877 220358 138030 220360
rect 157333 220418 157399 220421
rect 161473 220418 161539 220421
rect 157333 220416 161539 220418
rect 157333 220360 157338 220416
rect 157394 220360 161478 220416
rect 161534 220360 161539 220416
rect 157333 220358 161539 220360
rect 72877 220355 72943 220358
rect 157333 220355 157399 220358
rect 161473 220355 161539 220358
rect 147489 220282 147555 220285
rect 148225 220282 148291 220285
rect 147489 220280 148291 220282
rect 147489 220224 147494 220280
rect 147550 220224 148230 220280
rect 148286 220224 148291 220280
rect 147489 220222 148291 220224
rect 147489 220219 147555 220222
rect 148225 220219 148291 220222
rect 519537 220282 519603 220285
rect 544193 220282 544259 220285
rect 554078 220282 554084 220284
rect 519537 220280 534090 220282
rect 519537 220224 519542 220280
rect 519598 220224 534090 220280
rect 519537 220222 534090 220224
rect 519537 220219 519603 220222
rect 69749 220146 69815 220149
rect 140773 220146 140839 220149
rect 146385 220146 146451 220149
rect 69749 220144 138030 220146
rect 69749 220088 69754 220144
rect 69810 220088 138030 220144
rect 69749 220086 138030 220088
rect 69749 220083 69815 220086
rect 137970 219874 138030 220086
rect 140773 220144 146451 220146
rect 140773 220088 140778 220144
rect 140834 220088 146390 220144
rect 146446 220088 146451 220144
rect 140773 220086 146451 220088
rect 140773 220083 140839 220086
rect 146385 220083 146451 220086
rect 510981 220012 511047 220013
rect 510981 220008 511028 220012
rect 511092 220010 511098 220012
rect 512637 220010 512703 220013
rect 526437 220012 526503 220013
rect 526437 220010 526484 220012
rect 510981 219952 510986 220008
rect 510981 219948 511028 219952
rect 511092 219950 511138 220010
rect 512637 220008 524430 220010
rect 512637 219952 512642 220008
rect 512698 219952 524430 220008
rect 512637 219950 524430 219952
rect 526392 220008 526484 220010
rect 526392 219952 526442 220008
rect 526392 219950 526484 219952
rect 511092 219948 511098 219950
rect 510981 219947 511047 219948
rect 512637 219947 512703 219950
rect 151077 219874 151143 219877
rect 137970 219872 151143 219874
rect 137970 219816 151082 219872
rect 151138 219816 151143 219872
rect 137970 219814 151143 219816
rect 151077 219811 151143 219814
rect 494789 219738 494855 219741
rect 519537 219738 519603 219741
rect 519813 219740 519879 219741
rect 522573 219740 522639 219741
rect 519813 219738 519860 219740
rect 494789 219736 519603 219738
rect 494789 219680 494794 219736
rect 494850 219680 519542 219736
rect 519598 219680 519603 219736
rect 494789 219678 519603 219680
rect 519768 219736 519860 219738
rect 519768 219680 519818 219736
rect 519768 219678 519860 219680
rect 494789 219675 494855 219678
rect 519537 219675 519603 219678
rect 519813 219676 519860 219678
rect 519924 219676 519930 219740
rect 522573 219736 522620 219740
rect 522684 219738 522690 219740
rect 524370 219738 524430 219950
rect 526437 219948 526484 219950
rect 526548 219948 526554 220012
rect 530025 220010 530091 220013
rect 533705 220010 533771 220013
rect 530025 220008 533771 220010
rect 530025 219952 530030 220008
rect 530086 219952 533710 220008
rect 533766 219952 533771 220008
rect 530025 219950 533771 219952
rect 534030 220010 534090 220222
rect 544193 220280 554084 220282
rect 544193 220224 544198 220280
rect 544254 220224 554084 220280
rect 544193 220222 554084 220224
rect 544193 220219 544259 220222
rect 554078 220220 554084 220222
rect 554148 220220 554154 220284
rect 555233 220282 555299 220285
rect 557950 220282 558010 220460
rect 643185 220418 643251 220421
rect 668393 220418 668459 220421
rect 572854 220358 582390 220418
rect 572854 220282 572914 220358
rect 555233 220280 558010 220282
rect 555233 220224 555238 220280
rect 555294 220224 558010 220280
rect 555233 220222 558010 220224
rect 558134 220222 572914 220282
rect 555233 220219 555299 220222
rect 558134 220010 558194 220222
rect 572989 220146 573055 220149
rect 582097 220146 582163 220149
rect 572989 220144 582163 220146
rect 572989 220088 572994 220144
rect 573050 220088 582102 220144
rect 582158 220088 582163 220144
rect 572989 220086 582163 220088
rect 572989 220083 573055 220086
rect 582097 220083 582163 220086
rect 582330 220010 582390 220358
rect 643185 220416 668459 220418
rect 643185 220360 643190 220416
rect 643246 220360 668398 220416
rect 668454 220360 668459 220416
rect 643185 220358 668459 220360
rect 643185 220355 643251 220358
rect 668393 220355 668459 220358
rect 670693 220418 670759 220421
rect 672809 220418 672875 220421
rect 670693 220416 672875 220418
rect 670693 220360 670698 220416
rect 670754 220360 672814 220416
rect 672870 220360 672875 220416
rect 670693 220358 672875 220360
rect 670693 220355 670759 220358
rect 672809 220355 672875 220358
rect 599025 220282 599091 220285
rect 601785 220282 601851 220285
rect 606753 220282 606819 220285
rect 599025 220280 601851 220282
rect 599025 220224 599030 220280
rect 599086 220224 601790 220280
rect 601846 220224 601851 220280
rect 599025 220222 601851 220224
rect 599025 220219 599091 220222
rect 601785 220219 601851 220222
rect 606342 220280 606819 220282
rect 606342 220224 606758 220280
rect 606814 220224 606819 220280
rect 606342 220222 606819 220224
rect 606342 220010 606402 220222
rect 606753 220219 606819 220222
rect 674373 220282 674439 220285
rect 674373 220280 676292 220282
rect 674373 220224 674378 220280
rect 674434 220224 676292 220280
rect 674373 220222 676292 220224
rect 674373 220219 674439 220222
rect 641437 220146 641503 220149
rect 641437 220144 672228 220146
rect 641437 220088 641442 220144
rect 641498 220088 672228 220144
rect 641437 220086 672228 220088
rect 641437 220083 641503 220086
rect 617057 220010 617123 220013
rect 534030 219950 558194 220010
rect 558318 219950 572914 220010
rect 582330 219950 606402 220010
rect 606526 220008 617123 220010
rect 606526 219952 617062 220008
rect 617118 219952 617123 220008
rect 606526 219950 617123 219952
rect 672168 220010 672228 220086
rect 672168 219950 674850 220010
rect 526437 219947 526503 219948
rect 530025 219947 530091 219950
rect 533705 219947 533771 219950
rect 558318 219738 558378 219950
rect 572854 219874 572914 219950
rect 572854 219814 573098 219874
rect 522573 219680 522578 219736
rect 522573 219676 522620 219680
rect 522684 219678 522730 219738
rect 524370 219678 558378 219738
rect 558545 219738 558611 219741
rect 559097 219738 559163 219741
rect 558545 219736 559163 219738
rect 558545 219680 558550 219736
rect 558606 219680 559102 219736
rect 559158 219680 559163 219736
rect 558545 219678 559163 219680
rect 522684 219676 522690 219678
rect 519813 219675 519879 219676
rect 522573 219675 522639 219676
rect 558545 219675 558611 219678
rect 559097 219675 559163 219678
rect 559373 219738 559439 219741
rect 562542 219738 562548 219740
rect 559373 219736 562548 219738
rect 559373 219680 559378 219736
rect 559434 219680 562548 219736
rect 559373 219678 562548 219680
rect 559373 219675 559439 219678
rect 562542 219676 562548 219678
rect 562612 219676 562618 219740
rect 562869 219738 562935 219741
rect 568021 219738 568087 219741
rect 562869 219736 568087 219738
rect 562869 219680 562874 219736
rect 562930 219680 568026 219736
rect 568082 219680 568087 219736
rect 562869 219678 568087 219680
rect 562869 219675 562935 219678
rect 568021 219675 568087 219678
rect 568614 219676 568620 219740
rect 568684 219738 568690 219740
rect 572161 219738 572227 219741
rect 568684 219736 572227 219738
rect 568684 219680 572166 219736
rect 572222 219680 572227 219736
rect 568684 219678 572227 219680
rect 573038 219738 573098 219814
rect 606526 219738 606586 219950
rect 617057 219947 617123 219950
rect 668393 219874 668459 219877
rect 670693 219874 670759 219877
rect 671981 219876 672047 219877
rect 671981 219874 672028 219876
rect 668393 219872 670759 219874
rect 668393 219816 668398 219872
rect 668454 219816 670698 219872
rect 670754 219816 670759 219872
rect 668393 219814 670759 219816
rect 671936 219872 672028 219874
rect 671936 219816 671986 219872
rect 671936 219814 672028 219816
rect 668393 219811 668459 219814
rect 670693 219811 670759 219814
rect 671981 219812 672028 219814
rect 672092 219812 672098 219876
rect 671981 219811 672047 219812
rect 573038 219678 606586 219738
rect 606753 219738 606819 219741
rect 630949 219738 631015 219741
rect 606753 219736 631015 219738
rect 606753 219680 606758 219736
rect 606814 219680 630954 219736
rect 631010 219680 631015 219736
rect 606753 219678 631015 219680
rect 674790 219738 674850 219950
rect 675518 219948 675524 220012
rect 675588 220010 675594 220012
rect 676029 220010 676095 220013
rect 675588 220008 676095 220010
rect 675588 219952 676034 220008
rect 676090 219952 676095 220008
rect 675588 219950 676095 219952
rect 675588 219948 675594 219950
rect 676029 219947 676095 219950
rect 683481 219874 683547 219877
rect 683468 219872 683547 219874
rect 683468 219816 683486 219872
rect 683542 219816 683547 219872
rect 683468 219814 683547 219816
rect 683481 219811 683547 219814
rect 676029 219738 676095 219741
rect 674790 219736 676095 219738
rect 674790 219680 676034 219736
rect 676090 219680 676095 219736
rect 674790 219678 676095 219680
rect 568684 219676 568690 219678
rect 572161 219675 572227 219678
rect 606753 219675 606819 219678
rect 630949 219675 631015 219678
rect 676029 219675 676095 219678
rect 147029 219466 147095 219469
rect 148041 219466 148107 219469
rect 147029 219464 148107 219466
rect 147029 219408 147034 219464
rect 147090 219408 148046 219464
rect 148102 219408 148107 219464
rect 147029 219406 148107 219408
rect 147029 219403 147095 219406
rect 148041 219403 148107 219406
rect 484577 219466 484643 219469
rect 630765 219466 630831 219469
rect 484577 219464 630831 219466
rect 484577 219408 484582 219464
rect 484638 219408 630770 219464
rect 630826 219408 630831 219464
rect 484577 219406 630831 219408
rect 484577 219403 484643 219406
rect 630765 219403 630831 219406
rect 666829 219466 666895 219469
rect 666829 219464 676292 219466
rect 666829 219408 666834 219464
rect 666890 219408 676292 219464
rect 666829 219406 676292 219408
rect 666829 219403 666895 219406
rect 195053 219330 195119 219333
rect 196065 219330 196131 219333
rect 195053 219328 196131 219330
rect 195053 219272 195058 219328
rect 195114 219272 196070 219328
rect 196126 219272 196131 219328
rect 195053 219270 196131 219272
rect 195053 219267 195119 219270
rect 196065 219267 196131 219270
rect 137829 219194 137895 219197
rect 138105 219194 138171 219197
rect 137829 219192 138171 219194
rect 137829 219136 137834 219192
rect 137890 219136 138110 219192
rect 138166 219136 138171 219192
rect 137829 219134 138171 219136
rect 137829 219131 137895 219134
rect 138105 219131 138171 219134
rect 166257 219194 166323 219197
rect 167177 219194 167243 219197
rect 166257 219192 167243 219194
rect 166257 219136 166262 219192
rect 166318 219136 167182 219192
rect 167238 219136 167243 219192
rect 166257 219134 167243 219136
rect 166257 219131 166323 219134
rect 167177 219131 167243 219134
rect 490557 219194 490623 219197
rect 491109 219194 491175 219197
rect 490557 219192 491175 219194
rect 490557 219136 490562 219192
rect 490618 219136 491114 219192
rect 491170 219136 491175 219192
rect 490557 219134 491175 219136
rect 490557 219131 490623 219134
rect 491109 219131 491175 219134
rect 492949 219194 493015 219197
rect 493593 219194 493659 219197
rect 492949 219192 493659 219194
rect 492949 219136 492954 219192
rect 493010 219136 493598 219192
rect 493654 219136 493659 219192
rect 492949 219134 493659 219136
rect 492949 219131 493015 219134
rect 493593 219131 493659 219134
rect 497733 219194 497799 219197
rect 502517 219194 502583 219197
rect 497733 219192 502583 219194
rect 497733 219136 497738 219192
rect 497794 219136 502522 219192
rect 502578 219136 502583 219192
rect 497733 219134 502583 219136
rect 497733 219131 497799 219134
rect 502517 219131 502583 219134
rect 502701 219194 502767 219197
rect 505093 219194 505159 219197
rect 502701 219192 505159 219194
rect 502701 219136 502706 219192
rect 502762 219136 505098 219192
rect 505154 219136 505159 219192
rect 502701 219134 505159 219136
rect 502701 219131 502767 219134
rect 505093 219131 505159 219134
rect 505277 219194 505343 219197
rect 514753 219194 514819 219197
rect 505277 219192 514819 219194
rect 505277 219136 505282 219192
rect 505338 219136 514758 219192
rect 514814 219136 514819 219192
rect 505277 219134 514819 219136
rect 505277 219131 505343 219134
rect 514753 219131 514819 219134
rect 514937 219194 515003 219197
rect 547597 219194 547663 219197
rect 514937 219192 547663 219194
rect 514937 219136 514942 219192
rect 514998 219136 547602 219192
rect 547658 219136 547663 219192
rect 514937 219134 547663 219136
rect 514937 219131 515003 219134
rect 547597 219131 547663 219134
rect 548149 219194 548215 219197
rect 572662 219194 572668 219196
rect 548149 219192 572668 219194
rect 548149 219136 548154 219192
rect 548210 219136 572668 219192
rect 548149 219134 572668 219136
rect 548149 219131 548215 219134
rect 572662 219132 572668 219134
rect 572732 219132 572738 219196
rect 572846 219132 572852 219196
rect 572916 219194 572922 219196
rect 582097 219194 582163 219197
rect 572916 219192 582163 219194
rect 572916 219136 582102 219192
rect 582158 219136 582163 219192
rect 572916 219134 582163 219136
rect 572916 219132 572922 219134
rect 582097 219131 582163 219134
rect 582281 219194 582347 219197
rect 586145 219194 586211 219197
rect 582281 219192 586211 219194
rect 582281 219136 582286 219192
rect 582342 219136 586150 219192
rect 586206 219136 586211 219192
rect 582281 219134 586211 219136
rect 582281 219131 582347 219134
rect 586145 219131 586211 219134
rect 586329 219194 586395 219197
rect 599761 219194 599827 219197
rect 604085 219194 604151 219197
rect 586329 219192 599827 219194
rect 586329 219136 586334 219192
rect 586390 219136 599766 219192
rect 599822 219136 599827 219192
rect 586329 219134 599827 219136
rect 586329 219131 586395 219134
rect 599761 219131 599827 219134
rect 600638 219192 604151 219194
rect 600638 219136 604090 219192
rect 604146 219136 604151 219192
rect 600638 219134 604151 219136
rect 142245 219058 142311 219061
rect 145649 219058 145715 219061
rect 142245 219056 145715 219058
rect 142245 219000 142250 219056
rect 142306 219000 145654 219056
rect 145710 219000 145715 219056
rect 142245 218998 145715 219000
rect 142245 218995 142311 218998
rect 145649 218995 145715 218998
rect 152089 218922 152155 218925
rect 153837 218922 153903 218925
rect 152089 218920 153903 218922
rect 152089 218864 152094 218920
rect 152150 218864 153842 218920
rect 153898 218864 153903 218920
rect 152089 218862 153903 218864
rect 152089 218859 152155 218862
rect 153837 218859 153903 218862
rect 166441 218922 166507 218925
rect 166993 218922 167059 218925
rect 166441 218920 167059 218922
rect 166441 218864 166446 218920
rect 166502 218864 166998 218920
rect 167054 218864 167059 218920
rect 166441 218862 167059 218864
rect 166441 218859 166507 218862
rect 166993 218859 167059 218862
rect 490281 218922 490347 218925
rect 600638 218922 600698 219134
rect 604085 219131 604151 219134
rect 638861 219194 638927 219197
rect 675293 219194 675359 219197
rect 638861 219192 675359 219194
rect 638861 219136 638866 219192
rect 638922 219136 675298 219192
rect 675354 219136 675359 219192
rect 638861 219134 675359 219136
rect 638861 219131 638927 219134
rect 675293 219131 675359 219134
rect 675661 219058 675727 219061
rect 675661 219056 676292 219058
rect 675661 219000 675666 219056
rect 675722 219000 676292 219056
rect 675661 218998 676292 219000
rect 675661 218995 675727 218998
rect 490281 218920 572684 218922
rect 490281 218864 490286 218920
rect 490342 218888 572684 218920
rect 572808 218888 600698 218922
rect 490342 218864 600698 218888
rect 490281 218862 600698 218864
rect 600957 218922 601023 218925
rect 640057 218922 640123 218925
rect 675518 218922 675524 218924
rect 600957 218920 615510 218922
rect 600957 218864 600962 218920
rect 601018 218864 615510 218920
rect 600957 218862 615510 218864
rect 490281 218859 490347 218862
rect 572624 218828 572868 218862
rect 600957 218859 601023 218862
rect 147489 218786 147555 218789
rect 148593 218786 148659 218789
rect 147489 218784 148659 218786
rect 147489 218728 147494 218784
rect 147550 218728 148598 218784
rect 148654 218728 148659 218784
rect 147489 218726 148659 218728
rect 147489 218723 147555 218726
rect 148593 218723 148659 218726
rect 157241 218650 157307 218653
rect 157701 218650 157767 218653
rect 157241 218648 157767 218650
rect 157241 218592 157246 218648
rect 157302 218592 157706 218648
rect 157762 218592 157767 218648
rect 157241 218590 157767 218592
rect 157241 218587 157307 218590
rect 157701 218587 157767 218590
rect 166533 218650 166599 218653
rect 167177 218650 167243 218653
rect 166533 218648 167243 218650
rect 166533 218592 166538 218648
rect 166594 218592 167182 218648
rect 167238 218592 167243 218648
rect 166533 218590 167243 218592
rect 166533 218587 166599 218590
rect 167177 218587 167243 218590
rect 491109 218650 491175 218653
rect 504817 218650 504883 218653
rect 491109 218648 504883 218650
rect 491109 218592 491114 218648
rect 491170 218592 504822 218648
rect 504878 218592 504883 218648
rect 491109 218590 504883 218592
rect 491109 218587 491175 218590
rect 504817 218587 504883 218590
rect 505001 218650 505067 218653
rect 510153 218650 510219 218653
rect 548149 218650 548215 218653
rect 505001 218648 509986 218650
rect 505001 218592 505006 218648
rect 505062 218592 509986 218648
rect 505001 218590 509986 218592
rect 505001 218587 505067 218590
rect 166257 218378 166323 218381
rect 167361 218378 167427 218381
rect 166257 218376 167427 218378
rect 166257 218320 166262 218376
rect 166318 218320 167366 218376
rect 167422 218320 167427 218376
rect 166257 218318 167427 218320
rect 166257 218315 166323 218318
rect 167361 218315 167427 218318
rect 496905 218378 496971 218381
rect 500033 218378 500099 218381
rect 496905 218376 500099 218378
rect 496905 218320 496910 218376
rect 496966 218320 500038 218376
rect 500094 218320 500099 218376
rect 496905 218318 500099 218320
rect 496905 218315 496971 218318
rect 500033 218315 500099 218318
rect 500217 218378 500283 218381
rect 504633 218378 504699 218381
rect 500217 218376 504699 218378
rect 500217 218320 500222 218376
rect 500278 218320 504638 218376
rect 504694 218320 504699 218376
rect 500217 218318 504699 218320
rect 500217 218315 500283 218318
rect 504633 218315 504699 218318
rect 505277 218378 505343 218381
rect 509693 218378 509759 218381
rect 505277 218376 509759 218378
rect 505277 218320 505282 218376
rect 505338 218320 509698 218376
rect 509754 218320 509759 218376
rect 505277 218318 509759 218320
rect 509926 218378 509986 218590
rect 510153 218648 548215 218650
rect 510153 218592 510158 218648
rect 510214 218592 548154 218648
rect 548210 218592 548215 218648
rect 510153 218590 548215 218592
rect 510153 218587 510219 218590
rect 548149 218587 548215 218590
rect 548566 218590 562794 218650
rect 548566 218378 548626 218590
rect 509926 218318 548626 218378
rect 549253 218378 549319 218381
rect 553669 218378 553735 218381
rect 549253 218376 553735 218378
rect 549253 218320 549258 218376
rect 549314 218320 553674 218376
rect 553730 218320 553735 218376
rect 549253 218318 553735 218320
rect 505277 218315 505343 218318
rect 509693 218315 509759 218318
rect 549253 218315 549319 218318
rect 553669 218315 553735 218318
rect 554037 218378 554103 218381
rect 562174 218378 562180 218380
rect 554037 218376 562180 218378
rect 554037 218320 554042 218376
rect 554098 218320 562180 218376
rect 554037 218318 562180 218320
rect 554037 218315 554103 218318
rect 562174 218316 562180 218318
rect 562244 218316 562250 218380
rect 562734 218378 562794 218590
rect 562910 218588 562916 218652
rect 562980 218650 562986 218652
rect 572621 218650 572687 218653
rect 562980 218648 572687 218650
rect 562980 218592 572626 218648
rect 572682 218592 572687 218648
rect 562980 218590 572687 218592
rect 562980 218588 562986 218590
rect 572621 218587 572687 218590
rect 582327 218650 582393 218653
rect 614481 218650 614547 218653
rect 582327 218648 614547 218650
rect 582327 218592 582332 218648
rect 582388 218592 614486 218648
rect 614542 218592 614547 218648
rect 582327 218590 614547 218592
rect 615450 218650 615510 218862
rect 640057 218920 675524 218922
rect 640057 218864 640062 218920
rect 640118 218864 675524 218920
rect 640057 218862 675524 218864
rect 640057 218859 640123 218862
rect 675518 218860 675524 218862
rect 675588 218860 675594 218924
rect 631133 218650 631199 218653
rect 615450 218648 631199 218650
rect 615450 218592 631138 218648
rect 631194 218592 631199 218648
rect 615450 218590 631199 218592
rect 582327 218587 582393 218590
rect 614481 218587 614547 218590
rect 631133 218587 631199 218590
rect 649901 218650 649967 218653
rect 674741 218650 674807 218653
rect 649901 218648 674807 218650
rect 649901 218592 649906 218648
rect 649962 218592 674746 218648
rect 674802 218592 674807 218648
rect 649901 218590 674807 218592
rect 649901 218587 649967 218590
rect 674741 218587 674807 218590
rect 674966 218588 674972 218652
rect 675036 218650 675042 218652
rect 675036 218590 676292 218650
rect 675036 218588 675042 218590
rect 572805 218514 572871 218517
rect 582189 218514 582255 218517
rect 572805 218512 582255 218514
rect 572805 218456 572810 218512
rect 572866 218456 582194 218512
rect 582250 218456 582255 218512
rect 572805 218454 582255 218456
rect 572805 218451 572871 218454
rect 582189 218451 582255 218454
rect 586513 218378 586579 218381
rect 600957 218378 601023 218381
rect 562734 218344 572500 218378
rect 586513 218376 601023 218378
rect 574737 218344 574803 218347
rect 562734 218342 574803 218344
rect 562734 218318 574742 218342
rect 572440 218286 574742 218318
rect 574798 218286 574803 218342
rect 586513 218320 586518 218376
rect 586574 218320 600962 218376
rect 601018 218320 601023 218376
rect 586513 218318 601023 218320
rect 586513 218315 586579 218318
rect 600957 218315 601023 218318
rect 601141 218378 601207 218381
rect 629937 218378 630003 218381
rect 601141 218376 630003 218378
rect 601141 218320 601146 218376
rect 601202 218320 629942 218376
rect 629998 218320 630003 218376
rect 601141 218318 630003 218320
rect 601141 218315 601207 218318
rect 629937 218315 630003 218318
rect 572440 218284 574803 218286
rect 574737 218281 574803 218284
rect 571241 218208 571307 218211
rect 571241 218206 572362 218208
rect 571241 218150 571246 218206
rect 571302 218150 572362 218206
rect 575054 218180 575060 218244
rect 575124 218242 575130 218244
rect 586329 218242 586395 218245
rect 575124 218240 586395 218242
rect 575124 218184 586334 218240
rect 586390 218184 586395 218240
rect 575124 218182 586395 218184
rect 575124 218180 575130 218182
rect 586329 218179 586395 218182
rect 675886 218180 675892 218244
rect 675956 218242 675962 218244
rect 675956 218182 676292 218242
rect 675956 218180 675962 218182
rect 571241 218148 572362 218150
rect 571241 218145 571307 218148
rect 487797 218106 487863 218109
rect 562869 218106 562935 218109
rect 487797 218104 562935 218106
rect 487797 218048 487802 218104
rect 487858 218048 562874 218104
rect 562930 218048 562935 218104
rect 487797 218046 562935 218048
rect 572302 218106 572362 218148
rect 574461 218106 574527 218109
rect 572302 218104 574527 218106
rect 572302 218048 574466 218104
rect 574522 218048 574527 218104
rect 572302 218046 574527 218048
rect 487797 218043 487863 218046
rect 562869 218043 562935 218046
rect 574461 218043 574527 218046
rect 586513 218106 586579 218109
rect 626441 218106 626507 218109
rect 586513 218104 626507 218106
rect 586513 218048 586518 218104
rect 586574 218048 626446 218104
rect 626502 218048 626507 218104
rect 586513 218046 626507 218048
rect 586513 218043 586579 218046
rect 626441 218043 626507 218046
rect 35525 217970 35591 217973
rect 54477 217970 54543 217973
rect 35525 217968 54543 217970
rect 35525 217912 35530 217968
rect 35586 217912 54482 217968
rect 54538 217912 54543 217968
rect 35525 217910 54543 217912
rect 35525 217907 35591 217910
rect 54477 217907 54543 217910
rect 563278 217908 563284 217972
rect 563348 217970 563354 217972
rect 572161 217970 572227 217973
rect 563348 217968 572227 217970
rect 563348 217912 572166 217968
rect 572222 217912 572227 217968
rect 563348 217910 572227 217912
rect 563348 217908 563354 217910
rect 572161 217907 572227 217910
rect 498653 217834 498719 217837
rect 504817 217834 504883 217837
rect 505829 217834 505895 217837
rect 498653 217832 504650 217834
rect 498653 217776 498658 217832
rect 498714 217776 504650 217832
rect 498653 217774 504650 217776
rect 498653 217771 498719 217774
rect 503529 217562 503595 217565
rect 504398 217562 504404 217564
rect 503529 217560 504404 217562
rect 503529 217504 503534 217560
rect 503590 217504 504404 217560
rect 503529 217502 504404 217504
rect 503529 217499 503595 217502
rect 504398 217500 504404 217502
rect 504468 217500 504474 217564
rect 504590 217562 504650 217774
rect 504817 217832 505895 217834
rect 504817 217776 504822 217832
rect 504878 217776 505834 217832
rect 505890 217776 505895 217832
rect 504817 217774 505895 217776
rect 504817 217771 504883 217774
rect 505829 217771 505895 217774
rect 506013 217834 506079 217837
rect 508262 217834 508268 217836
rect 506013 217832 508268 217834
rect 506013 217776 506018 217832
rect 506074 217776 508268 217832
rect 506013 217774 508268 217776
rect 506013 217771 506079 217774
rect 508262 217772 508268 217774
rect 508332 217772 508338 217836
rect 508497 217834 508563 217837
rect 533613 217834 533679 217837
rect 562726 217834 562732 217836
rect 508497 217832 533679 217834
rect 508497 217776 508502 217832
rect 508558 217776 533618 217832
rect 533674 217776 533679 217832
rect 508497 217774 533679 217776
rect 508497 217771 508563 217774
rect 533613 217771 533679 217774
rect 534214 217774 562732 217834
rect 534214 217562 534274 217774
rect 562726 217772 562732 217774
rect 562796 217772 562802 217836
rect 591481 217834 591547 217837
rect 572302 217832 591547 217834
rect 572302 217776 591486 217832
rect 591542 217776 591547 217832
rect 572302 217774 591547 217776
rect 563237 217698 563303 217701
rect 572302 217698 572362 217774
rect 591481 217771 591547 217774
rect 591665 217834 591731 217837
rect 601141 217834 601207 217837
rect 591665 217832 601207 217834
rect 591665 217776 591670 217832
rect 591726 217776 601146 217832
rect 601202 217776 601207 217832
rect 591665 217774 601207 217776
rect 591665 217771 591731 217774
rect 601141 217771 601207 217774
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 563237 217696 572362 217698
rect 563237 217640 563242 217696
rect 563298 217640 572362 217696
rect 563237 217638 572362 217640
rect 563237 217635 563303 217638
rect 504590 217502 534274 217562
rect 534441 217562 534507 217565
rect 563094 217562 563100 217564
rect 534441 217560 563100 217562
rect 534441 217504 534446 217560
rect 534502 217504 563100 217560
rect 534441 217502 563100 217504
rect 534441 217499 534507 217502
rect 563094 217500 563100 217502
rect 563164 217500 563170 217564
rect 572437 217562 572503 217565
rect 574277 217562 574343 217565
rect 572437 217560 574343 217562
rect 572437 217504 572442 217560
rect 572498 217504 574282 217560
rect 574338 217504 574343 217560
rect 572437 217502 574343 217504
rect 572437 217499 572503 217502
rect 574277 217499 574343 217502
rect 574921 217562 574987 217565
rect 591021 217562 591087 217565
rect 597921 217562 597987 217565
rect 574921 217560 591087 217562
rect 574921 217504 574926 217560
rect 574982 217504 591026 217560
rect 591082 217504 591087 217560
rect 574921 217502 591087 217504
rect 574921 217499 574987 217502
rect 591021 217499 591087 217502
rect 591254 217560 597987 217562
rect 591254 217504 597926 217560
rect 597982 217504 597987 217560
rect 591254 217502 597987 217504
rect 565997 217460 566063 217463
rect 567694 217460 567700 217462
rect 565997 217458 567700 217460
rect 565675 217428 565741 217429
rect 565670 217364 565676 217428
rect 565740 217426 565746 217428
rect 565740 217366 565832 217426
rect 565997 217402 566002 217458
rect 566058 217402 567700 217458
rect 565997 217400 567700 217402
rect 565997 217397 566063 217400
rect 567694 217398 567700 217400
rect 567764 217398 567770 217462
rect 565740 217364 565746 217366
rect 565675 217363 565741 217364
rect 493593 217292 493659 217293
rect 493542 217290 493548 217292
rect 493502 217230 493548 217290
rect 493612 217288 493659 217292
rect 493654 217232 493659 217288
rect 493542 217228 493548 217230
rect 493612 217228 493659 217232
rect 493593 217227 493659 217228
rect 497549 217290 497615 217293
rect 590837 217290 590903 217293
rect 497549 217288 565554 217290
rect 497549 217232 497554 217288
rect 497610 217232 565554 217288
rect 497549 217230 565554 217232
rect 497549 217227 497615 217230
rect 565494 217188 565554 217230
rect 565908 217288 590903 217290
rect 565908 217232 590842 217288
rect 590898 217232 590903 217288
rect 565908 217230 590903 217232
rect 492121 217154 492187 217157
rect 565494 217154 565738 217188
rect 565908 217154 565968 217230
rect 590837 217227 590903 217230
rect 492121 217152 492506 217154
rect 492121 217096 492126 217152
rect 492182 217096 492506 217152
rect 565494 217128 565968 217154
rect 492121 217094 492506 217096
rect 565678 217094 565968 217128
rect 492121 217091 492187 217094
rect 492446 216746 492506 217094
rect 508262 216956 508268 217020
rect 508332 217018 508338 217020
rect 591254 217018 591314 217502
rect 597921 217499 597987 217502
rect 644933 217562 644999 217565
rect 674925 217562 674991 217565
rect 644933 217560 674991 217562
rect 644933 217504 644938 217560
rect 644994 217504 674930 217560
rect 674986 217504 674991 217560
rect 644933 217502 674991 217504
rect 644933 217499 644999 217502
rect 674925 217499 674991 217502
rect 675518 217364 675524 217428
rect 675588 217426 675594 217428
rect 675588 217366 676292 217426
rect 675588 217364 675594 217366
rect 591481 217290 591547 217293
rect 598473 217290 598539 217293
rect 591481 217288 598539 217290
rect 591481 217232 591486 217288
rect 591542 217232 598478 217288
rect 598534 217232 598539 217288
rect 591481 217230 598539 217232
rect 591481 217227 591547 217230
rect 598473 217227 598539 217230
rect 642081 217290 642147 217293
rect 675150 217290 675156 217292
rect 642081 217288 675156 217290
rect 642081 217232 642086 217288
rect 642142 217232 675156 217288
rect 642081 217230 675156 217232
rect 642081 217227 642147 217230
rect 675150 217228 675156 217230
rect 675220 217228 675226 217292
rect 508332 216958 565554 217018
rect 508332 216956 508338 216958
rect 565494 216882 565554 216958
rect 566046 216958 591314 217018
rect 592033 217018 592099 217021
rect 595161 217018 595227 217021
rect 592033 217016 595227 217018
rect 592033 216960 592038 217016
rect 592094 216960 595166 217016
rect 595222 216960 595227 217016
rect 592033 216958 595227 216960
rect 566046 216882 566106 216958
rect 592033 216955 592099 216958
rect 595161 216955 595227 216958
rect 675702 216956 675708 217020
rect 675772 217018 675778 217020
rect 675772 216958 676292 217018
rect 675772 216956 675778 216958
rect 565494 216822 566106 216882
rect 674925 216882 674991 216885
rect 675334 216882 675340 216884
rect 674925 216880 675340 216882
rect 674925 216824 674930 216880
rect 674986 216824 675340 216880
rect 674925 216822 675340 216824
rect 674925 216819 674991 216822
rect 675334 216820 675340 216822
rect 675404 216820 675410 216884
rect 590837 216746 590903 216749
rect 492446 216686 565370 216746
rect 565310 216610 565370 216686
rect 566230 216744 590903 216746
rect 566230 216688 590842 216744
rect 590898 216688 590903 216744
rect 566230 216686 590903 216688
rect 566230 216610 566290 216686
rect 590837 216683 590903 216686
rect 591021 216746 591087 216749
rect 595621 216746 595687 216749
rect 591021 216744 595687 216746
rect 591021 216688 591026 216744
rect 591082 216688 595626 216744
rect 595682 216688 595687 216744
rect 591021 216686 595687 216688
rect 591021 216683 591087 216686
rect 595621 216683 595687 216686
rect 595805 216746 595871 216749
rect 595805 216744 596190 216746
rect 595805 216688 595810 216744
rect 595866 216688 596190 216744
rect 595805 216686 596190 216688
rect 595805 216683 595871 216686
rect 565310 216550 566290 216610
rect 596130 216610 596190 216686
rect 597553 216610 597619 216613
rect 596130 216608 597619 216610
rect 596130 216552 597558 216608
rect 597614 216552 597619 216608
rect 596130 216550 597619 216552
rect 597553 216547 597619 216550
rect 674741 216610 674807 216613
rect 674741 216608 676292 216610
rect 674741 216552 674746 216608
rect 674802 216552 676292 216608
rect 674741 216550 676292 216552
rect 674741 216547 674807 216550
rect 519302 216474 519308 216476
rect 509926 216414 519308 216474
rect 504398 216140 504404 216204
rect 504468 216202 504474 216204
rect 509926 216202 509986 216414
rect 519302 216412 519308 216414
rect 519372 216412 519378 216476
rect 519854 216412 519860 216476
rect 519924 216474 519930 216476
rect 564934 216474 564940 216476
rect 519924 216414 564940 216474
rect 519924 216412 519930 216414
rect 564934 216412 564940 216414
rect 565004 216412 565010 216476
rect 566590 216412 566596 216476
rect 566660 216474 566666 216476
rect 595989 216474 596055 216477
rect 566660 216472 596055 216474
rect 566660 216416 595994 216472
rect 596050 216416 596055 216472
rect 566660 216414 596055 216416
rect 566660 216412 566666 216414
rect 595989 216411 596055 216414
rect 655421 216474 655487 216477
rect 669405 216474 669471 216477
rect 655421 216472 669471 216474
rect 655421 216416 655426 216472
rect 655482 216416 669410 216472
rect 669466 216416 669471 216472
rect 655421 216414 669471 216416
rect 655421 216411 655487 216414
rect 669405 216411 669471 216414
rect 504468 216142 509986 216202
rect 504468 216140 504474 216142
rect 511022 216140 511028 216204
rect 511092 216202 511098 216204
rect 599025 216202 599091 216205
rect 511092 216200 599091 216202
rect 511092 216144 599030 216200
rect 599086 216144 599091 216200
rect 511092 216142 599091 216144
rect 511092 216140 511098 216142
rect 599025 216139 599091 216142
rect 600957 216202 601023 216205
rect 673361 216202 673427 216205
rect 600957 216200 615510 216202
rect 600957 216144 600962 216200
rect 601018 216144 615510 216200
rect 600957 216142 615510 216144
rect 600957 216139 601023 216142
rect 519302 215868 519308 215932
rect 519372 215930 519378 215932
rect 536046 215930 536052 215932
rect 519372 215870 536052 215930
rect 519372 215868 519378 215870
rect 536046 215868 536052 215870
rect 536116 215868 536122 215932
rect 537158 215870 572730 215930
rect 522614 215596 522620 215660
rect 522684 215658 522690 215660
rect 537158 215658 537218 215870
rect 546718 215658 546724 215660
rect 522684 215598 537218 215658
rect 539366 215598 546724 215658
rect 522684 215596 522690 215598
rect 538806 215522 538812 215524
rect 537342 215462 538812 215522
rect 526478 215324 526484 215388
rect 526548 215386 526554 215388
rect 537342 215386 537402 215462
rect 538806 215460 538812 215462
rect 538876 215460 538882 215524
rect 539174 215460 539180 215524
rect 539244 215522 539250 215524
rect 539366 215522 539426 215598
rect 546718 215596 546724 215598
rect 546788 215596 546794 215660
rect 547638 215596 547644 215660
rect 547708 215658 547714 215660
rect 548190 215658 548196 215660
rect 547708 215598 548196 215658
rect 547708 215596 547714 215598
rect 548190 215596 548196 215598
rect 548260 215596 548266 215660
rect 548374 215596 548380 215660
rect 548444 215658 548450 215660
rect 556470 215658 556476 215660
rect 548444 215598 556476 215658
rect 548444 215596 548450 215598
rect 556470 215596 556476 215598
rect 556540 215596 556546 215660
rect 558862 215596 558868 215660
rect 558932 215658 558938 215660
rect 566406 215658 566412 215660
rect 558932 215598 566412 215658
rect 558932 215596 558938 215598
rect 566406 215596 566412 215598
rect 566476 215596 566482 215660
rect 572478 215658 572484 215660
rect 566598 215598 572484 215658
rect 539244 215462 539426 215522
rect 546910 215462 547338 215522
rect 539244 215460 539250 215462
rect 526548 215326 537402 215386
rect 526548 215324 526554 215326
rect 539910 215324 539916 215388
rect 539980 215386 539986 215388
rect 546910 215386 546970 215462
rect 539980 215326 546970 215386
rect 547278 215386 547338 215462
rect 556846 215462 558608 215522
rect 547278 215326 555664 215386
rect 539980 215324 539986 215326
rect 555604 215310 555664 215326
rect 556846 215310 556906 215462
rect 558548 215386 558608 215462
rect 566598 215386 566658 215598
rect 572478 215596 572484 215598
rect 572548 215596 572554 215660
rect 572670 215658 572730 215870
rect 572846 215868 572852 215932
rect 572916 215930 572922 215932
rect 582097 215930 582163 215933
rect 572916 215928 582163 215930
rect 572916 215872 582102 215928
rect 582158 215872 582163 215928
rect 572916 215870 582163 215872
rect 572916 215868 572922 215870
rect 582097 215867 582163 215870
rect 583702 215868 583708 215932
rect 583772 215930 583778 215932
rect 611353 215930 611419 215933
rect 583772 215928 611419 215930
rect 583772 215872 611358 215928
rect 611414 215872 611419 215928
rect 583772 215870 611419 215872
rect 615450 215930 615510 216142
rect 673361 216200 676292 216202
rect 673361 216144 673366 216200
rect 673422 216144 676292 216200
rect 673361 216142 676292 216144
rect 673361 216139 673427 216142
rect 620553 215930 620619 215933
rect 615450 215928 620619 215930
rect 615450 215872 620558 215928
rect 620614 215872 620619 215928
rect 615450 215870 620619 215872
rect 583772 215868 583778 215870
rect 611353 215867 611419 215870
rect 620553 215867 620619 215870
rect 643001 215930 643067 215933
rect 674925 215930 674991 215933
rect 643001 215928 674991 215930
rect 643001 215872 643006 215928
rect 643062 215872 674930 215928
rect 674986 215872 674991 215928
rect 643001 215870 674991 215872
rect 643001 215867 643067 215870
rect 674925 215867 674991 215870
rect 675293 215794 675359 215797
rect 675293 215792 676292 215794
rect 675293 215736 675298 215792
rect 675354 215736 676292 215792
rect 675293 215734 676292 215736
rect 675293 215731 675359 215734
rect 618897 215658 618963 215661
rect 572670 215656 618963 215658
rect 572670 215600 618902 215656
rect 618958 215600 618963 215656
rect 572670 215598 618963 215600
rect 618897 215595 618963 215598
rect 646589 215658 646655 215661
rect 675109 215658 675175 215661
rect 646589 215656 675175 215658
rect 646589 215600 646594 215656
rect 646650 215600 675114 215656
rect 675170 215600 675175 215656
rect 646589 215598 675175 215600
rect 646589 215595 646655 215598
rect 675109 215595 675175 215598
rect 567878 215386 567884 215388
rect 558548 215326 566658 215386
rect 566782 215326 567884 215386
rect 555604 215250 556906 215310
rect 536046 215052 536052 215116
rect 536116 215114 536122 215116
rect 538990 215114 538996 215116
rect 536116 215054 538996 215114
rect 536116 215052 536122 215054
rect 538990 215052 538996 215054
rect 539060 215052 539066 215116
rect 540094 215052 540100 215116
rect 540164 215114 540170 215116
rect 546902 215114 546908 215116
rect 540164 215054 546908 215114
rect 540164 215052 540170 215054
rect 546902 215052 546908 215054
rect 546972 215052 546978 215116
rect 548190 215052 548196 215116
rect 548260 215114 548266 215116
rect 566782 215114 566842 215326
rect 567878 215324 567884 215326
rect 567948 215324 567954 215388
rect 568070 215326 576594 215386
rect 548260 215054 566842 215114
rect 548260 215052 548266 215054
rect 566958 215052 566964 215116
rect 567028 215114 567034 215116
rect 568070 215114 568130 215326
rect 567028 215054 568130 215114
rect 567028 215052 567034 215054
rect 568246 215052 568252 215116
rect 568316 215114 568322 215116
rect 575473 215114 575539 215117
rect 568316 215112 575539 215114
rect 568316 215056 575478 215112
rect 575534 215056 575539 215112
rect 568316 215054 575539 215056
rect 576534 215114 576594 215326
rect 576710 215324 576716 215388
rect 576780 215386 576786 215388
rect 586697 215386 586763 215389
rect 595805 215386 595871 215389
rect 576780 215326 586530 215386
rect 576780 215324 576786 215326
rect 576853 215114 576919 215117
rect 576534 215112 576919 215114
rect 576534 215056 576858 215112
rect 576914 215056 576919 215112
rect 576534 215054 576919 215056
rect 586470 215114 586530 215326
rect 586697 215384 595871 215386
rect 586697 215328 586702 215384
rect 586758 215328 595810 215384
rect 595866 215328 595871 215384
rect 586697 215326 595871 215328
rect 586697 215323 586763 215326
rect 595805 215323 595871 215326
rect 595989 215386 596055 215389
rect 600957 215386 601023 215389
rect 595989 215384 601023 215386
rect 595989 215328 595994 215384
rect 596050 215328 600962 215384
rect 601018 215328 601023 215384
rect 595989 215326 601023 215328
rect 595989 215323 596055 215326
rect 600957 215323 601023 215326
rect 666461 215386 666527 215389
rect 666461 215384 676292 215386
rect 666461 215328 666466 215384
rect 666522 215328 676292 215384
rect 666461 215326 676292 215328
rect 666461 215323 666527 215326
rect 595713 215114 595779 215117
rect 586470 215112 595779 215114
rect 586470 215056 595718 215112
rect 595774 215056 595779 215112
rect 586470 215054 595779 215056
rect 568316 215052 568322 215054
rect 575473 215051 575539 215054
rect 576853 215051 576919 215054
rect 595713 215051 595779 215054
rect 664621 215114 664687 215117
rect 675845 215114 675911 215117
rect 664621 215112 675911 215114
rect 664621 215056 664626 215112
rect 664682 215056 675850 215112
rect 675906 215056 675911 215112
rect 676070 215086 676076 215150
rect 676140 215114 676146 215150
rect 676140 215086 676230 215114
rect 664621 215054 675911 215056
rect 676078 215054 676230 215086
rect 664621 215051 664687 215054
rect 675845 215051 675911 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 41492 214918 44883 214920
rect 44817 214915 44883 214918
rect 575606 214916 575612 214980
rect 575676 214978 575682 214980
rect 576301 214978 576367 214981
rect 575676 214976 576367 214978
rect 575676 214920 576306 214976
rect 576362 214920 576367 214976
rect 575676 214918 576367 214920
rect 676170 214978 676230 215054
rect 676170 214918 676292 214978
rect 575676 214916 575682 214918
rect 576301 214915 576367 214918
rect 651005 214842 651071 214845
rect 672165 214842 672231 214845
rect 651005 214840 672231 214842
rect 651005 214784 651010 214840
rect 651066 214784 672170 214840
rect 672226 214784 672231 214840
rect 651005 214782 672231 214784
rect 651005 214779 651071 214782
rect 672165 214779 672231 214782
rect 672717 214706 672783 214709
rect 673126 214706 673132 214708
rect 672717 214704 673132 214706
rect 672717 214648 672722 214704
rect 672778 214648 673132 214704
rect 672717 214646 673132 214648
rect 672717 214643 672783 214646
rect 673126 214644 673132 214646
rect 673196 214644 673202 214708
rect 647141 214570 647207 214573
rect 667013 214570 667079 214573
rect 647141 214568 667079 214570
rect 35758 214301 35818 214540
rect 647141 214512 647146 214568
rect 647202 214512 667018 214568
rect 667074 214512 667079 214568
rect 647141 214510 667079 214512
rect 647141 214507 647207 214510
rect 667013 214507 667079 214510
rect 675886 214508 675892 214572
rect 675956 214570 675962 214572
rect 675956 214510 676292 214570
rect 675956 214508 675962 214510
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 35574 214132 35634 214235
rect 575982 214026 576042 214404
rect 669405 214162 669471 214165
rect 669405 214160 676292 214162
rect 669405 214104 669410 214160
rect 669466 214104 676292 214160
rect 669405 214102 676292 214104
rect 669405 214099 669471 214102
rect 578601 214026 578667 214029
rect 575982 214024 578667 214026
rect 575982 213968 578606 214024
rect 578662 213968 578667 214024
rect 575982 213966 578667 213968
rect 578601 213963 578667 213966
rect 43529 213754 43595 213757
rect 41492 213752 43595 213754
rect 41492 213696 43534 213752
rect 43590 213696 43595 213752
rect 41492 213694 43595 213696
rect 43529 213691 43595 213694
rect 664805 213754 664871 213757
rect 672073 213754 672139 213757
rect 664805 213752 671906 213754
rect 664805 213696 664810 213752
rect 664866 213696 671906 213752
rect 664805 213694 671906 213696
rect 664805 213691 664871 213694
rect 661493 213482 661559 213485
rect 671846 213482 671906 213694
rect 672073 213752 676292 213754
rect 672073 213696 672078 213752
rect 672134 213696 676292 213752
rect 672073 213694 676292 213696
rect 672073 213691 672139 213694
rect 675845 213482 675911 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 671846 213480 675911 213482
rect 671846 213424 675850 213480
rect 675906 213424 675911 213480
rect 671846 213422 675911 213424
rect 661493 213419 661559 213422
rect 45001 213346 45067 213349
rect 41492 213344 45067 213346
rect 41492 213288 45006 213344
rect 45062 213288 45067 213344
rect 41492 213286 45067 213288
rect 45001 213283 45067 213286
rect 642173 213210 642239 213213
rect 669270 213210 669330 213422
rect 675845 213419 675911 213422
rect 683297 213346 683363 213349
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 683297 213283 683363 213286
rect 675845 213210 675911 213213
rect 642173 213208 663810 213210
rect 642173 213152 642178 213208
rect 642234 213152 663810 213208
rect 642173 213150 663810 213152
rect 669270 213208 675911 213210
rect 669270 213152 675850 213208
rect 675906 213152 675911 213208
rect 669270 213150 675911 213152
rect 642173 213147 642239 213150
rect 42977 212938 43043 212941
rect 41492 212936 43043 212938
rect 41492 212880 42982 212936
rect 43038 212880 43043 212936
rect 41492 212878 43043 212880
rect 663750 212938 663810 213150
rect 675845 213147 675911 213150
rect 673545 212938 673611 212941
rect 663750 212936 673611 212938
rect 663750 212880 673550 212936
rect 673606 212880 673611 212936
rect 663750 212878 673611 212880
rect 42977 212875 43043 212878
rect 673545 212875 673611 212878
rect 675017 212938 675083 212941
rect 675661 212938 675727 212941
rect 675017 212936 675727 212938
rect 675017 212880 675022 212936
rect 675078 212880 675666 212936
rect 675722 212880 675727 212936
rect 675017 212878 675727 212880
rect 675017 212875 675083 212878
rect 675661 212875 675727 212878
rect 683070 212533 683130 212908
rect 47945 212530 48011 212533
rect 41492 212528 48011 212530
rect 41492 212472 47950 212528
rect 48006 212472 48011 212528
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 41492 212470 48011 212472
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 47945 212467 48011 212470
rect 683113 212467 683179 212470
rect 42793 212122 42859 212125
rect 41492 212120 42859 212122
rect 41492 212064 42798 212120
rect 42854 212064 42859 212120
rect 41492 212062 42859 212064
rect 42793 212059 42859 212062
rect 575982 211714 576042 212228
rect 674046 212060 674052 212124
rect 674116 212122 674122 212124
rect 674116 212062 676292 212122
rect 674116 212060 674122 212062
rect 579429 211714 579495 211717
rect 575982 211712 579495 211714
rect 35758 211445 35818 211684
rect 575982 211656 579434 211712
rect 579490 211656 579495 211712
rect 575982 211654 579495 211656
rect 579429 211651 579495 211654
rect 35758 211440 35867 211445
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211382 35867 211384
rect 35801 211379 35867 211382
rect 675886 211380 675892 211444
rect 675956 211442 675962 211444
rect 676438 211442 676444 211444
rect 675956 211382 676444 211442
rect 675956 211380 675962 211382
rect 676438 211380 676444 211382
rect 676508 211380 676514 211444
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 44173 211243 44239 211246
rect 669446 211108 669452 211172
rect 669516 211170 669522 211172
rect 670601 211170 670667 211173
rect 683113 211170 683179 211173
rect 669516 211168 670667 211170
rect 669516 211112 670606 211168
rect 670662 211112 670667 211168
rect 669516 211110 670667 211112
rect 669516 211108 669522 211110
rect 670601 211107 670667 211110
rect 670926 211168 683179 211170
rect 670926 211112 683118 211168
rect 683174 211112 683179 211168
rect 670926 211110 683179 211112
rect 43253 210898 43319 210901
rect 41492 210896 43319 210898
rect 41492 210840 43258 210896
rect 43314 210840 43319 210896
rect 41492 210838 43319 210840
rect 43253 210835 43319 210838
rect 670601 210898 670667 210901
rect 670926 210898 670986 211110
rect 683113 211107 683179 211110
rect 670601 210896 670986 210898
rect 670601 210840 670606 210896
rect 670662 210840 670986 210896
rect 670601 210838 670986 210840
rect 670601 210835 670667 210838
rect 44173 210490 44239 210493
rect 41492 210488 44239 210490
rect 41492 210432 44178 210488
rect 44234 210432 44239 210488
rect 41492 210430 44239 210432
rect 44173 210427 44239 210430
rect 674966 210428 674972 210492
rect 675036 210490 675042 210492
rect 675886 210490 675892 210492
rect 675036 210430 675892 210490
rect 675036 210428 675042 210430
rect 675886 210428 675892 210430
rect 675956 210428 675962 210492
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 41462 209812 41522 210052
rect 575982 209946 576042 210052
rect 578785 209946 578851 209949
rect 575982 209944 578851 209946
rect 575982 209888 578790 209944
rect 578846 209888 578851 209944
rect 575982 209886 578851 209888
rect 578785 209883 578851 209886
rect 672901 209946 672967 209949
rect 678930 209946 678990 210294
rect 683297 210291 683363 210294
rect 672901 209944 678990 209946
rect 672901 209888 672906 209944
rect 672962 209888 678990 209944
rect 672901 209886 678990 209888
rect 672901 209883 672967 209886
rect 41454 209748 41460 209812
rect 41524 209748 41530 209812
rect 673913 209674 673979 209677
rect 676857 209674 676923 209677
rect 673913 209672 676923 209674
rect 41278 209402 41338 209644
rect 673913 209616 673918 209672
rect 673974 209616 676862 209672
rect 676918 209616 676923 209672
rect 673913 209614 676923 209616
rect 673913 209611 673979 209614
rect 676857 209611 676923 209614
rect 42793 209402 42859 209405
rect 41278 209400 42859 209402
rect 41278 209344 42798 209400
rect 42854 209344 42859 209400
rect 41278 209342 42859 209344
rect 42793 209339 42859 209342
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 41689 208994 41755 208997
rect 49325 208994 49391 208997
rect 41689 208992 49391 208994
rect 41689 208936 41694 208992
rect 41750 208936 49330 208992
rect 49386 208936 49391 208992
rect 41689 208934 49391 208936
rect 41689 208931 41755 208934
rect 49325 208931 49391 208934
rect 41462 208586 41522 208828
rect 44357 208586 44423 208589
rect 41462 208584 44423 208586
rect 41462 208528 44362 208584
rect 44418 208528 44423 208584
rect 41462 208526 44423 208528
rect 44357 208523 44423 208526
rect 40726 208180 40786 208420
rect 40718 208116 40724 208180
rect 40788 208116 40794 208180
rect 43437 208042 43503 208045
rect 41492 208040 43503 208042
rect 41492 207984 43442 208040
rect 43498 207984 43503 208040
rect 41492 207982 43503 207984
rect 43437 207979 43503 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40033 207770 40099 207773
rect 42006 207770 42012 207772
rect 40033 207768 42012 207770
rect 40033 207712 40038 207768
rect 40094 207712 42012 207768
rect 40033 207710 42012 207712
rect 40033 207707 40099 207710
rect 42006 207708 42012 207710
rect 42076 207708 42082 207772
rect 40910 207364 40970 207604
rect 40902 207300 40908 207364
rect 40972 207300 40978 207364
rect 575982 207362 576042 207876
rect 579429 207362 579495 207365
rect 575982 207360 579495 207362
rect 575982 207304 579434 207360
rect 579490 207304 579495 207360
rect 575982 207302 579495 207304
rect 579429 207299 579495 207302
rect 676121 207226 676187 207229
rect 669270 207224 676187 207226
rect 40542 206956 40602 207196
rect 666326 207090 666386 207196
rect 669270 207168 676126 207224
rect 676182 207168 676187 207224
rect 669270 207166 676187 207168
rect 669270 207090 669330 207166
rect 676121 207163 676187 207166
rect 666326 207030 669330 207090
rect 40534 206892 40540 206956
rect 40604 206892 40610 206956
rect 673545 206954 673611 206957
rect 677777 206954 677843 206957
rect 673545 206952 677843 206954
rect 673545 206896 673550 206952
rect 673606 206896 677782 206952
rect 677838 206896 677843 206952
rect 673545 206894 677843 206896
rect 673545 206891 673611 206894
rect 677777 206891 677843 206894
rect 43989 206818 44055 206821
rect 41492 206816 44055 206818
rect 41492 206760 43994 206816
rect 44050 206760 44055 206816
rect 41492 206758 44055 206760
rect 43989 206755 44055 206758
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 43253 206274 43319 206277
rect 49509 206274 49575 206277
rect 43253 206272 49575 206274
rect 43253 206216 43258 206272
rect 43314 206216 49514 206272
rect 49570 206216 49575 206272
rect 43253 206214 49575 206216
rect 43253 206211 43319 206214
rect 49509 206211 49575 206214
rect 44541 206002 44607 206005
rect 41492 206000 44607 206002
rect 41492 205944 44546 206000
rect 44602 205944 44607 206000
rect 41492 205942 44607 205944
rect 44541 205939 44607 205942
rect 578233 205866 578299 205869
rect 575798 205864 578299 205866
rect 575798 205808 578238 205864
rect 578294 205808 578299 205864
rect 575798 205806 578299 205808
rect 575798 205700 575858 205806
rect 578233 205803 578299 205806
rect 43805 205594 43871 205597
rect 41492 205592 43871 205594
rect 41492 205536 43810 205592
rect 43866 205536 43871 205592
rect 41492 205534 43871 205536
rect 43805 205531 43871 205534
rect 675753 205594 675819 205597
rect 676622 205594 676628 205596
rect 675753 205592 676628 205594
rect 675753 205536 675758 205592
rect 675814 205536 676628 205592
rect 675753 205534 676628 205536
rect 675753 205531 675819 205534
rect 676622 205532 676628 205534
rect 676692 205532 676698 205596
rect 43621 205186 43687 205189
rect 41492 205184 43687 205186
rect 41492 205128 43626 205184
rect 43682 205128 43687 205184
rect 41492 205126 43687 205128
rect 43621 205123 43687 205126
rect 674741 205050 674807 205053
rect 675477 205050 675543 205053
rect 674741 205048 675543 205050
rect 674741 204992 674746 205048
rect 674802 204992 675482 205048
rect 675538 204992 675543 205048
rect 674741 204990 675543 204992
rect 674741 204987 674807 204990
rect 675477 204987 675543 204990
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 35574 204101 35634 204340
rect 35574 204096 35683 204101
rect 35574 204040 35622 204096
rect 35678 204040 35683 204096
rect 35574 204038 35683 204040
rect 35617 204035 35683 204038
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 41462 203282 41522 203524
rect 50705 203282 50771 203285
rect 41462 203280 50771 203282
rect 41462 203224 50710 203280
rect 50766 203224 50771 203280
rect 41462 203222 50771 203224
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 666326 203282 666386 203932
rect 673913 203282 673979 203285
rect 666326 203280 673979 203282
rect 666326 203224 673918 203280
rect 673974 203224 673979 203280
rect 666326 203222 673979 203224
rect 50705 203219 50771 203222
rect 578325 203219 578391 203222
rect 673913 203219 673979 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 674833 202738 674899 202741
rect 675385 202738 675451 202741
rect 674833 202736 675451 202738
rect 674833 202680 674838 202736
rect 674894 202680 675390 202736
rect 675446 202680 675451 202736
rect 674833 202678 675451 202680
rect 674833 202675 674899 202678
rect 675385 202675 675451 202678
rect 35617 202194 35683 202197
rect 43437 202194 43503 202197
rect 35617 202192 43503 202194
rect 35617 202136 35622 202192
rect 35678 202136 43442 202192
rect 43498 202136 43503 202192
rect 35617 202134 43503 202136
rect 35617 202131 35683 202134
rect 43437 202131 43503 202134
rect 666326 201650 666386 202300
rect 673361 201922 673427 201925
rect 675477 201922 675543 201925
rect 673361 201920 675543 201922
rect 673361 201864 673366 201920
rect 673422 201864 675482 201920
rect 675538 201864 675543 201920
rect 673361 201862 675543 201864
rect 673361 201859 673427 201862
rect 675477 201859 675543 201862
rect 673545 201650 673611 201653
rect 666326 201648 673611 201650
rect 666326 201592 673550 201648
rect 673606 201592 673611 201648
rect 666326 201590 673611 201592
rect 673545 201587 673611 201590
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 575982 200834 576042 201348
rect 666461 200970 666527 200973
rect 675017 200970 675083 200973
rect 666461 200968 675083 200970
rect 666461 200912 666466 200968
rect 666522 200912 675022 200968
rect 675078 200912 675083 200968
rect 666461 200910 675083 200912
rect 666461 200907 666527 200910
rect 675017 200907 675083 200910
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672073 200698 672139 200701
rect 675201 200698 675267 200701
rect 672073 200696 675267 200698
rect 672073 200640 672078 200696
rect 672134 200640 675206 200696
rect 675262 200640 675267 200696
rect 672073 200638 675267 200640
rect 672073 200635 672139 200638
rect 675201 200635 675267 200638
rect 675753 200698 675819 200701
rect 676438 200698 676444 200700
rect 675753 200696 676444 200698
rect 675753 200640 675758 200696
rect 675814 200640 676444 200696
rect 675753 200638 676444 200640
rect 675753 200635 675819 200638
rect 676438 200636 676444 200638
rect 676508 200636 676514 200700
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 575982 198930 576042 199172
rect 669313 199066 669379 199069
rect 666356 199064 669379 199066
rect 666356 199008 669318 199064
rect 669374 199008 669379 199064
rect 666356 199006 669379 199008
rect 669313 199003 669379 199006
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 590377 198250 590443 198253
rect 675569 198252 675635 198253
rect 675518 198250 675524 198252
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 675478 198190 675524 198250
rect 675588 198248 675635 198252
rect 675630 198192 675635 198248
rect 590377 198187 590443 198190
rect 675518 198188 675524 198190
rect 675588 198188 675635 198192
rect 675569 198187 675635 198188
rect 37917 197842 37983 197845
rect 41822 197842 41828 197844
rect 37917 197840 41828 197842
rect 37917 197784 37922 197840
rect 37978 197784 41828 197840
rect 37917 197782 41828 197784
rect 37917 197779 37983 197782
rect 41822 197780 41828 197782
rect 41892 197780 41898 197844
rect 669129 197434 669195 197437
rect 666356 197432 669195 197434
rect 666356 197376 669134 197432
rect 669190 197376 669195 197432
rect 666356 197374 669195 197376
rect 669129 197371 669195 197374
rect 40718 197100 40724 197164
rect 40788 197162 40794 197164
rect 41781 197162 41847 197165
rect 40788 197160 41847 197162
rect 40788 197104 41786 197160
rect 41842 197104 41847 197160
rect 40788 197102 41847 197104
rect 40788 197100 40794 197102
rect 41781 197099 41847 197102
rect 669405 197162 669471 197165
rect 675385 197162 675451 197165
rect 669405 197160 675451 197162
rect 669405 197104 669410 197160
rect 669466 197104 675390 197160
rect 675446 197104 675451 197160
rect 669405 197102 675451 197104
rect 669405 197099 669471 197102
rect 675385 197099 675451 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49325 196482 49391 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49325 196480 52164 196482
rect 49325 196424 49330 196480
rect 49386 196424 52164 196480
rect 49325 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49325 196419 49391 196422
rect 578509 196419 578575 196422
rect 669221 196074 669287 196077
rect 672257 196074 672323 196077
rect 669221 196072 672323 196074
rect 669221 196016 669226 196072
rect 669282 196016 672262 196072
rect 672318 196016 672323 196072
rect 669221 196014 672323 196016
rect 669221 196011 669287 196014
rect 672257 196011 672323 196014
rect 41873 195804 41939 195805
rect 41822 195802 41828 195804
rect 41782 195742 41828 195802
rect 41892 195800 41939 195804
rect 41934 195744 41939 195800
rect 41822 195740 41828 195742
rect 41892 195740 41939 195744
rect 41873 195739 41939 195740
rect 40902 195468 40908 195532
rect 40972 195530 40978 195532
rect 42609 195530 42675 195533
rect 40972 195528 42675 195530
rect 40972 195472 42614 195528
rect 42670 195472 42675 195528
rect 40972 195470 42675 195472
rect 40972 195468 40978 195470
rect 42609 195467 42675 195470
rect 41454 195196 41460 195260
rect 41524 195258 41530 195260
rect 41781 195258 41847 195261
rect 41524 195256 41847 195258
rect 41524 195200 41786 195256
rect 41842 195200 41847 195256
rect 41524 195198 41847 195200
rect 41524 195196 41530 195198
rect 41781 195195 41847 195198
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 40534 194516 40540 194580
rect 40604 194578 40610 194580
rect 41638 194578 41644 194580
rect 40604 194518 41644 194578
rect 40604 194516 40610 194518
rect 41638 194516 41644 194518
rect 41708 194516 41714 194580
rect 49509 194442 49575 194445
rect 49509 194440 52164 194442
rect 49509 194384 49514 194440
rect 49570 194384 52164 194440
rect 49509 194382 52164 194384
rect 49509 194379 49575 194382
rect 669405 194170 669471 194173
rect 666356 194168 669471 194170
rect 666356 194112 669410 194168
rect 669466 194112 669471 194168
rect 666356 194110 669471 194112
rect 669405 194107 669471 194110
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42425 193218 42491 193221
rect 43989 193218 44055 193221
rect 42425 193216 44055 193218
rect 42425 193160 42430 193216
rect 42486 193160 43994 193216
rect 44050 193160 44055 193216
rect 42425 193158 44055 193160
rect 42425 193155 42491 193158
rect 43989 193155 44055 193158
rect 675661 193218 675727 193221
rect 675886 193218 675892 193220
rect 675661 193216 675892 193218
rect 675661 193160 675666 193216
rect 675722 193160 675892 193216
rect 675661 193158 675892 193160
rect 675661 193155 675727 193158
rect 675886 193156 675892 193158
rect 675956 193156 675962 193220
rect 42374 192884 42380 192948
rect 42444 192946 42450 192948
rect 42609 192946 42675 192949
rect 42444 192944 42675 192946
rect 42444 192888 42614 192944
rect 42670 192888 42675 192944
rect 42444 192886 42675 192888
rect 42444 192884 42450 192886
rect 42609 192883 42675 192886
rect 47945 192402 48011 192405
rect 47945 192400 52164 192402
rect 47945 192344 47950 192400
rect 48006 192344 52164 192400
rect 47945 192342 52164 192344
rect 47945 192339 48011 192342
rect 575982 192266 576042 192644
rect 667933 192538 667999 192541
rect 666356 192536 667999 192538
rect 666356 192480 667938 192536
rect 667994 192480 667999 192536
rect 666356 192478 667999 192480
rect 667933 192475 667999 192478
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 43621 191722 43687 191725
rect 42333 191720 43687 191722
rect 42333 191664 42338 191720
rect 42394 191664 43626 191720
rect 43682 191664 43687 191720
rect 42333 191662 43687 191664
rect 42333 191659 42399 191662
rect 43621 191659 43687 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43805 190498 43871 190501
rect 42425 190496 43871 190498
rect 42425 190440 42430 190496
rect 42486 190440 43810 190496
rect 43866 190440 43871 190496
rect 42425 190438 43871 190440
rect 42425 190435 42491 190438
rect 43805 190435 43871 190438
rect 48773 190498 48839 190501
rect 48773 190496 52164 190498
rect 48773 190440 48778 190496
rect 48834 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 48773 190438 52164 190440
rect 48773 190435 48839 190438
rect 670601 190362 670667 190365
rect 675293 190362 675359 190365
rect 670601 190360 675359 190362
rect 670601 190304 670606 190360
rect 670662 190304 675298 190360
rect 675354 190304 675359 190360
rect 670601 190302 675359 190304
rect 670601 190299 670667 190302
rect 675293 190299 675359 190302
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 44357 189954 44423 189957
rect 42425 189952 44423 189954
rect 42425 189896 42430 189952
rect 42486 189896 44362 189952
rect 44418 189896 44423 189952
rect 42425 189894 44423 189896
rect 42425 189891 42491 189894
rect 44357 189891 44423 189894
rect 667933 189274 667999 189277
rect 666356 189272 667999 189274
rect 666356 189216 667938 189272
rect 667994 189216 667999 189272
rect 666356 189214 667999 189216
rect 667933 189211 667999 189214
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 44541 187642 44607 187645
rect 669221 187642 669287 187645
rect 42425 187640 44607 187642
rect 42425 187584 42430 187640
rect 42486 187584 44546 187640
rect 44602 187584 44607 187640
rect 42425 187582 44607 187584
rect 666356 187640 669287 187642
rect 666356 187584 669226 187640
rect 669282 187584 669287 187640
rect 666356 187582 669287 187584
rect 42425 187579 42491 187582
rect 44541 187579 44607 187582
rect 669221 187579 669287 187582
rect 41781 187236 41847 187237
rect 41781 187232 41828 187236
rect 41892 187234 41898 187236
rect 41781 187176 41786 187232
rect 41781 187172 41828 187176
rect 41892 187174 41938 187234
rect 41892 187172 41898 187174
rect 41781 187171 41847 187172
rect 666185 186962 666251 186965
rect 683113 186962 683179 186965
rect 666185 186960 683179 186962
rect 666185 186904 666190 186960
rect 666246 186904 683118 186960
rect 683174 186904 683179 186960
rect 666185 186902 683179 186904
rect 666185 186899 666251 186902
rect 683113 186899 683179 186902
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 42333 186148 42399 186149
rect 42333 186146 42380 186148
rect 42288 186144 42380 186146
rect 42288 186088 42338 186144
rect 42288 186086 42380 186088
rect 42333 186084 42380 186086
rect 42444 186084 42450 186148
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 42333 186083 42399 186084
rect 41965 185876 42031 185877
rect 41965 185872 42012 185876
rect 42076 185874 42082 185876
rect 41965 185816 41970 185872
rect 41965 185812 42012 185816
rect 42076 185814 42122 185874
rect 42076 185812 42082 185814
rect 41965 185811 42031 185812
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 42425 184922 42491 184925
rect 44173 184922 44239 184925
rect 42425 184920 44239 184922
rect 42425 184864 42430 184920
rect 42486 184864 44178 184920
rect 44234 184864 44239 184920
rect 42425 184862 44239 184864
rect 42425 184859 42491 184862
rect 44173 184859 44239 184862
rect 579521 184378 579587 184381
rect 669221 184378 669287 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 666356 184376 669287 184378
rect 666356 184320 669226 184376
rect 669282 184320 669287 184376
rect 666356 184318 669287 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 669221 184315 669287 184318
rect 589457 183562 589523 183565
rect 672073 183562 672139 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672073 183560 672948 183562
rect 672073 183504 672078 183560
rect 672134 183504 672948 183560
rect 672073 183502 672948 183504
rect 589457 183499 589523 183502
rect 672073 183499 672139 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 43253 183154 43319 183157
rect 42425 183152 43319 183154
rect 42425 183096 42430 183152
rect 42486 183096 43258 183152
rect 43314 183096 43319 183152
rect 42425 183094 43319 183096
rect 42425 183091 42491 183094
rect 43253 183091 43319 183094
rect 668117 182746 668183 182749
rect 666356 182744 668183 182746
rect 666356 182688 668122 182744
rect 668178 182688 668183 182744
rect 666356 182686 668183 182688
rect 668117 182683 668183 182686
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667381 181386 667447 181389
rect 676489 181386 676555 181389
rect 667381 181384 676555 181386
rect 667381 181328 667386 181384
rect 667442 181328 676494 181384
rect 676550 181328 676555 181384
rect 667381 181326 676555 181328
rect 667381 181323 667447 181326
rect 676489 181323 676555 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 674097 179482 674163 179485
rect 666356 179480 674163 179482
rect 666356 179424 674102 179480
rect 674158 179424 674163 179480
rect 666356 179422 674163 179424
rect 674097 179419 674163 179422
rect 667749 178802 667815 178805
rect 683113 178802 683179 178805
rect 667749 178800 675770 178802
rect 667749 178744 667754 178800
rect 667810 178744 675770 178800
rect 667749 178742 675770 178744
rect 667749 178739 667815 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 675710 177986 675770 178742
rect 683070 178800 683179 178802
rect 683070 178744 683118 178800
rect 683174 178744 683179 178800
rect 683070 178739 683179 178744
rect 683070 178500 683130 178739
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 675710 177926 675954 177986
rect 672441 177850 672507 177853
rect 666356 177848 672507 177850
rect 666356 177792 672446 177848
rect 672502 177792 672507 177848
rect 666356 177790 672507 177792
rect 672441 177787 672507 177790
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 675894 177714 675954 177926
rect 675894 177654 676292 177714
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 674557 177306 674623 177309
rect 674557 177304 676292 177306
rect 674557 177248 674562 177304
rect 674618 177248 676292 177304
rect 674557 177246 676292 177248
rect 674557 177243 674623 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 674189 176898 674255 176901
rect 674189 176896 676292 176898
rect 674189 176840 674194 176896
rect 674250 176840 676292 176896
rect 674189 176838 676292 176840
rect 674189 176835 674255 176838
rect 671889 176490 671955 176493
rect 671889 176488 676292 176490
rect 671889 176432 671894 176488
rect 671950 176432 676292 176488
rect 671889 176430 676292 176432
rect 671889 176427 671955 176430
rect 674649 176082 674715 176085
rect 674649 176080 676292 176082
rect 674649 176024 674654 176080
rect 674710 176024 676292 176080
rect 674649 176022 676292 176024
rect 674649 176019 674715 176022
rect 674373 175674 674439 175677
rect 674373 175672 676292 175674
rect 674373 175616 674378 175672
rect 674434 175616 676292 175672
rect 674373 175614 676292 175616
rect 674373 175611 674439 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 672533 175266 672599 175269
rect 672533 175264 676292 175266
rect 575982 175130 576042 175236
rect 672533 175208 672538 175264
rect 672594 175208 676292 175264
rect 672533 175206 676292 175208
rect 672533 175203 672599 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 666829 174858 666895 174861
rect 666829 174856 676292 174858
rect 666829 174800 666834 174856
rect 666890 174800 676292 174856
rect 666829 174798 676292 174800
rect 666829 174795 666895 174798
rect 667933 174586 667999 174589
rect 666356 174584 667999 174586
rect 666356 174528 667938 174584
rect 667994 174528 667999 174584
rect 666356 174526 667999 174528
rect 667933 174523 667999 174526
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 678237 173226 678303 173229
rect 678237 173224 678316 173226
rect 678237 173168 678242 173224
rect 678298 173168 678316 173224
rect 678237 173166 678316 173168
rect 678237 173163 678303 173166
rect 673085 172954 673151 172957
rect 666356 172952 673151 172954
rect 666356 172896 673090 172952
rect 673146 172896 673151 172952
rect 666356 172894 673151 172896
rect 673085 172891 673151 172894
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 675886 171940 675892 172004
rect 675956 172002 675962 172004
rect 675956 171942 676292 172002
rect 675956 171940 675962 171942
rect 680997 171594 681063 171597
rect 680997 171592 681076 171594
rect 680997 171536 681002 171592
rect 681058 171536 681076 171592
rect 680997 171534 681076 171536
rect 680997 171531 681063 171534
rect 679617 171186 679683 171189
rect 679604 171184 679683 171186
rect 679604 171128 679622 171184
rect 679678 171128 679683 171184
rect 679604 171126 679683 171128
rect 679617 171123 679683 171126
rect 579521 171050 579587 171053
rect 575798 171048 579587 171050
rect 575798 170992 579526 171048
rect 579582 170992 579587 171048
rect 575798 170990 579587 170992
rect 575798 170884 575858 170990
rect 579521 170987 579587 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589457 170506 589523 170509
rect 589457 170504 592572 170506
rect 589457 170448 589462 170504
rect 589518 170448 592572 170504
rect 589457 170446 592572 170448
rect 589457 170443 589523 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 673177 169962 673243 169965
rect 673177 169960 676292 169962
rect 673177 169904 673182 169960
rect 673238 169904 676292 169960
rect 673177 169902 676292 169904
rect 673177 169899 673243 169902
rect 668025 169690 668091 169693
rect 666356 169688 668091 169690
rect 666356 169632 668030 169688
rect 668086 169632 668091 169688
rect 666356 169630 668091 169632
rect 668025 169627 668091 169630
rect 674373 169554 674439 169557
rect 674373 169552 676292 169554
rect 674373 169496 674378 169552
rect 674434 169496 676292 169552
rect 674373 169494 676292 169496
rect 674373 169491 674439 169494
rect 578325 169282 578391 169285
rect 575798 169280 578391 169282
rect 575798 169224 578330 169280
rect 578386 169224 578391 169280
rect 575798 169222 578391 169224
rect 575798 168708 575858 169222
rect 578325 169219 578391 169222
rect 672349 169146 672415 169149
rect 672349 169144 676292 169146
rect 672349 169088 672354 169144
rect 672410 169088 676292 169144
rect 672349 169086 676292 169088
rect 672349 169083 672415 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 674005 168738 674071 168741
rect 674005 168736 676292 168738
rect 674005 168680 674010 168736
rect 674066 168680 676292 168736
rect 674005 168678 676292 168680
rect 674005 168675 674071 168678
rect 673729 168466 673795 168469
rect 667982 168464 673795 168466
rect 667982 168408 673734 168464
rect 673790 168408 673795 168464
rect 667982 168406 673795 168408
rect 667982 168330 668042 168406
rect 673729 168403 673795 168406
rect 666326 168270 668042 168330
rect 673870 168270 676292 168330
rect 666326 168028 666386 168270
rect 669773 168194 669839 168197
rect 673870 168194 673930 168270
rect 669773 168192 673930 168194
rect 669773 168136 669778 168192
rect 669834 168136 673930 168192
rect 669773 168134 673930 168136
rect 669773 168131 669839 168134
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675518 167452 675524 167516
rect 675588 167514 675594 167516
rect 675588 167454 676292 167514
rect 675588 167452 675594 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578969 166970 579035 166973
rect 575798 166968 579035 166970
rect 575798 166912 578974 166968
rect 579030 166912 579035 166968
rect 575798 166910 579035 166912
rect 575798 166532 575858 166910
rect 578969 166907 579035 166910
rect 671889 166970 671955 166973
rect 676170 166970 676230 167046
rect 671889 166968 676230 166970
rect 671889 166912 671894 166968
rect 671950 166912 676230 166968
rect 671889 166910 676230 166912
rect 671889 166907 671955 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 670325 165610 670391 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 670325 165608 676095 165610
rect 670325 165552 670330 165608
rect 670386 165552 676034 165608
rect 676090 165552 676095 165608
rect 670325 165550 676095 165552
rect 589457 165547 589523 165550
rect 670325 165547 670391 165550
rect 676029 165547 676095 165550
rect 667933 164794 667999 164797
rect 666356 164792 667999 164794
rect 666356 164736 667938 164792
rect 667994 164736 667999 164792
rect 666356 164734 667999 164736
rect 667933 164731 667999 164734
rect 578877 164522 578943 164525
rect 575798 164520 578943 164522
rect 575798 164464 578882 164520
rect 578938 164464 578943 164520
rect 575798 164462 578943 164464
rect 575798 164356 575858 164462
rect 578877 164459 578943 164462
rect 669129 164250 669195 164253
rect 673126 164250 673132 164252
rect 669129 164248 673132 164250
rect 669129 164192 669134 164248
rect 669190 164192 673132 164248
rect 669129 164190 673132 164192
rect 669129 164187 669195 164190
rect 673126 164188 673132 164190
rect 673196 164188 673202 164252
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668301 163162 668367 163165
rect 666356 163160 668367 163162
rect 666356 163104 668306 163160
rect 668362 163104 668367 163160
rect 666356 163102 668367 163104
rect 668301 163099 668367 163102
rect 579429 162482 579495 162485
rect 575798 162480 579495 162482
rect 575798 162424 579434 162480
rect 579490 162424 579495 162480
rect 575798 162422 579495 162424
rect 575798 162180 575858 162422
rect 579429 162419 579495 162422
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675334 161876 675340 161940
rect 675404 161938 675410 161940
rect 675937 161938 676003 161941
rect 675404 161936 676003 161938
rect 675404 161880 675942 161936
rect 675998 161880 676003 161936
rect 675404 161878 676003 161880
rect 675404 161876 675410 161878
rect 675937 161875 676003 161878
rect 676121 161394 676187 161397
rect 676078 161392 676187 161394
rect 676078 161336 676126 161392
rect 676182 161336 676187 161392
rect 676078 161331 676187 161336
rect 589457 160714 589523 160717
rect 675753 160714 675819 160717
rect 676078 160714 676138 161331
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 675753 160712 676138 160714
rect 675753 160656 675758 160712
rect 675814 160656 676138 160712
rect 675753 160654 676138 160656
rect 589457 160651 589523 160654
rect 675753 160651 675819 160654
rect 575982 159898 576042 160004
rect 579245 159898 579311 159901
rect 668945 159898 669011 159901
rect 575982 159896 579311 159898
rect 575982 159840 579250 159896
rect 579306 159840 579311 159896
rect 575982 159838 579311 159840
rect 666356 159896 669011 159898
rect 666356 159840 668950 159896
rect 669006 159840 669011 159896
rect 666356 159838 669011 159840
rect 579245 159835 579311 159838
rect 668945 159835 669011 159838
rect 675753 159354 675819 159357
rect 676438 159354 676444 159356
rect 675753 159352 676444 159354
rect 675753 159296 675758 159352
rect 675814 159296 676444 159352
rect 675753 159294 676444 159296
rect 675753 159291 675819 159294
rect 676438 159292 676444 159294
rect 676508 159292 676514 159356
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 579153 158266 579219 158269
rect 671705 158266 671771 158269
rect 575798 158264 579219 158266
rect 575798 158208 579158 158264
rect 579214 158208 579219 158264
rect 575798 158206 579219 158208
rect 666356 158264 671771 158266
rect 666356 158208 671710 158264
rect 671766 158208 671771 158264
rect 666356 158206 671771 158208
rect 575798 157828 575858 158206
rect 579153 158203 579219 158206
rect 671705 158203 671771 158206
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589457 157450 589523 157453
rect 589457 157448 592572 157450
rect 589457 157392 589462 157448
rect 589518 157392 592572 157448
rect 589457 157390 592572 157392
rect 589457 157387 589523 157390
rect 675385 157044 675451 157045
rect 675334 156980 675340 157044
rect 675404 157042 675451 157044
rect 675404 157040 675496 157042
rect 675446 156984 675496 157040
rect 675404 156982 675496 156984
rect 675404 156980 675451 156982
rect 675385 156979 675451 156980
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 579521 155954 579587 155957
rect 575798 155952 579587 155954
rect 575798 155896 579526 155952
rect 579582 155896 579587 155952
rect 575798 155894 579587 155896
rect 575798 155652 575858 155894
rect 579521 155891 579587 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 674373 155410 674439 155413
rect 675109 155410 675175 155413
rect 674373 155408 675175 155410
rect 674373 155352 674378 155408
rect 674434 155352 675114 155408
rect 675170 155352 675175 155408
rect 674373 155350 675175 155352
rect 674373 155347 674439 155350
rect 675109 155347 675175 155350
rect 666326 154594 666386 154972
rect 674230 154594 674236 154596
rect 666326 154534 674236 154594
rect 674230 154532 674236 154534
rect 674300 154532 674306 154596
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578233 154050 578299 154053
rect 575798 154048 578299 154050
rect 575798 153992 578238 154048
rect 578294 153992 578299 154048
rect 575798 153990 578299 153992
rect 575798 153476 575858 153990
rect 578233 153987 578299 153990
rect 668761 153370 668827 153373
rect 666356 153368 668827 153370
rect 666356 153312 668766 153368
rect 668822 153312 668827 153368
rect 666356 153310 668827 153312
rect 668761 153307 668827 153310
rect 672349 153098 672415 153101
rect 675109 153098 675175 153101
rect 672349 153096 675175 153098
rect 672349 153040 672354 153096
rect 672410 153040 675114 153096
rect 675170 153040 675175 153096
rect 672349 153038 675175 153040
rect 672349 153035 672415 153038
rect 675109 153035 675175 153038
rect 675753 153098 675819 153101
rect 676254 153098 676260 153100
rect 675753 153096 676260 153098
rect 675753 153040 675758 153096
rect 675814 153040 676260 153096
rect 675753 153038 676260 153040
rect 675753 153035 675819 153038
rect 676254 153036 676260 153038
rect 676324 153036 676330 153100
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 673177 151738 673243 151741
rect 675109 151738 675175 151741
rect 673177 151736 675175 151738
rect 673177 151680 673182 151736
rect 673238 151680 675114 151736
rect 675170 151680 675175 151736
rect 673177 151678 675175 151680
rect 673177 151675 673243 151678
rect 675109 151675 675175 151678
rect 674005 151058 674071 151061
rect 675109 151058 675175 151061
rect 674005 151056 675175 151058
rect 674005 151000 674010 151056
rect 674066 151000 675114 151056
rect 675170 151000 675175 151056
rect 674005 150998 675175 151000
rect 674005 150995 674071 150998
rect 675109 150995 675175 150998
rect 589457 150922 589523 150925
rect 589457 150920 592572 150922
rect 589457 150864 589462 150920
rect 589518 150864 592572 150920
rect 589457 150862 592572 150864
rect 589457 150859 589523 150862
rect 671521 150106 671587 150109
rect 666356 150104 671587 150106
rect 666356 150048 671526 150104
rect 671582 150048 671587 150104
rect 666356 150046 671587 150048
rect 671521 150043 671587 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589181 149290 589247 149293
rect 589181 149288 592572 149290
rect 589181 149232 589186 149288
rect 589242 149232 592572 149288
rect 589181 149230 592572 149232
rect 589181 149227 589247 149230
rect 668761 149154 668827 149157
rect 672717 149154 672783 149157
rect 668761 149152 672783 149154
rect 668761 149096 668766 149152
rect 668822 149096 672722 149152
rect 672778 149096 672783 149152
rect 668761 149094 672783 149096
rect 668761 149091 668827 149094
rect 672717 149091 672783 149094
rect 668485 148474 668551 148477
rect 666356 148472 668551 148474
rect 666356 148416 668490 148472
rect 668546 148416 668551 148472
rect 666356 148414 668551 148416
rect 668485 148411 668551 148414
rect 675661 148474 675727 148477
rect 675886 148474 675892 148476
rect 675661 148472 675892 148474
rect 675661 148416 675666 148472
rect 675722 148416 675892 148472
rect 675661 148414 675892 148416
rect 675661 148411 675727 148414
rect 675886 148412 675892 148414
rect 675956 148412 675962 148476
rect 589365 147658 589431 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 589365 147656 592572 147658
rect 589365 147600 589370 147656
rect 589426 147600 592572 147656
rect 589365 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 589365 147595 589431 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675661 147660 675727 147661
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 579521 147250 579587 147253
rect 575798 147248 579587 147250
rect 575798 147192 579526 147248
rect 579582 147192 579587 147248
rect 575798 147190 579587 147192
rect 575798 146948 575858 147190
rect 579521 147187 579587 147190
rect 589457 146026 589523 146029
rect 675753 146026 675819 146029
rect 676070 146026 676076 146028
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 675753 146024 676076 146026
rect 675753 145968 675758 146024
rect 675814 145968 676076 146024
rect 675753 145966 676076 145968
rect 589457 145963 589523 145966
rect 675753 145963 675819 145966
rect 676070 145964 676076 145966
rect 676140 145964 676146 146028
rect 668485 145210 668551 145213
rect 666356 145208 668551 145210
rect 666356 145152 668490 145208
rect 668546 145152 668551 145208
rect 666356 145150 668551 145152
rect 668485 145147 668551 145150
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589917 144394 589983 144397
rect 589917 144392 592572 144394
rect 589917 144336 589922 144392
rect 589978 144336 592572 144392
rect 589917 144334 592572 144336
rect 589917 144331 589983 144334
rect 669262 143578 669268 143580
rect 666356 143518 669268 143578
rect 669262 143516 669268 143518
rect 669332 143516 669338 143580
rect 578601 143034 578667 143037
rect 575798 143032 578667 143034
rect 575798 142976 578606 143032
rect 578662 142976 578667 143032
rect 575798 142974 578667 142976
rect 575798 142596 575858 142974
rect 578601 142971 578667 142974
rect 589457 142762 589523 142765
rect 589457 142760 592572 142762
rect 589457 142704 589462 142760
rect 589518 142704 592572 142760
rect 589457 142702 592572 142704
rect 589457 142699 589523 142702
rect 589089 141130 589155 141133
rect 589089 141128 592572 141130
rect 589089 141072 589094 141128
rect 589150 141072 592572 141128
rect 589089 141070 592572 141072
rect 589089 141067 589155 141070
rect 579521 140586 579587 140589
rect 575798 140584 579587 140586
rect 575798 140528 579526 140584
rect 579582 140528 579587 140584
rect 575798 140526 579587 140528
rect 575798 140420 575858 140526
rect 579521 140523 579587 140526
rect 672073 140314 672139 140317
rect 666356 140312 672139 140314
rect 666356 140256 672078 140312
rect 672134 140256 672139 140312
rect 666356 140254 672139 140256
rect 672073 140251 672139 140254
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578693 138818 578759 138821
rect 575798 138816 578759 138818
rect 575798 138760 578698 138816
rect 578754 138760 578759 138816
rect 575798 138758 578759 138760
rect 575798 138244 575858 138758
rect 578693 138755 578759 138758
rect 669129 138682 669195 138685
rect 666356 138680 669195 138682
rect 666356 138624 669134 138680
rect 669190 138624 669195 138680
rect 666356 138622 669195 138624
rect 669129 138619 669195 138622
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589273 136234 589339 136237
rect 589273 136232 592572 136234
rect 589273 136176 589278 136232
rect 589334 136176 592572 136232
rect 589273 136174 592572 136176
rect 589273 136171 589339 136174
rect 667565 135962 667631 135965
rect 683113 135962 683179 135965
rect 667565 135960 683179 135962
rect 667565 135904 667570 135960
rect 667626 135904 683118 135960
rect 683174 135904 683179 135960
rect 667565 135902 683179 135904
rect 667565 135899 667631 135902
rect 683113 135899 683179 135902
rect 668025 135418 668091 135421
rect 666356 135416 668091 135418
rect 666356 135360 668030 135416
rect 668086 135360 668091 135416
rect 666356 135358 668091 135360
rect 668025 135355 668091 135358
rect 589457 134602 589523 134605
rect 667197 134602 667263 134605
rect 675845 134602 675911 134605
rect 589457 134600 592572 134602
rect 589457 134544 589462 134600
rect 589518 134544 592572 134600
rect 589457 134542 592572 134544
rect 667197 134600 675911 134602
rect 667197 134544 667202 134600
rect 667258 134544 675850 134600
rect 675906 134544 675911 134600
rect 667197 134542 675911 134544
rect 589457 134539 589523 134542
rect 667197 134539 667263 134542
rect 675845 134539 675911 134542
rect 578325 134466 578391 134469
rect 575798 134464 578391 134466
rect 575798 134408 578330 134464
rect 578386 134408 578391 134464
rect 575798 134406 578391 134408
rect 575798 133892 575858 134406
rect 578325 134403 578391 134406
rect 670734 133786 670740 133788
rect 666356 133726 670740 133786
rect 670734 133724 670740 133726
rect 670804 133724 670810 133788
rect 667013 133106 667079 133109
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 667013 133104 676322 133106
rect 667013 133048 667018 133104
rect 667074 133048 676322 133104
rect 667013 133046 676322 133048
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 667013 133043 667079 133046
rect 676446 133043 676555 133048
rect 588537 132970 588603 132973
rect 588537 132968 592572 132970
rect 588537 132912 588542 132968
rect 588598 132912 592572 132968
rect 676446 132940 676506 133043
rect 588537 132910 592572 132912
rect 588537 132907 588603 132910
rect 683113 132698 683179 132701
rect 682886 132696 683179 132698
rect 682886 132640 683118 132696
rect 683174 132640 683179 132696
rect 682886 132638 683179 132640
rect 682886 132532 682946 132638
rect 683113 132635 683179 132638
rect 578233 132290 578299 132293
rect 575798 132288 578299 132290
rect 575798 132232 578238 132288
rect 578294 132232 578299 132288
rect 575798 132230 578299 132232
rect 575798 131716 575858 132230
rect 578233 132227 578299 132230
rect 674189 132154 674255 132157
rect 674189 132152 676292 132154
rect 674189 132096 674194 132152
rect 674250 132096 676292 132152
rect 674189 132094 676292 132096
rect 674189 132091 674255 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 590101 131338 590167 131341
rect 674649 131338 674715 131341
rect 590101 131336 592572 131338
rect 590101 131280 590106 131336
rect 590162 131280 592572 131336
rect 590101 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 590101 131275 590167 131278
rect 674649 131275 674715 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130522 667980 130524
rect 666356 130462 667980 130522
rect 667974 130460 667980 130462
rect 668044 130460 668050 130524
rect 672533 130522 672599 130525
rect 672533 130520 676292 130522
rect 672533 130464 672538 130520
rect 672594 130464 676292 130520
rect 672533 130462 676292 130464
rect 672533 130459 672599 130462
rect 675937 130114 676003 130117
rect 675937 130112 676292 130114
rect 675937 130056 675942 130112
rect 675998 130056 676292 130112
rect 675937 130054 676292 130056
rect 675937 130051 676003 130054
rect 579521 129706 579587 129709
rect 575798 129704 579587 129706
rect 575798 129648 579526 129704
rect 579582 129648 579587 129704
rect 575798 129646 579587 129648
rect 575798 129540 575858 129646
rect 579521 129643 579587 129646
rect 589457 129706 589523 129709
rect 673361 129706 673427 129709
rect 589457 129704 592572 129706
rect 589457 129648 589462 129704
rect 589518 129648 592572 129704
rect 589457 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 589457 129643 589523 129646
rect 673361 129643 673427 129646
rect 674097 129298 674163 129301
rect 674097 129296 676292 129298
rect 674097 129240 674102 129296
rect 674158 129240 676292 129296
rect 674097 129238 676292 129240
rect 674097 129235 674163 129238
rect 673494 128890 673500 128892
rect 666356 128830 673500 128890
rect 673494 128828 673500 128830
rect 673564 128828 673570 128892
rect 676630 128620 676690 128860
rect 676622 128556 676628 128620
rect 676692 128556 676698 128620
rect 668945 128346 669011 128349
rect 674046 128346 674052 128348
rect 668945 128344 674052 128346
rect 668945 128288 668950 128344
rect 669006 128288 674052 128344
rect 668945 128286 674052 128288
rect 668945 128283 669011 128286
rect 674046 128284 674052 128286
rect 674116 128284 674122 128348
rect 674281 128346 674347 128349
rect 675937 128346 676003 128349
rect 674281 128344 676003 128346
rect 674281 128288 674286 128344
rect 674342 128288 675942 128344
rect 675998 128288 676003 128344
rect 674281 128286 676003 128288
rect 674281 128283 674347 128286
rect 675937 128283 676003 128286
rect 676070 128148 676076 128212
rect 676140 128210 676146 128212
rect 676262 128210 676322 128452
rect 676140 128150 676322 128210
rect 676140 128148 676146 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 682334 127805 682394 128044
rect 578325 127802 578391 127805
rect 575798 127800 578391 127802
rect 575798 127744 578330 127800
rect 578386 127744 578391 127800
rect 575798 127742 578391 127744
rect 682334 127800 682443 127805
rect 682334 127744 682382 127800
rect 682438 127744 682443 127800
rect 682334 127742 682443 127744
rect 575798 127364 575858 127742
rect 578325 127739 578391 127742
rect 682377 127739 682443 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 676254 126924 676260 126988
rect 676324 126924 676330 126988
rect 676262 126820 676322 126924
rect 590285 126442 590351 126445
rect 675017 126442 675083 126445
rect 590285 126440 592572 126442
rect 590285 126384 590290 126440
rect 590346 126384 592572 126440
rect 590285 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 590285 126379 590351 126382
rect 675017 126379 675083 126382
rect 673269 126034 673335 126037
rect 673269 126032 676292 126034
rect 673269 125976 673274 126032
rect 673330 125976 676292 126032
rect 673269 125974 676292 125976
rect 673269 125971 673335 125974
rect 668761 125626 668827 125629
rect 666356 125624 668827 125626
rect 666356 125568 668766 125624
rect 668822 125568 668827 125624
rect 666356 125566 668827 125568
rect 668761 125563 668827 125566
rect 674649 125626 674715 125629
rect 674649 125624 676292 125626
rect 674649 125568 674654 125624
rect 674710 125568 676292 125624
rect 674649 125566 676292 125568
rect 674649 125563 674715 125566
rect 579245 125354 579311 125357
rect 575798 125352 579311 125354
rect 575798 125296 579250 125352
rect 579306 125296 579311 125352
rect 575798 125294 579311 125296
rect 575798 125188 575858 125294
rect 579245 125291 579311 125294
rect 674465 125218 674531 125221
rect 674465 125216 676292 125218
rect 674465 125160 674470 125216
rect 674526 125160 676292 125216
rect 674465 125158 676292 125160
rect 674465 125155 674531 125158
rect 589457 124810 589523 124813
rect 589457 124808 592572 124810
rect 589457 124752 589462 124808
rect 589518 124752 592572 124808
rect 589457 124750 592572 124752
rect 589457 124747 589523 124750
rect 676446 124540 676506 124780
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 672349 124402 672415 124405
rect 672349 124400 676292 124402
rect 672349 124344 672354 124400
rect 672410 124344 676292 124400
rect 672349 124342 676292 124344
rect 672349 124339 672415 124342
rect 672901 123994 672967 123997
rect 666356 123992 672967 123994
rect 666356 123936 672906 123992
rect 672962 123936 672967 123992
rect 666356 123934 672967 123936
rect 672901 123931 672967 123934
rect 673085 123994 673151 123997
rect 673085 123992 676292 123994
rect 673085 123936 673090 123992
rect 673146 123936 676292 123992
rect 673085 123934 676292 123936
rect 673085 123931 673151 123934
rect 579245 123586 579311 123589
rect 575798 123584 579311 123586
rect 575798 123528 579250 123584
rect 579306 123528 579311 123584
rect 575798 123526 579311 123528
rect 575798 123012 575858 123526
rect 579245 123523 579311 123526
rect 673361 123586 673427 123589
rect 673361 123584 676292 123586
rect 673361 123528 673366 123584
rect 673422 123528 676292 123584
rect 673361 123526 676292 123528
rect 673361 123523 673427 123526
rect 589457 123178 589523 123181
rect 672809 123178 672875 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672809 123176 676292 123178
rect 672809 123120 672814 123176
rect 672870 123120 676292 123176
rect 672809 123118 676292 123120
rect 589457 123115 589523 123118
rect 672809 123115 672875 123118
rect 669589 122770 669655 122773
rect 669589 122768 676292 122770
rect 669589 122712 669594 122768
rect 669650 122712 676292 122768
rect 669589 122710 676292 122712
rect 669589 122707 669655 122710
rect 675702 122300 675708 122364
rect 675772 122362 675778 122364
rect 675772 122302 676292 122362
rect 675772 122300 675778 122302
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589457 121546 589523 121549
rect 589457 121544 592572 121546
rect 589457 121488 589462 121544
rect 589518 121488 592572 121544
rect 589457 121486 592572 121488
rect 589457 121483 589523 121486
rect 669221 121410 669287 121413
rect 672809 121410 672875 121413
rect 669221 121408 672875 121410
rect 669221 121352 669226 121408
rect 669282 121352 672814 121408
rect 672870 121352 672875 121408
rect 669221 121350 672875 121352
rect 669221 121347 669287 121350
rect 672809 121347 672875 121350
rect 579061 121138 579127 121141
rect 575798 121136 579127 121138
rect 575798 121080 579066 121136
rect 579122 121080 579127 121136
rect 575798 121078 579127 121080
rect 575798 120836 575858 121078
rect 579061 121075 579127 121078
rect 672533 121138 672599 121141
rect 675894 121138 675954 121622
rect 672533 121136 675954 121138
rect 672533 121080 672538 121136
rect 672594 121080 675954 121136
rect 672533 121078 675954 121080
rect 672533 121075 672599 121078
rect 668945 120730 669011 120733
rect 666356 120728 669011 120730
rect 666356 120672 668950 120728
rect 669006 120672 669011 120728
rect 666356 120670 669011 120672
rect 668945 120667 669011 120670
rect 589917 119914 589983 119917
rect 589917 119912 592572 119914
rect 589917 119856 589922 119912
rect 589978 119856 592572 119912
rect 589917 119854 592572 119856
rect 589917 119851 589983 119854
rect 668209 119098 668275 119101
rect 666356 119096 668275 119098
rect 666356 119040 668214 119096
rect 668270 119040 668275 119096
rect 666356 119038 668275 119040
rect 668209 119035 668275 119038
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 588721 118282 588787 118285
rect 588721 118280 592572 118282
rect 588721 118224 588726 118280
rect 588782 118224 592572 118280
rect 588721 118222 592572 118224
rect 588721 118219 588787 118222
rect 668025 117466 668091 117469
rect 666356 117464 668091 117466
rect 666356 117408 668030 117464
rect 668086 117408 668091 117464
rect 666356 117406 668091 117408
rect 668025 117403 668091 117406
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 671889 115834 671955 115837
rect 666356 115832 671955 115834
rect 666356 115776 671894 115832
rect 671950 115776 671955 115832
rect 666356 115774 671955 115776
rect 671889 115771 671955 115774
rect 589641 115018 589707 115021
rect 589641 115016 592572 115018
rect 589641 114960 589646 115016
rect 589702 114960 592572 115016
rect 589641 114958 592572 114960
rect 589641 114955 589707 114958
rect 579521 114474 579587 114477
rect 575798 114472 579587 114474
rect 575798 114416 579526 114472
rect 579582 114416 579587 114472
rect 575798 114414 579587 114416
rect 575798 114308 575858 114414
rect 579521 114411 579587 114414
rect 669221 114202 669287 114205
rect 666356 114200 669287 114202
rect 666356 114144 669226 114200
rect 669282 114144 669287 114200
rect 666356 114142 669287 114144
rect 669221 114139 669287 114142
rect 589549 113386 589615 113389
rect 589549 113384 592572 113386
rect 589549 113328 589554 113384
rect 589610 113328 592572 113384
rect 589549 113326 592572 113328
rect 589549 113323 589615 113326
rect 675293 113114 675359 113117
rect 676622 113114 676628 113116
rect 675293 113112 676628 113114
rect 675293 113056 675298 113112
rect 675354 113056 676628 113112
rect 675293 113054 676628 113056
rect 675293 113051 675359 113054
rect 676622 113052 676628 113054
rect 676692 113052 676698 113116
rect 579521 112706 579587 112709
rect 575798 112704 579587 112706
rect 575798 112648 579526 112704
rect 579582 112648 579587 112704
rect 575798 112646 579587 112648
rect 575798 112132 575858 112646
rect 579521 112643 579587 112646
rect 668209 112570 668275 112573
rect 666356 112568 668275 112570
rect 666356 112512 668214 112568
rect 668270 112512 668275 112568
rect 666356 112510 668275 112512
rect 668209 112507 668275 112510
rect 668301 111890 668367 111893
rect 674097 111890 674163 111893
rect 668301 111888 674163 111890
rect 668301 111832 668306 111888
rect 668362 111832 674102 111888
rect 674158 111832 674163 111888
rect 668301 111830 674163 111832
rect 668301 111827 668367 111830
rect 674097 111827 674163 111830
rect 589457 111754 589523 111757
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 589457 111691 589523 111694
rect 673085 111482 673151 111485
rect 675109 111482 675175 111485
rect 673085 111480 675175 111482
rect 673085 111424 673090 111480
rect 673146 111424 675114 111480
rect 675170 111424 675175 111480
rect 673085 111422 675175 111424
rect 673085 111419 673151 111422
rect 675109 111419 675175 111422
rect 672533 110938 672599 110941
rect 666356 110936 672599 110938
rect 666356 110880 672538 110936
rect 672594 110880 672599 110936
rect 666356 110878 672599 110880
rect 672533 110875 672599 110878
rect 579429 110258 579495 110261
rect 575798 110256 579495 110258
rect 575798 110200 579434 110256
rect 579490 110200 579495 110256
rect 575798 110198 579495 110200
rect 575798 109956 575858 110198
rect 579429 110195 579495 110198
rect 672349 110258 672415 110261
rect 674649 110258 674715 110261
rect 672349 110256 674715 110258
rect 672349 110200 672354 110256
rect 672410 110200 674654 110256
rect 674710 110200 674715 110256
rect 672349 110198 674715 110200
rect 672349 110195 672415 110198
rect 674649 110195 674715 110198
rect 589273 110122 589339 110125
rect 589273 110120 592572 110122
rect 589273 110064 589278 110120
rect 589334 110064 592572 110120
rect 589273 110062 592572 110064
rect 589273 110059 589339 110062
rect 668025 109306 668091 109309
rect 666356 109304 668091 109306
rect 666356 109248 668030 109304
rect 668086 109248 668091 109304
rect 666356 109246 668091 109248
rect 668025 109243 668091 109246
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 671521 107674 671587 107677
rect 666356 107672 671587 107674
rect 666356 107616 671526 107672
rect 671582 107616 671587 107672
rect 666356 107614 671587 107616
rect 671521 107611 671587 107614
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 672809 106450 672875 106453
rect 675109 106450 675175 106453
rect 672809 106448 675175 106450
rect 672809 106392 672814 106448
rect 672870 106392 675114 106448
rect 675170 106392 675175 106448
rect 672809 106390 675175 106392
rect 672809 106387 672875 106390
rect 675109 106387 675175 106390
rect 675753 106178 675819 106181
rect 676438 106178 676444 106180
rect 675753 106176 676444 106178
rect 675753 106120 675758 106176
rect 675814 106120 676444 106176
rect 675753 106118 676444 106120
rect 675753 106115 675819 106118
rect 676438 106116 676444 106118
rect 676508 106116 676514 106180
rect 666645 106042 666711 106045
rect 667197 106042 667263 106045
rect 666356 106040 667263 106042
rect 666356 105984 666650 106040
rect 666706 105984 667202 106040
rect 667258 105984 667263 106040
rect 666356 105982 667263 105984
rect 666645 105979 666711 105982
rect 667197 105979 667263 105982
rect 578325 105906 578391 105909
rect 575798 105904 578391 105906
rect 575798 105848 578330 105904
rect 578386 105848 578391 105904
rect 575798 105846 578391 105848
rect 575798 105604 575858 105846
rect 578325 105843 578391 105846
rect 673361 105634 673427 105637
rect 675109 105634 675175 105637
rect 673361 105632 675175 105634
rect 673361 105576 673366 105632
rect 673422 105576 675114 105632
rect 675170 105576 675175 105632
rect 673361 105574 675175 105576
rect 673361 105571 673427 105574
rect 675109 105571 675175 105574
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 668301 104410 668367 104413
rect 666356 104408 668367 104410
rect 666356 104352 668306 104408
rect 668362 104352 668367 104408
rect 666356 104350 668367 104352
rect 668301 104347 668367 104350
rect 590101 103594 590167 103597
rect 590101 103592 592572 103594
rect 590101 103536 590106 103592
rect 590162 103536 592572 103592
rect 590101 103534 592572 103536
rect 590101 103531 590167 103534
rect 575982 103322 576042 103428
rect 579521 103322 579587 103325
rect 575982 103320 579587 103322
rect 575982 103264 579526 103320
rect 579582 103264 579587 103320
rect 575982 103262 579587 103264
rect 579521 103259 579587 103262
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 666326 102234 666386 102748
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 668485 102234 668551 102237
rect 674281 102234 674347 102237
rect 666326 102232 674347 102234
rect 666326 102176 668490 102232
rect 668546 102176 674286 102232
rect 674342 102176 674347 102232
rect 666326 102174 674347 102176
rect 668485 102171 668551 102174
rect 674281 102171 674347 102174
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579245 101826 579311 101829
rect 575798 101824 579311 101826
rect 575798 101768 579250 101824
rect 579306 101768 579311 101824
rect 575798 101766 579311 101768
rect 575798 101252 575858 101766
rect 579245 101763 579311 101766
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 579521 97474 579587 97477
rect 575798 97472 579587 97474
rect 575798 97416 579526 97472
rect 579582 97416 579587 97472
rect 575798 97414 579587 97416
rect 575798 96900 575858 97414
rect 579521 97411 579587 97414
rect 634854 96596 634860 96660
rect 634924 96658 634930 96660
rect 635733 96658 635799 96661
rect 634924 96656 635799 96658
rect 634924 96600 635738 96656
rect 635794 96600 635799 96656
rect 634924 96598 635799 96600
rect 634924 96596 634930 96598
rect 635733 96595 635799 96598
rect 637021 96658 637087 96661
rect 637246 96658 637252 96660
rect 637021 96656 637252 96658
rect 637021 96600 637026 96656
rect 637082 96600 637252 96656
rect 637021 96598 637252 96600
rect 637021 96595 637087 96598
rect 637246 96596 637252 96598
rect 637316 96596 637322 96660
rect 626441 95434 626507 95437
rect 626441 95432 628268 95434
rect 626441 95376 626446 95432
rect 626502 95376 628268 95432
rect 626441 95374 628268 95376
rect 626441 95371 626507 95374
rect 643185 95162 643251 95165
rect 642958 95160 643251 95162
rect 642958 95104 643190 95160
rect 643246 95104 643251 95160
rect 642958 95102 643251 95104
rect 579521 95026 579587 95029
rect 575798 95024 579587 95026
rect 575798 94968 579526 95024
rect 579582 94968 579587 95024
rect 575798 94966 579587 94968
rect 575798 94724 575858 94966
rect 579521 94963 579587 94966
rect 642958 94588 643018 95102
rect 643185 95099 643251 95102
rect 626257 94482 626323 94485
rect 626257 94480 628268 94482
rect 626257 94424 626262 94480
rect 626318 94424 628268 94480
rect 626257 94422 628268 94424
rect 626257 94419 626323 94422
rect 655237 94210 655303 94213
rect 655237 94208 656788 94210
rect 655237 94152 655242 94208
rect 655298 94152 656788 94208
rect 655237 94150 656788 94152
rect 655237 94147 655303 94150
rect 626441 93530 626507 93533
rect 626441 93528 628268 93530
rect 626441 93472 626446 93528
rect 626502 93472 628268 93528
rect 626441 93470 628268 93472
rect 626441 93467 626507 93470
rect 655053 93394 655119 93397
rect 665173 93394 665239 93397
rect 655053 93392 656788 93394
rect 655053 93336 655058 93392
rect 655114 93336 656788 93392
rect 655053 93334 656788 93336
rect 663596 93392 665239 93394
rect 663596 93336 665178 93392
rect 665234 93336 665239 93392
rect 663596 93334 665239 93336
rect 655053 93331 655119 93334
rect 665173 93331 665239 93334
rect 578509 93122 578575 93125
rect 663241 93122 663307 93125
rect 575798 93120 578575 93122
rect 575798 93064 578514 93120
rect 578570 93064 578575 93120
rect 575798 93062 578575 93064
rect 575798 92548 575858 93062
rect 578509 93059 578575 93062
rect 663198 93120 663307 93122
rect 663198 93064 663246 93120
rect 663302 93064 663307 93120
rect 663198 93059 663307 93064
rect 625613 92578 625679 92581
rect 654869 92578 654935 92581
rect 625613 92576 628268 92578
rect 625613 92520 625618 92576
rect 625674 92520 628268 92576
rect 625613 92518 628268 92520
rect 654869 92576 656788 92578
rect 654869 92520 654874 92576
rect 654930 92520 656788 92576
rect 663198 92548 663258 93059
rect 654869 92518 656788 92520
rect 625613 92515 625679 92518
rect 654869 92515 654935 92518
rect 644933 92170 644999 92173
rect 642988 92168 644999 92170
rect 642988 92112 644938 92168
rect 644994 92112 644999 92168
rect 642988 92110 644999 92112
rect 644933 92107 644999 92110
rect 663701 92034 663767 92037
rect 663382 92032 663767 92034
rect 663382 91976 663706 92032
rect 663762 91976 663767 92032
rect 663382 91974 663767 91976
rect 663382 91732 663442 91974
rect 663701 91971 663767 91974
rect 625429 91626 625495 91629
rect 625429 91624 628268 91626
rect 625429 91568 625434 91624
rect 625490 91568 628268 91624
rect 625429 91566 628268 91568
rect 625429 91563 625495 91566
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 579061 90946 579127 90949
rect 575798 90944 579127 90946
rect 575798 90888 579066 90944
rect 579122 90888 579127 90944
rect 575798 90886 579127 90888
rect 575798 90372 575858 90886
rect 579061 90883 579127 90886
rect 626441 90674 626507 90677
rect 654133 90674 654199 90677
rect 665357 90674 665423 90677
rect 626441 90672 628268 90674
rect 626441 90616 626446 90672
rect 626502 90616 628268 90672
rect 626441 90614 628268 90616
rect 654133 90672 656788 90674
rect 654133 90616 654138 90672
rect 654194 90616 656788 90672
rect 654133 90614 656788 90616
rect 663596 90672 665423 90674
rect 663596 90616 665362 90672
rect 665418 90616 665423 90672
rect 663596 90614 665423 90616
rect 626441 90611 626507 90614
rect 654133 90611 654199 90614
rect 665357 90611 665423 90614
rect 655789 89858 655855 89861
rect 664621 89858 664687 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664687 89858
rect 663596 89800 664626 89856
rect 664682 89800 664687 89856
rect 663596 89798 664687 89800
rect 655789 89795 655855 89798
rect 664621 89795 664687 89798
rect 625245 89722 625311 89725
rect 643369 89722 643435 89725
rect 625245 89720 628268 89722
rect 625245 89664 625250 89720
rect 625306 89664 628268 89720
rect 625245 89662 628268 89664
rect 642988 89720 643435 89722
rect 642988 89664 643374 89720
rect 643430 89664 643435 89720
rect 642988 89662 643435 89664
rect 625245 89659 625311 89662
rect 643369 89659 643435 89662
rect 664161 89042 664227 89045
rect 663596 89040 664227 89042
rect 663596 88984 664166 89040
rect 664222 88984 664227 89040
rect 663596 88982 664227 88984
rect 664161 88979 664227 88982
rect 626441 88906 626507 88909
rect 626441 88904 628268 88906
rect 626441 88848 626446 88904
rect 626502 88848 628268 88904
rect 626441 88846 628268 88848
rect 626441 88843 626507 88846
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643553 87138 643619 87141
rect 642988 87136 643619 87138
rect 642988 87080 643558 87136
rect 643614 87080 643619 87136
rect 642988 87078 643619 87080
rect 643553 87075 643619 87078
rect 625613 87002 625679 87005
rect 625613 87000 628268 87002
rect 625613 86944 625618 87000
rect 625674 86944 628268 87000
rect 625613 86942 628268 86944
rect 625613 86939 625679 86942
rect 578509 86458 578575 86461
rect 575798 86456 578575 86458
rect 575798 86400 578514 86456
rect 578570 86400 578575 86456
rect 575798 86398 578575 86400
rect 575798 86020 575858 86398
rect 578509 86395 578575 86398
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 644749 84690 644815 84693
rect 642988 84688 644815 84690
rect 642988 84632 644754 84688
rect 644810 84632 644815 84688
rect 642988 84630 644815 84632
rect 644749 84627 644815 84630
rect 625613 84146 625679 84149
rect 625613 84144 628268 84146
rect 625613 84088 625618 84144
rect 625674 84088 628268 84144
rect 625613 84086 628268 84088
rect 625613 84083 625679 84086
rect 579337 84010 579403 84013
rect 575798 84008 579403 84010
rect 575798 83952 579342 84008
rect 579398 83952 579403 84008
rect 575798 83950 579403 83952
rect 575798 83844 575858 83950
rect 579337 83947 579403 83950
rect 624417 82922 624483 82925
rect 628238 82922 628298 83164
rect 624417 82920 628298 82922
rect 624417 82864 624422 82920
rect 624478 82864 628298 82920
rect 624417 82862 628298 82864
rect 624417 82859 624483 82862
rect 643737 82786 643803 82789
rect 642958 82784 643803 82786
rect 642958 82728 643742 82784
rect 643798 82728 643803 82784
rect 642958 82726 643803 82728
rect 579245 82242 579311 82245
rect 575798 82240 579311 82242
rect 575798 82184 579250 82240
rect 579306 82184 579311 82240
rect 642958 82212 643018 82726
rect 643737 82723 643803 82726
rect 575798 82182 579311 82184
rect 575798 81668 575858 82182
rect 579245 82179 579311 82182
rect 628606 81701 628666 82212
rect 628606 81696 628715 81701
rect 628606 81640 628654 81696
rect 628710 81640 628715 81696
rect 628606 81638 628715 81640
rect 628649 81635 628715 81638
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 629201 80819 629267 80822
rect 633893 80474 633959 80477
rect 634854 80474 634860 80476
rect 633893 80472 634860 80474
rect 633893 80416 633898 80472
rect 633954 80416 634860 80472
rect 633893 80414 634860 80416
rect 633893 80411 633959 80414
rect 634854 80412 634860 80414
rect 634924 80412 634930 80476
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 579061 77890 579127 77893
rect 575798 77888 579127 77890
rect 575798 77832 579066 77888
rect 579122 77832 579127 77888
rect 575798 77830 579127 77832
rect 575798 77316 575858 77830
rect 579061 77827 579127 77830
rect 585777 77890 585843 77893
rect 637062 77890 637068 77892
rect 585777 77888 637068 77890
rect 585777 77832 585782 77888
rect 585838 77832 637068 77888
rect 585777 77830 637068 77832
rect 585777 77827 585843 77830
rect 637062 77828 637068 77830
rect 637132 77890 637138 77892
rect 639597 77890 639663 77893
rect 637132 77888 639663 77890
rect 637132 77832 639602 77888
rect 639658 77832 639663 77888
rect 637132 77830 639663 77832
rect 637132 77828 637138 77830
rect 639597 77827 639663 77830
rect 579245 75578 579311 75581
rect 575798 75576 579311 75578
rect 575798 75520 579250 75576
rect 579306 75520 579311 75576
rect 575798 75518 579311 75520
rect 575798 75140 575858 75518
rect 579245 75515 579311 75518
rect 647049 74490 647115 74493
rect 646668 74488 647115 74490
rect 646668 74432 647054 74488
rect 647110 74432 647115 74488
rect 646668 74430 647115 74432
rect 647049 74427 647115 74430
rect 578601 73130 578667 73133
rect 575798 73128 578667 73130
rect 575798 73072 578606 73128
rect 578662 73072 578667 73128
rect 575798 73070 578667 73072
rect 575798 72964 575858 73070
rect 578601 73067 578667 73070
rect 646865 72994 646931 72997
rect 646668 72992 646931 72994
rect 646668 72936 646870 72992
rect 646926 72936 646931 72992
rect 646668 72934 646931 72936
rect 646865 72931 646931 72934
rect 648981 71498 649047 71501
rect 646668 71496 649047 71498
rect 646668 71440 648986 71496
rect 649042 71440 649047 71496
rect 646668 71438 649047 71440
rect 648981 71435 649047 71438
rect 579061 71362 579127 71365
rect 575798 71360 579127 71362
rect 575798 71304 579066 71360
rect 579122 71304 579127 71360
rect 575798 71302 579127 71304
rect 575798 70788 575858 71302
rect 579061 71299 579127 71302
rect 647325 70002 647391 70005
rect 646668 70000 647391 70002
rect 646668 69944 647330 70000
rect 647386 69944 647391 70000
rect 646668 69942 647391 69944
rect 647325 69939 647391 69942
rect 646221 68914 646287 68917
rect 646221 68912 646330 68914
rect 646221 68856 646226 68912
rect 646282 68856 646330 68912
rect 646221 68851 646330 68856
rect 575982 68098 576042 68612
rect 646270 68476 646330 68851
rect 579521 68098 579587 68101
rect 575982 68096 579587 68098
rect 575982 68040 579526 68096
rect 579582 68040 579587 68096
rect 575982 68038 579587 68040
rect 579521 68035 579587 68038
rect 649165 67010 649231 67013
rect 646668 67008 649231 67010
rect 646668 66952 649170 67008
rect 649226 66952 649231 67008
rect 646668 66950 649231 66952
rect 649165 66947 649231 66950
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 647509 65514 647575 65517
rect 646668 65512 647575 65514
rect 646668 65456 647514 65512
rect 647570 65456 647575 65512
rect 646668 65454 647575 65456
rect 647509 65451 647575 65454
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 646086 63988 646146 64363
rect 575982 61842 576042 62084
rect 578509 61842 578575 61845
rect 575982 61840 578575 61842
rect 575982 61784 578514 61840
rect 578570 61784 578575 61840
rect 575982 61782 578575 61784
rect 578509 61779 578575 61782
rect 579521 60346 579587 60349
rect 575798 60344 579587 60346
rect 575798 60288 579526 60344
rect 579582 60288 579587 60344
rect 575798 60286 579587 60288
rect 575798 59908 575858 60286
rect 579521 60283 579587 60286
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 579521 56130 579587 56133
rect 575798 56128 579587 56130
rect 575798 56072 579526 56128
rect 579582 56072 579587 56128
rect 575798 56070 579587 56072
rect 575798 55556 575858 56070
rect 579521 56067 579587 56070
rect 461710 54980 461716 55044
rect 461780 55042 461786 55044
rect 581637 55042 581703 55045
rect 461780 55040 581703 55042
rect 461780 54984 581642 55040
rect 581698 54984 581703 55040
rect 461780 54982 581703 54984
rect 461780 54980 461786 54982
rect 581637 54979 581703 54982
rect 584397 54770 584463 54773
rect 459878 54768 584463 54770
rect 459878 54712 584402 54768
rect 584458 54712 584463 54768
rect 459878 54710 584463 54712
rect 459878 53685 459938 54710
rect 584397 54707 584463 54710
rect 462630 54436 462636 54500
rect 462700 54498 462706 54500
rect 604453 54498 604519 54501
rect 462700 54496 604519 54498
rect 462700 54440 604458 54496
rect 604514 54440 604519 54496
rect 462700 54438 604519 54440
rect 462700 54436 462706 54438
rect 604453 54435 604519 54438
rect 580257 54226 580323 54229
rect 460798 54224 580323 54226
rect 460798 54168 580262 54224
rect 580318 54168 580323 54224
rect 460798 54166 580323 54168
rect 460798 53685 460858 54166
rect 580257 54163 580323 54166
rect 461710 53892 461716 53956
rect 461780 53892 461786 53956
rect 462630 53892 462636 53956
rect 462700 53892 462706 53956
rect 461718 53685 461778 53892
rect 462638 53685 462698 53892
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462589 53680 462698 53685
rect 462589 53624 462594 53680
rect 462650 53624 462698 53680
rect 462589 53622 462698 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53619 462655 53622
rect 461899 52866 461965 52869
rect 465717 52866 465783 52869
rect 461899 52864 465783 52866
rect 461899 52808 461904 52864
rect 461960 52808 465722 52864
rect 465778 52808 465783 52864
rect 461899 52806 465783 52808
rect 461899 52803 461965 52806
rect 465717 52803 465783 52806
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 553669 50282 553735 50285
rect 529860 50280 553735 50282
rect 529860 50224 553674 50280
rect 553730 50224 553735 50280
rect 529860 50222 553735 50224
rect 529860 50220 529866 50222
rect 553669 50219 553735 50222
rect 308990 49676 308996 49740
rect 309060 49738 309066 49740
rect 309685 49738 309751 49741
rect 309060 49736 309751 49738
rect 309060 49680 309690 49736
rect 309746 49680 309751 49736
rect 309060 49678 309751 49680
rect 309060 49676 309066 49678
rect 309685 49675 309751 49678
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 663977 48514 664043 48517
rect 662094 48512 664043 48514
rect 661480 48456 663982 48512
rect 664038 48456 664043 48512
rect 661480 48454 664043 48456
rect 661480 48452 662154 48454
rect 663977 48451 664043 48454
rect 526478 48044 526484 48108
rect 526548 48106 526554 48108
rect 552013 48106 552079 48109
rect 526548 48104 552079 48106
rect 526548 48048 552018 48104
rect 552074 48048 552079 48104
rect 526548 48046 552079 48048
rect 526548 48044 526554 48046
rect 552013 48043 552079 48046
rect 520958 47772 520964 47836
rect 521028 47834 521034 47836
rect 547873 47834 547939 47837
rect 663793 47834 663859 47837
rect 521028 47832 547939 47834
rect 521028 47776 547878 47832
rect 547934 47776 547939 47832
rect 661910 47832 663859 47834
rect 661910 47791 663798 47832
rect 521028 47774 547939 47776
rect 521028 47772 521034 47774
rect 547873 47771 547939 47774
rect 661388 47776 663798 47791
rect 663854 47776 663859 47832
rect 661388 47774 663859 47776
rect 661388 47731 661970 47774
rect 663793 47771 663859 47774
rect 515438 47500 515444 47564
rect 515508 47562 515514 47564
rect 544009 47562 544075 47565
rect 515508 47560 544075 47562
rect 515508 47504 544014 47560
rect 544070 47504 544075 47560
rect 515508 47502 544075 47504
rect 515508 47500 515514 47502
rect 544009 47499 544075 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 461342 44372 461348 44436
rect 461412 44434 461418 44436
rect 461945 44434 462011 44437
rect 461412 44432 462011 44434
rect 461412 44376 461950 44432
rect 462006 44376 462011 44432
rect 461412 44374 462011 44376
rect 461412 44372 461418 44374
rect 461945 44371 462011 44374
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462497 44434 462563 44437
rect 462332 44432 462563 44434
rect 462332 44376 462502 44432
rect 462558 44376 462563 44432
rect 462332 44374 462563 44376
rect 462332 44372 462338 44374
rect 462497 44371 462563 44374
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 310421 44162 310487 44165
rect 364885 44162 364951 44165
rect 463693 44162 463759 44165
rect 310421 44160 354690 44162
rect 310421 44104 310426 44160
rect 310482 44104 354690 44160
rect 310421 44102 354690 44104
rect 310421 44099 310487 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 354630 43890 354690 44102
rect 364885 44160 463759 44162
rect 364885 44104 364890 44160
rect 364946 44104 463698 44160
rect 463754 44104 463759 44160
rect 364885 44102 463759 44104
rect 364885 44099 364951 44102
rect 463693 44099 463759 44102
rect 440182 43890 440188 43892
rect 354630 43830 440188 43890
rect 440182 43828 440188 43830
rect 440252 43828 440258 43892
rect 440918 43828 440924 43892
rect 440988 43890 440994 43892
rect 462957 43890 463023 43893
rect 440988 43888 463023 43890
rect 440988 43832 462962 43888
rect 463018 43832 463023 43888
rect 440988 43830 463023 43832
rect 440988 43828 440994 43830
rect 462957 43827 463023 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463693 42938 463759 42941
rect 461761 42936 463759 42938
rect 461761 42880 461766 42936
rect 461822 42880 463698 42936
rect 463754 42880 463759 42936
rect 461761 42878 463759 42880
rect 461761 42875 461827 42878
rect 463693 42875 463759 42878
rect 308949 42804 309015 42805
rect 518801 42804 518867 42805
rect 308949 42800 308996 42804
rect 309060 42802 309066 42804
rect 518750 42802 518756 42804
rect 308949 42744 308954 42800
rect 308949 42740 308996 42744
rect 309060 42742 309106 42802
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 309060 42740 309066 42742
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 308949 42739 309015 42740
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 443545 42258 443611 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 443545 42256 461183 42258
rect 443545 42200 443550 42256
rect 443606 42200 461122 42256
rect 461178 42200 461183 42256
rect 443545 42198 461183 42200
rect 443545 42195 443611 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 443545 41578 443611 41581
rect 427770 41576 443611 41578
rect 427770 41520 443550 41576
rect 443606 41520 443611 41576
rect 427770 41518 443611 41520
rect 443545 41515 443611 41518
rect 141693 40492 141759 40493
rect 141693 40488 141740 40492
rect 141804 40490 141810 40492
rect 141693 40432 141698 40488
rect 141693 40428 141740 40432
rect 141804 40430 141850 40490
rect 141804 40428 141810 40430
rect 141693 40427 141759 40428
<< via3 >>
rect 89484 997188 89548 997252
rect 195284 997188 195348 997252
rect 189764 997052 189828 997116
rect 243492 997188 243556 997252
rect 243860 996916 243924 996980
rect 89852 996236 89916 996300
rect 140084 996236 140148 996300
rect 89300 995556 89364 995620
rect 89484 995616 89548 995620
rect 89484 995560 89534 995616
rect 89534 995560 89548 995616
rect 89484 995556 89548 995560
rect 132356 995964 132420 996028
rect 132540 995692 132604 995756
rect 188108 996372 188172 996436
rect 194916 996644 194980 996708
rect 192340 996372 192404 996436
rect 191604 995964 191668 996028
rect 188108 995752 188172 995756
rect 188108 995696 188122 995752
rect 188122 995696 188172 995752
rect 188108 995692 188172 995696
rect 189764 995692 189828 995756
rect 192340 995616 192404 995620
rect 192340 995560 192354 995616
rect 192354 995560 192404 995616
rect 192340 995556 192404 995560
rect 287836 997188 287900 997252
rect 524092 997732 524156 997796
rect 385908 997188 385972 997252
rect 511028 997248 511092 997252
rect 511028 997192 511042 997248
rect 511042 997192 511092 997248
rect 511028 997188 511092 997192
rect 532556 997188 532620 997252
rect 553532 997188 553596 997252
rect 630260 997188 630324 997252
rect 295380 996916 295444 996980
rect 633940 996916 634004 996980
rect 291516 996644 291580 996708
rect 388668 996644 388732 996708
rect 529796 996644 529860 996708
rect 396580 996372 396644 996436
rect 385356 996236 385420 996300
rect 243492 995752 243556 995756
rect 243492 995696 243506 995752
rect 243506 995696 243556 995752
rect 243492 995692 243556 995696
rect 243860 995752 243924 995756
rect 243860 995696 243874 995752
rect 243874 995696 243924 995752
rect 243860 995692 243924 995696
rect 292252 996100 292316 996164
rect 484348 996236 484412 996300
rect 295380 995752 295444 995756
rect 295380 995696 295394 995752
rect 295394 995696 295444 995752
rect 295380 995692 295444 995696
rect 132356 995344 132420 995348
rect 132356 995288 132406 995344
rect 132406 995288 132420 995344
rect 132356 995284 132420 995288
rect 140820 995284 140884 995348
rect 292436 995556 292500 995620
rect 364196 995828 364260 995892
rect 388484 995692 388548 995756
rect 388668 995752 388732 995756
rect 388668 995696 388718 995752
rect 388718 995696 388732 995752
rect 388668 995692 388732 995696
rect 484348 995692 484412 995756
rect 393452 995420 393516 995484
rect 396580 995480 396644 995484
rect 396580 995424 396594 995480
rect 396594 995424 396644 995480
rect 396580 995420 396644 995424
rect 385356 995038 385420 995042
rect 385356 994982 385406 995038
rect 385406 994982 385420 995038
rect 388484 995012 388548 995076
rect 532004 995692 532068 995756
rect 532556 995692 532620 995756
rect 538260 996644 538324 996708
rect 627868 996644 627932 996708
rect 529796 995616 529860 995620
rect 529796 995560 529846 995616
rect 529846 995560 529860 995616
rect 529796 995556 529860 995560
rect 522804 995012 522868 995076
rect 627868 995752 627932 995756
rect 627868 995696 627918 995752
rect 627918 995696 627932 995752
rect 627868 995692 627932 995696
rect 630260 995752 630324 995756
rect 630260 995696 630310 995752
rect 630310 995696 630324 995752
rect 630260 995692 630324 995696
rect 633940 995752 634004 995756
rect 633940 995696 633990 995752
rect 633990 995696 634004 995752
rect 633940 995692 634004 995696
rect 636700 995692 636764 995756
rect 385356 994978 385420 994982
rect 385908 994936 385972 994940
rect 385908 994880 385958 994936
rect 385958 994880 385972 994936
rect 385908 994876 385972 994880
rect 191604 994740 191668 994804
rect 287836 994800 287900 994804
rect 287836 994744 287850 994800
rect 287850 994744 287900 994800
rect 287836 994740 287900 994744
rect 291516 994800 291580 994804
rect 291516 994744 291530 994800
rect 291530 994744 291580 994800
rect 291516 994740 291580 994744
rect 538260 994468 538324 994532
rect 132540 993788 132604 993852
rect 141924 993380 141988 993444
rect 142292 993380 142356 993444
rect 41460 967132 41524 967196
rect 676076 965092 676140 965156
rect 676628 963596 676692 963660
rect 675340 963384 675404 963388
rect 675340 963328 675390 963384
rect 675390 963328 675404 963384
rect 675340 963324 675404 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 41276 959788 41340 959852
rect 675156 959304 675220 959308
rect 675156 959248 675206 959304
rect 675206 959248 675220 959304
rect 675156 959244 675220 959248
rect 40540 959108 40604 959172
rect 41828 957808 41892 957812
rect 41828 957752 41842 957808
rect 41842 957752 41892 957808
rect 41828 957748 41892 957752
rect 676812 957748 676876 957812
rect 676996 956388 677060 956452
rect 40724 955436 40788 955500
rect 675340 954484 675404 954548
rect 41828 952852 41892 952916
rect 41460 952444 41524 952508
rect 41644 952172 41708 952236
rect 41276 951628 41340 951692
rect 676628 951492 676692 951556
rect 675156 951144 675220 951148
rect 675156 951088 675206 951144
rect 675206 951088 675220 951144
rect 675156 951084 675220 951088
rect 676076 950676 676140 950740
rect 40356 944012 40420 944076
rect 42196 944012 42260 944076
rect 40724 943740 40788 943804
rect 42012 943740 42076 943804
rect 41828 939388 41892 939452
rect 41828 936532 41892 936596
rect 41828 935716 41892 935780
rect 676996 931908 677060 931972
rect 676812 931500 676876 931564
rect 42012 911916 42076 911980
rect 42196 911644 42260 911708
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 676076 875876 676140 875940
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 673868 873156 673932 873220
rect 676812 870844 676876 870908
rect 675340 863152 675404 863156
rect 675340 863096 675354 863152
rect 675354 863096 675404 863152
rect 675340 863092 675404 863096
rect 39988 814234 40052 814298
rect 41828 813180 41892 813244
rect 42196 808692 42260 808756
rect 42012 805564 42076 805628
rect 40724 805488 40788 805492
rect 40724 805432 40774 805488
rect 40774 805432 40788 805488
rect 40724 805428 40788 805432
rect 41644 805292 41708 805356
rect 40908 805020 40972 805084
rect 40540 804748 40604 804812
rect 42196 804748 42260 804812
rect 40908 795364 40972 795428
rect 40724 794140 40788 794204
rect 40540 792508 40604 792572
rect 41644 788972 41708 789036
rect 41828 788624 41892 788628
rect 41828 788568 41842 788624
rect 41842 788568 41892 788624
rect 41828 788564 41892 788568
rect 41460 786796 41524 786860
rect 675524 777004 675588 777068
rect 675524 775704 675588 775708
rect 675524 775648 675574 775704
rect 675574 775648 675588 775704
rect 675524 775644 675588 775648
rect 675708 775568 675772 775572
rect 675708 775512 675758 775568
rect 675758 775512 675772 775568
rect 675708 775508 675772 775512
rect 676996 774420 677060 774484
rect 675708 774284 675772 774348
rect 676076 772652 676140 772716
rect 673868 770884 673932 770948
rect 41460 769796 41524 769860
rect 675156 768164 675220 768228
rect 676076 766532 676140 766596
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 40724 764900 40788 764964
rect 41644 764492 41708 764556
rect 676996 761968 677060 761972
rect 676996 761912 677046 761968
rect 677046 761912 677060 761968
rect 676996 761908 677060 761912
rect 676812 761832 676876 761836
rect 676812 761776 676826 761832
rect 676826 761776 676876 761832
rect 676812 761772 676876 761776
rect 41828 757692 41892 757756
rect 42012 756332 42076 756396
rect 40908 754836 40972 754900
rect 42012 754080 42076 754084
rect 42012 754024 42026 754080
rect 42026 754024 42076 754080
rect 42012 754020 42076 754024
rect 42196 753204 42260 753268
rect 42196 751768 42260 751772
rect 42196 751712 42210 751768
rect 42210 751712 42260 751768
rect 42196 751708 42260 751712
rect 40724 750348 40788 750412
rect 40540 747356 40604 747420
rect 41644 745044 41708 745108
rect 41828 744772 41892 744836
rect 41460 743684 41524 743748
rect 674420 742460 674484 742524
rect 674236 741508 674300 741572
rect 674604 739604 674668 739668
rect 672028 732864 672092 732868
rect 672028 732808 672042 732864
rect 672042 732808 672092 732864
rect 672028 732804 672092 732808
rect 673316 732864 673380 732868
rect 673316 732808 673366 732864
rect 673366 732808 673380 732864
rect 673316 732804 673380 732808
rect 675892 729948 675956 730012
rect 676812 729948 676876 730012
rect 673316 728512 673380 728516
rect 673316 728456 673366 728512
rect 673366 728456 673380 728512
rect 673316 728452 673380 728456
rect 672028 728180 672092 728244
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 41828 722332 41892 722396
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 718524 40604 718588
rect 41828 718524 41892 718588
rect 42012 714716 42076 714780
rect 41828 714444 41892 714508
rect 41276 714232 41340 714236
rect 41276 714176 41326 714232
rect 41326 714176 41340 714232
rect 41276 714172 41340 714176
rect 42380 713220 42444 713284
rect 41276 712132 41340 712196
rect 675892 711996 675956 712060
rect 41828 709880 41892 709884
rect 41828 709824 41878 709880
rect 41878 709824 41892 709880
rect 41828 709820 41892 709824
rect 40724 707372 40788 707436
rect 42380 707372 42444 707436
rect 40540 706420 40604 706484
rect 41644 702340 41708 702404
rect 41460 700436 41524 700500
rect 42196 699952 42260 699956
rect 42196 699896 42210 699952
rect 42210 699896 42260 699952
rect 42196 699892 42260 699896
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676996 694044 677060 694108
rect 675340 686428 675404 686492
rect 41828 683572 41892 683636
rect 674420 682620 674484 682684
rect 674236 682348 674300 682412
rect 41828 681048 41892 681052
rect 41828 680992 41842 681048
rect 41842 680992 41892 681048
rect 41828 680988 41892 680992
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 42564 673100 42628 673164
rect 42380 672828 42444 672892
rect 41828 671196 41892 671260
rect 674604 670108 674668 670172
rect 42196 669292 42260 669356
rect 674972 669292 675036 669356
rect 42564 668476 42628 668540
rect 40724 668204 40788 668268
rect 42012 667720 42076 667724
rect 42012 667664 42026 667720
rect 42026 667664 42076 667720
rect 42012 667660 42076 667664
rect 42380 666572 42444 666636
rect 40540 663988 40604 664052
rect 674420 663988 674484 664052
rect 41460 659636 41524 659700
rect 41644 658548 41708 658612
rect 41828 658276 41892 658340
rect 44220 653108 44284 653172
rect 675340 652836 675404 652900
rect 674972 651476 675036 651540
rect 675156 649768 675220 649772
rect 675156 649712 675206 649768
rect 675206 649712 675220 649768
rect 675156 649708 675220 649712
rect 674420 648892 674484 648956
rect 674420 647592 674484 647596
rect 674420 647536 674470 647592
rect 674470 647536 674484 647592
rect 674420 647532 674484 647536
rect 675156 647532 675220 647596
rect 674972 647320 675036 647324
rect 674972 647264 675022 647320
rect 675022 647264 675036 647320
rect 674972 647260 675036 647264
rect 674052 645084 674116 645148
rect 676812 644268 676876 644332
rect 675156 644056 675220 644060
rect 675156 644000 675206 644056
rect 675206 644000 675220 644056
rect 675156 643996 675220 644000
rect 671476 643452 671540 643516
rect 41644 640596 41708 640660
rect 676628 640188 676692 640252
rect 41460 639372 41524 639436
rect 675156 638012 675220 638076
rect 676628 637876 676692 637940
rect 675340 637604 675404 637668
rect 41828 637332 41892 637396
rect 40724 634884 40788 634948
rect 40540 634476 40604 634540
rect 675340 631348 675404 631412
rect 676076 631348 676140 631412
rect 42564 626588 42628 626652
rect 42196 625228 42260 625292
rect 42564 625016 42628 625020
rect 42564 624960 42578 625016
rect 42578 624960 42628 625016
rect 42564 624956 42628 624960
rect 42196 623324 42260 623388
rect 40724 622100 40788 622164
rect 40540 619788 40604 619852
rect 676996 619108 677060 619172
rect 673868 616116 673932 616180
rect 42012 615904 42076 615908
rect 42012 615848 42062 615904
rect 42062 615848 42076 615904
rect 42012 615844 42076 615848
rect 41460 615436 41524 615500
rect 41828 614136 41892 614140
rect 41828 614080 41878 614136
rect 41878 614080 41892 614136
rect 41828 614076 41892 614080
rect 44220 614076 44284 614140
rect 675524 607744 675588 607748
rect 675524 607688 675538 607744
rect 675538 607688 675588 607744
rect 675524 607684 675588 607688
rect 674420 602924 674484 602988
rect 42012 597212 42076 597276
rect 41828 596396 41892 596460
rect 676076 593404 676140 593468
rect 676996 593404 677060 593468
rect 41828 593132 41892 593196
rect 42196 592316 42260 592380
rect 675340 592316 675404 592380
rect 675524 592104 675588 592108
rect 675524 592048 675574 592104
rect 675574 592048 675588 592104
rect 675524 592044 675588 592048
rect 43852 591500 43916 591564
rect 40540 589656 40604 589660
rect 40540 589600 40554 589656
rect 40554 589600 40604 589656
rect 40540 589596 40604 589600
rect 40724 589596 40788 589660
rect 41828 589596 41892 589660
rect 40908 589324 40972 589388
rect 42196 589324 42260 589388
rect 676076 586196 676140 586260
rect 42012 585380 42076 585444
rect 41828 585108 41892 585172
rect 41092 584564 41156 584628
rect 42012 580484 42076 580548
rect 41092 580212 41156 580276
rect 40724 578172 40788 578236
rect 40908 577492 40972 577556
rect 42380 577416 42444 577420
rect 42380 577360 42430 577416
rect 42430 577360 42444 577416
rect 42380 577356 42444 577360
rect 40540 576812 40604 576876
rect 676996 575996 677060 576060
rect 676812 572732 676876 572796
rect 42380 572596 42444 572660
rect 41828 572188 41892 572252
rect 41460 571916 41524 571980
rect 671476 571100 671540 571164
rect 41644 570964 41708 571028
rect 675340 563136 675404 563140
rect 675340 563080 675390 563136
rect 675390 563080 675404 563136
rect 675340 563076 675404 563080
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676812 557500 676876 557564
rect 42012 553012 42076 553076
rect 42196 551788 42260 551852
rect 677180 550700 677244 550764
rect 675524 546484 675588 546548
rect 676076 546484 676140 546548
rect 41644 546348 41708 546412
rect 675340 545940 675404 546004
rect 40540 545668 40604 545732
rect 40724 545396 40788 545460
rect 40540 536964 40604 537028
rect 40724 535196 40788 535260
rect 41460 530572 41524 530636
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 41644 529076 41708 529140
rect 674420 527036 674484 527100
rect 676812 503644 676876 503708
rect 677364 492416 677428 492420
rect 677364 492360 677378 492416
rect 677378 492360 677428 492416
rect 677364 492356 677428 492360
rect 675892 490452 675956 490516
rect 675892 488820 675956 488884
rect 673684 475356 673748 475420
rect 674052 475356 674116 475420
rect 673684 464748 673748 464812
rect 673868 455092 673932 455156
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 41460 418780 41524 418844
rect 40724 418508 40788 418572
rect 40540 418236 40604 418300
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 676996 402868 677060 402932
rect 41828 401840 41892 401844
rect 41828 401784 41842 401840
rect 41842 401784 41892 401840
rect 41828 401780 41892 401784
rect 676812 401236 676876 401300
rect 41460 398788 41524 398852
rect 675892 398788 675956 398852
rect 676260 396748 676324 396812
rect 676628 395116 676692 395180
rect 676444 394708 676508 394772
rect 676076 393076 676140 393140
rect 675708 387636 675772 387700
rect 676260 384916 676324 384980
rect 41460 381788 41524 381852
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 675892 377436 675956 377500
rect 676628 377164 676692 377228
rect 41644 376892 41708 376956
rect 41276 373220 41340 373284
rect 676076 372948 676140 373012
rect 674788 372540 674852 372604
rect 41828 371860 41892 371924
rect 41276 368460 41340 368524
rect 40724 363564 40788 363628
rect 40540 360028 40604 360092
rect 41828 359408 41892 359412
rect 41828 359352 41842 359408
rect 41842 359352 41892 359408
rect 41828 359348 41892 359352
rect 41460 358668 41524 358732
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43852 354240 43916 354244
rect 43852 354184 43902 354240
rect 43902 354184 43916 354240
rect 43852 354180 43916 354184
rect 675340 354180 675404 354244
rect 44220 353772 44284 353836
rect 675708 352956 675772 353020
rect 675892 351732 675956 351796
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675892 349208 675956 349212
rect 675892 349152 675942 349208
rect 675942 349152 675956 349208
rect 675892 349148 675956 349152
rect 44404 342892 44468 342956
rect 44220 342484 44284 342548
rect 44588 342076 44652 342140
rect 44404 341260 44468 341324
rect 43668 340444 43732 340508
rect 676628 340308 676692 340372
rect 675340 339008 675404 339012
rect 675340 338952 675390 339008
rect 675390 338952 675404 339008
rect 675340 338948 675404 338952
rect 40724 337724 40788 337788
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 42748 337588 42812 337652
rect 42932 336772 42996 336836
rect 676444 336636 676508 336700
rect 43116 336092 43180 336156
rect 40540 335684 40604 335748
rect 42564 335412 42628 335476
rect 41276 335276 41340 335340
rect 42564 334596 42628 334660
rect 43116 334656 43180 334660
rect 43116 334600 43166 334656
rect 43166 334600 43180 334656
rect 43116 334596 43180 334600
rect 40908 333644 40972 333708
rect 676260 332148 676324 332212
rect 41644 329020 41708 329084
rect 42012 328340 42076 328404
rect 676076 328340 676140 328404
rect 40724 326708 40788 326772
rect 40908 325348 40972 325412
rect 41460 324668 41524 324732
rect 40540 321132 40604 321196
rect 43116 316372 43180 316436
rect 41828 315616 41892 315620
rect 41828 315560 41878 315616
rect 41878 315560 41892 315616
rect 41828 315556 41892 315560
rect 42932 312700 42996 312764
rect 42012 312624 42076 312628
rect 42012 312568 42062 312624
rect 42062 312568 42076 312624
rect 42012 312564 42076 312568
rect 44220 311476 44284 311540
rect 44404 311264 44468 311268
rect 44404 311208 44418 311264
rect 44418 311208 44468 311264
rect 44404 311204 44468 311208
rect 44588 311128 44652 311132
rect 44588 311072 44602 311128
rect 44602 311072 44652 311128
rect 44588 311068 44652 311072
rect 675708 308756 675772 308820
rect 675892 306716 675956 306780
rect 675892 302636 675956 302700
rect 676444 301608 676508 301612
rect 676444 301552 676458 301608
rect 676458 301552 676508 301608
rect 676444 301548 676508 301552
rect 676628 301472 676692 301476
rect 676628 301416 676678 301472
rect 676678 301416 676692 301472
rect 676628 301412 676692 301416
rect 43668 297604 43732 297668
rect 675708 297332 675772 297396
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676260 295156 676324 295220
rect 40540 292528 40604 292592
rect 40908 292528 40972 292592
rect 41828 292496 41892 292500
rect 41828 292440 41842 292496
rect 41842 292440 41892 292496
rect 41828 292436 41892 292440
rect 676444 291484 676508 291548
rect 41828 290456 41892 290460
rect 41828 290400 41842 290456
rect 41842 290400 41892 290456
rect 41828 290396 41892 290400
rect 676628 286996 676692 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 40724 278428 40788 278492
rect 40908 277884 40972 277948
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 674972 263604 675036 263668
rect 676076 262380 676140 262444
rect 676996 261564 677060 261628
rect 676812 259932 676876 259996
rect 40724 251364 40788 251428
rect 676996 250276 677060 250340
rect 40540 249732 40604 249796
rect 674788 249596 674852 249660
rect 676076 249596 676140 249660
rect 676812 245244 676876 245308
rect 675156 244972 675220 245036
rect 675340 244700 675404 244764
rect 675156 240272 675220 240276
rect 675156 240216 675206 240272
rect 675206 240216 675220 240272
rect 675156 240212 675220 240216
rect 40724 240076 40788 240140
rect 42012 238036 42076 238100
rect 675340 236872 675404 236876
rect 675340 236816 675390 236872
rect 675390 236816 675404 236872
rect 675340 236812 675404 236816
rect 40540 235860 40604 235924
rect 674236 233140 674300 233204
rect 673684 231372 673748 231436
rect 673132 230284 673196 230348
rect 673316 230344 673380 230348
rect 673316 230288 673366 230344
rect 673366 230288 673380 230344
rect 673316 230284 673380 230288
rect 667980 229800 668044 229804
rect 667980 229744 667994 229800
rect 667994 229744 668044 229800
rect 667980 229740 668044 229744
rect 668164 229740 668228 229804
rect 668164 229196 668228 229260
rect 672948 228712 673012 228716
rect 672948 228656 672962 228712
rect 672962 228656 673012 228712
rect 672948 228652 673012 228656
rect 675156 228516 675220 228580
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 671108 227216 671172 227220
rect 671108 227160 671122 227216
rect 671122 227160 671172 227216
rect 671108 227156 671172 227160
rect 675340 226748 675404 226812
rect 672028 226612 672092 226676
rect 673500 226476 673564 226540
rect 671660 226340 671724 226404
rect 672028 226068 672092 226132
rect 673684 225116 673748 225180
rect 671660 224980 671724 225044
rect 673500 224844 673564 224908
rect 673132 224300 673196 224364
rect 671108 224028 671172 224092
rect 673316 224028 673380 224092
rect 673500 223620 673564 223684
rect 565676 222592 565740 222596
rect 565676 222536 565726 222592
rect 565726 222536 565740 222592
rect 565676 222532 565740 222536
rect 572484 221988 572548 222052
rect 672028 221036 672092 221100
rect 670740 220900 670804 220964
rect 572484 220628 572548 220692
rect 540100 220492 540164 220556
rect 563652 220492 563716 220556
rect 511028 220008 511092 220012
rect 511028 219952 511042 220008
rect 511042 219952 511092 220008
rect 511028 219948 511092 219952
rect 526484 220008 526548 220012
rect 526484 219952 526498 220008
rect 526498 219952 526548 220008
rect 519860 219736 519924 219740
rect 519860 219680 519874 219736
rect 519874 219680 519924 219736
rect 519860 219676 519924 219680
rect 522620 219736 522684 219740
rect 526484 219948 526548 219952
rect 554084 220220 554148 220284
rect 522620 219680 522634 219736
rect 522634 219680 522684 219736
rect 522620 219676 522684 219680
rect 562548 219676 562612 219740
rect 568620 219676 568684 219740
rect 672028 219872 672092 219876
rect 672028 219816 672042 219872
rect 672042 219816 672092 219872
rect 672028 219812 672092 219816
rect 675524 219948 675588 220012
rect 572668 219132 572732 219196
rect 572852 219132 572916 219196
rect 562180 218316 562244 218380
rect 562916 218588 562980 218652
rect 675524 218860 675588 218924
rect 674972 218588 675036 218652
rect 575060 218180 575124 218244
rect 675892 218180 675956 218244
rect 563284 217908 563348 217972
rect 504404 217500 504468 217564
rect 508268 217772 508332 217836
rect 562732 217772 562796 217836
rect 563100 217500 563164 217564
rect 565676 217424 565740 217428
rect 565676 217368 565680 217424
rect 565680 217368 565736 217424
rect 565736 217368 565740 217424
rect 565676 217364 565740 217368
rect 567700 217398 567764 217462
rect 493548 217288 493612 217292
rect 493548 217232 493598 217288
rect 493598 217232 493612 217288
rect 493548 217228 493612 217232
rect 508268 216956 508332 217020
rect 675524 217364 675588 217428
rect 675156 217228 675220 217292
rect 675708 216956 675772 217020
rect 675340 216820 675404 216884
rect 504404 216140 504468 216204
rect 519308 216412 519372 216476
rect 519860 216412 519924 216476
rect 564940 216412 565004 216476
rect 566596 216412 566660 216476
rect 511028 216140 511092 216204
rect 519308 215868 519372 215932
rect 536052 215868 536116 215932
rect 522620 215596 522684 215660
rect 526484 215324 526548 215388
rect 538812 215460 538876 215524
rect 539180 215460 539244 215524
rect 546724 215596 546788 215660
rect 547644 215596 547708 215660
rect 548196 215596 548260 215660
rect 548380 215596 548444 215660
rect 556476 215596 556540 215660
rect 558868 215596 558932 215660
rect 566412 215596 566476 215660
rect 539916 215324 539980 215388
rect 572484 215596 572548 215660
rect 572852 215868 572916 215932
rect 583708 215868 583772 215932
rect 536052 215052 536116 215116
rect 538996 215052 539060 215116
rect 540100 215052 540164 215116
rect 546908 215052 546972 215116
rect 548196 215052 548260 215116
rect 567884 215324 567948 215388
rect 566964 215052 567028 215116
rect 568252 215052 568316 215116
rect 576716 215324 576780 215388
rect 676076 215086 676140 215150
rect 575612 214916 575676 214980
rect 673132 214644 673196 214708
rect 675892 214508 675956 214572
rect 674052 212060 674116 212124
rect 675892 211380 675956 211444
rect 676444 211380 676508 211444
rect 669452 211108 669516 211172
rect 674972 210428 675036 210492
rect 675892 210428 675956 210492
rect 41460 209748 41524 209812
rect 40724 208116 40788 208180
rect 42012 207708 42076 207772
rect 40908 207300 40972 207364
rect 40540 206892 40604 206956
rect 676628 205532 676692 205596
rect 676444 200636 676508 200700
rect 675524 198248 675588 198252
rect 675524 198192 675574 198248
rect 675574 198192 675588 198248
rect 675524 198188 675588 198192
rect 41828 197780 41892 197844
rect 40724 197100 40788 197164
rect 676260 197100 676324 197164
rect 41828 195800 41892 195804
rect 41828 195744 41878 195800
rect 41878 195744 41892 195800
rect 41828 195740 41892 195744
rect 40908 195468 40972 195532
rect 41460 195196 41524 195260
rect 40540 194516 40604 194580
rect 41644 194516 41708 194580
rect 675892 193156 675956 193220
rect 42380 192884 42444 192948
rect 676076 191524 676140 191588
rect 41828 187232 41892 187236
rect 41828 187176 41842 187232
rect 41842 187176 41892 187232
rect 41828 187172 41892 187176
rect 42380 186144 42444 186148
rect 42380 186088 42394 186144
rect 42394 186088 42444 186144
rect 42380 186084 42444 186088
rect 42012 185872 42076 185876
rect 42012 185816 42026 185872
rect 42026 185816 42076 185872
rect 42012 185812 42076 185816
rect 672948 183500 673012 183564
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675892 171940 675956 172004
rect 675524 167452 675588 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 673132 164188 673196 164252
rect 675340 161876 675404 161940
rect 676444 159292 676508 159356
rect 675340 157040 675404 157044
rect 675340 156984 675390 157040
rect 675390 156984 675404 157040
rect 675340 156980 675404 156984
rect 676628 156300 676692 156364
rect 674236 154532 674300 154596
rect 676260 153036 676324 153100
rect 675892 148412 675956 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 676076 145964 676140 146028
rect 669268 143516 669332 143580
rect 670740 133724 670804 133788
rect 667980 130460 668044 130524
rect 673500 128828 673564 128892
rect 676628 128556 676692 128620
rect 674052 128284 674116 128348
rect 676076 128148 676140 128212
rect 675892 127196 675956 127260
rect 676260 126924 676324 126988
rect 676444 124476 676508 124540
rect 675708 122300 675772 122364
rect 676628 113052 676692 113116
rect 675892 108020 675956 108084
rect 676444 106116 676508 106180
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676260 101356 676324 101420
rect 634860 96596 634924 96660
rect 637252 96596 637316 96660
rect 634860 80412 634924 80476
rect 637068 77828 637132 77892
rect 461716 54980 461780 55044
rect 462636 54436 462700 54500
rect 461716 53892 461780 53956
rect 462636 53892 462700 53956
rect 194364 50220 194428 50284
rect 529796 50220 529860 50284
rect 308996 49676 309060 49740
rect 518756 48860 518820 48924
rect 526484 48044 526548 48108
rect 520964 47772 521028 47836
rect 515444 47500 515508 47564
rect 522068 47228 522132 47292
rect 461348 44372 461412 44436
rect 462268 44372 462332 44436
rect 141740 43964 141804 44028
rect 440188 43828 440252 43892
rect 440924 43828 440988 43892
rect 308996 42800 309060 42804
rect 308996 42744 309010 42800
rect 309010 42744 309060 42800
rect 308996 42740 309060 42744
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529796 42060 529860 42124
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
rect 141740 40488 141804 40492
rect 141740 40432 141754 40488
rect 141754 40432 141804 40488
rect 141740 40428 141804 40432
<< metal4 >>
rect 524091 997796 524157 997797
rect 524091 997732 524092 997796
rect 524156 997732 524157 997796
rect 524091 997731 524157 997732
rect 524094 997338 524154 997731
rect 89483 997252 89549 997253
rect 89483 997188 89484 997252
rect 89548 997188 89549 997252
rect 195283 997252 195349 997253
rect 195283 997250 195284 997252
rect 89483 997187 89549 997188
rect 194918 997190 195284 997250
rect 89486 995621 89546 997187
rect 189763 997116 189829 997117
rect 189763 997052 189764 997116
rect 189828 997052 189829 997116
rect 189763 997051 189829 997052
rect 188107 996436 188173 996437
rect 188107 996372 188108 996436
rect 188172 996372 188173 996436
rect 188107 996371 188173 996372
rect 89851 996300 89917 996301
rect 89851 996236 89852 996300
rect 89916 996236 89917 996300
rect 89851 996235 89917 996236
rect 140083 996300 140149 996301
rect 140083 996236 140084 996300
rect 140148 996236 140149 996300
rect 140083 996235 140149 996236
rect 89854 995890 89914 996235
rect 132355 996028 132421 996029
rect 132355 995964 132356 996028
rect 132420 995964 132421 996028
rect 132355 995963 132421 995964
rect 89670 995830 89914 995890
rect 89299 995620 89365 995621
rect 89299 995556 89300 995620
rect 89364 995556 89365 995620
rect 89299 995555 89365 995556
rect 89483 995620 89549 995621
rect 89483 995556 89484 995620
rect 89548 995556 89549 995620
rect 89483 995555 89549 995556
rect 89302 995210 89362 995555
rect 89670 995210 89730 995830
rect 132358 995349 132418 995963
rect 140086 995890 140146 996235
rect 140086 995830 140882 995890
rect 132539 995756 132605 995757
rect 132539 995692 132540 995756
rect 132604 995692 132605 995756
rect 132539 995691 132605 995692
rect 132355 995348 132421 995349
rect 132355 995284 132356 995348
rect 132420 995284 132421 995348
rect 132355 995283 132421 995284
rect 89302 995150 89730 995210
rect 132542 993853 132602 995691
rect 140822 995349 140882 995830
rect 188110 995757 188170 996371
rect 189766 995757 189826 997051
rect 194918 996709 194978 997190
rect 195283 997188 195284 997190
rect 195348 997188 195349 997252
rect 195283 997187 195349 997188
rect 243491 997252 243557 997253
rect 243491 997188 243492 997252
rect 243556 997188 243557 997252
rect 243491 997187 243557 997188
rect 287835 997252 287901 997253
rect 287835 997188 287836 997252
rect 287900 997188 287901 997252
rect 287835 997187 287901 997188
rect 385907 997252 385973 997253
rect 385907 997188 385908 997252
rect 385972 997188 385973 997252
rect 385907 997187 385973 997188
rect 194915 996708 194981 996709
rect 194915 996644 194916 996708
rect 194980 996644 194981 996708
rect 194915 996643 194981 996644
rect 192339 996436 192405 996437
rect 192339 996372 192340 996436
rect 192404 996372 192405 996436
rect 192339 996371 192405 996372
rect 191603 996028 191669 996029
rect 191603 995964 191604 996028
rect 191668 995964 191669 996028
rect 191603 995963 191669 995964
rect 188107 995756 188173 995757
rect 188107 995692 188108 995756
rect 188172 995692 188173 995756
rect 188107 995691 188173 995692
rect 189763 995756 189829 995757
rect 189763 995692 189764 995756
rect 189828 995692 189829 995756
rect 189763 995691 189829 995692
rect 140819 995348 140885 995349
rect 140819 995284 140820 995348
rect 140884 995284 140885 995348
rect 140819 995283 140885 995284
rect 191606 994805 191666 995963
rect 192342 995621 192402 996371
rect 243494 995757 243554 997187
rect 243859 996980 243925 996981
rect 243859 996916 243860 996980
rect 243924 996916 243925 996980
rect 243859 996915 243925 996916
rect 243862 995757 243922 996915
rect 243491 995756 243557 995757
rect 243491 995692 243492 995756
rect 243556 995692 243557 995756
rect 243491 995691 243557 995692
rect 243859 995756 243925 995757
rect 243859 995692 243860 995756
rect 243924 995692 243925 995756
rect 243859 995691 243925 995692
rect 192339 995620 192405 995621
rect 192339 995556 192340 995620
rect 192404 995556 192405 995620
rect 192339 995555 192405 995556
rect 287838 994805 287898 997187
rect 295379 996980 295445 996981
rect 295379 996916 295380 996980
rect 295444 996916 295445 996980
rect 295379 996915 295445 996916
rect 291515 996708 291581 996709
rect 291515 996644 291516 996708
rect 291580 996644 291581 996708
rect 291515 996643 291581 996644
rect 291518 994805 291578 996643
rect 292251 996164 292317 996165
rect 292251 996100 292252 996164
rect 292316 996100 292317 996164
rect 292251 996099 292317 996100
rect 292254 995890 292314 996099
rect 292254 995830 292498 995890
rect 292438 995621 292498 995830
rect 295382 995757 295442 996915
rect 385355 996300 385421 996301
rect 385355 996236 385356 996300
rect 385420 996236 385421 996300
rect 385355 996235 385421 996236
rect 364195 995892 364261 995893
rect 364195 995828 364196 995892
rect 364260 995828 364261 995892
rect 364195 995827 364261 995828
rect 295379 995756 295445 995757
rect 295379 995692 295380 995756
rect 295444 995692 295445 995756
rect 295379 995691 295445 995692
rect 292435 995620 292501 995621
rect 292435 995556 292436 995620
rect 292500 995556 292501 995620
rect 292435 995555 292501 995556
rect 191603 994804 191669 994805
rect 191603 994740 191604 994804
rect 191668 994740 191669 994804
rect 191603 994739 191669 994740
rect 287835 994804 287901 994805
rect 287835 994740 287836 994804
rect 287900 994740 287901 994804
rect 287835 994739 287901 994740
rect 291515 994804 291581 994805
rect 291515 994740 291516 994804
rect 291580 994740 291581 994804
rect 291515 994739 291581 994740
rect 132539 993852 132605 993853
rect 132539 993788 132540 993852
rect 132604 993788 132605 993852
rect 132539 993787 132605 993788
rect 141926 993790 142354 993850
rect 141926 993445 141986 993790
rect 142294 993445 142354 993790
rect 141923 993444 141989 993445
rect 141923 993380 141924 993444
rect 141988 993380 141989 993444
rect 141923 993379 141989 993380
rect 142291 993444 142357 993445
rect 142291 993380 142292 993444
rect 142356 993380 142357 993444
rect 142291 993379 142357 993380
rect 364198 993258 364258 995827
rect 385358 995043 385418 996235
rect 385355 995042 385421 995043
rect 385355 994978 385356 995042
rect 385420 994978 385421 995042
rect 385355 994977 385421 994978
rect 385910 994941 385970 997187
rect 532555 997252 532621 997253
rect 532555 997188 532556 997252
rect 532620 997188 532621 997252
rect 532555 997187 532621 997188
rect 388667 996708 388733 996709
rect 388667 996644 388668 996708
rect 388732 996644 388733 996708
rect 388667 996643 388733 996644
rect 388670 995757 388730 996643
rect 396579 996436 396645 996437
rect 396579 996372 396580 996436
rect 396644 996372 396645 996436
rect 396579 996371 396645 996372
rect 388483 995756 388549 995757
rect 388483 995692 388484 995756
rect 388548 995692 388549 995756
rect 388483 995691 388549 995692
rect 388667 995756 388733 995757
rect 388667 995692 388668 995756
rect 388732 995692 388733 995756
rect 388667 995691 388733 995692
rect 388486 995077 388546 995691
rect 396582 995485 396642 996371
rect 484347 996300 484413 996301
rect 484347 996236 484348 996300
rect 484412 996236 484413 996300
rect 484347 996235 484413 996236
rect 484350 995757 484410 996235
rect 484347 995756 484413 995757
rect 484347 995692 484348 995756
rect 484412 995692 484413 995756
rect 484347 995691 484413 995692
rect 393451 995484 393517 995485
rect 393451 995420 393452 995484
rect 393516 995420 393517 995484
rect 393451 995419 393517 995420
rect 396579 995484 396645 995485
rect 396579 995420 396580 995484
rect 396644 995420 396645 995484
rect 396579 995419 396645 995420
rect 393454 995210 393514 995419
rect 393086 995150 393514 995210
rect 388483 995076 388549 995077
rect 388483 995012 388484 995076
rect 388548 995012 388549 995076
rect 388483 995011 388549 995012
rect 385907 994940 385973 994941
rect 385907 994876 385908 994940
rect 385972 994876 385973 994940
rect 385907 994875 385973 994876
rect 393086 993258 393146 995150
rect 522806 995077 522866 997102
rect 529795 996708 529861 996709
rect 529795 996644 529796 996708
rect 529860 996644 529861 996708
rect 529795 996643 529861 996644
rect 529798 995621 529858 996643
rect 532006 995757 532066 997102
rect 532558 995757 532618 997187
rect 630259 997252 630325 997253
rect 630259 997188 630260 997252
rect 630324 997188 630325 997252
rect 630259 997187 630325 997188
rect 538259 996708 538325 996709
rect 538259 996644 538260 996708
rect 538324 996644 538325 996708
rect 538259 996643 538325 996644
rect 627867 996708 627933 996709
rect 627867 996644 627868 996708
rect 627932 996644 627933 996708
rect 627867 996643 627933 996644
rect 532003 995756 532069 995757
rect 532003 995692 532004 995756
rect 532068 995692 532069 995756
rect 532003 995691 532069 995692
rect 532555 995756 532621 995757
rect 532555 995692 532556 995756
rect 532620 995692 532621 995756
rect 532555 995691 532621 995692
rect 529795 995620 529861 995621
rect 529795 995556 529796 995620
rect 529860 995556 529861 995620
rect 529795 995555 529861 995556
rect 522803 995076 522869 995077
rect 522803 995012 522804 995076
rect 522868 995012 522869 995076
rect 522803 995011 522869 995012
rect 538262 994533 538322 996643
rect 627870 995757 627930 996643
rect 630262 995757 630322 997187
rect 633939 996980 634005 996981
rect 633939 996916 633940 996980
rect 634004 996916 634005 996980
rect 633939 996915 634005 996916
rect 633942 995757 634002 996915
rect 636702 995757 636762 997102
rect 627867 995756 627933 995757
rect 627867 995692 627868 995756
rect 627932 995692 627933 995756
rect 627867 995691 627933 995692
rect 630259 995756 630325 995757
rect 630259 995692 630260 995756
rect 630324 995692 630325 995756
rect 630259 995691 630325 995692
rect 633939 995756 634005 995757
rect 633939 995692 633940 995756
rect 634004 995692 634005 995756
rect 633939 995691 634005 995692
rect 636699 995756 636765 995757
rect 636699 995692 636700 995756
rect 636764 995692 636765 995756
rect 636699 995691 636765 995692
rect 538259 994532 538325 994533
rect 538259 994468 538260 994532
rect 538324 994468 538325 994532
rect 538259 994467 538325 994468
rect 41459 967196 41525 967197
rect 41459 967132 41460 967196
rect 41524 967132 41525 967196
rect 41459 967131 41525 967132
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 946710 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 40358 946650 40602 946710
rect 40358 944077 40418 946650
rect 40355 944076 40421 944077
rect 40355 944012 40356 944076
rect 40420 944012 40421 944076
rect 40355 944011 40421 944012
rect 40726 943805 40786 955435
rect 41278 951693 41338 959787
rect 41462 952509 41522 967131
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675339 963388 675405 963389
rect 675339 963324 675340 963388
rect 675404 963324 675405 963388
rect 675339 963323 675405 963324
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 959130 41890 962099
rect 675155 959308 675221 959309
rect 675155 959244 675156 959308
rect 675220 959244 675221 959308
rect 675155 959243 675221 959244
rect 41646 959070 41890 959130
rect 41459 952508 41525 952509
rect 41459 952444 41460 952508
rect 41524 952444 41525 952508
rect 41459 952443 41525 952444
rect 41646 952237 41706 959070
rect 41827 957812 41893 957813
rect 41827 957748 41828 957812
rect 41892 957748 41893 957812
rect 41827 957747 41893 957748
rect 41830 952917 41890 957747
rect 41827 952916 41893 952917
rect 41827 952852 41828 952916
rect 41892 952852 41893 952916
rect 41827 952851 41893 952852
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 41275 951692 41341 951693
rect 41275 951628 41276 951692
rect 41340 951628 41341 951692
rect 41275 951627 41341 951628
rect 675158 951149 675218 959243
rect 675342 954549 675402 963323
rect 675339 954548 675405 954549
rect 675339 954484 675340 954548
rect 675404 954484 675405 954548
rect 675339 954483 675405 954484
rect 675155 951148 675221 951149
rect 675155 951084 675156 951148
rect 675220 951084 675221 951148
rect 675155 951083 675221 951084
rect 676078 950741 676138 965091
rect 676627 963660 676693 963661
rect 676627 963596 676628 963660
rect 676692 963596 676693 963660
rect 676627 963595 676693 963596
rect 676630 951557 676690 963595
rect 676811 957812 676877 957813
rect 676811 957748 676812 957812
rect 676876 957748 676877 957812
rect 676811 957747 676877 957748
rect 676627 951556 676693 951557
rect 676627 951492 676628 951556
rect 676692 951492 676693 951556
rect 676627 951491 676693 951492
rect 676075 950740 676141 950741
rect 676075 950676 676076 950740
rect 676140 950676 676141 950740
rect 676075 950675 676141 950676
rect 42195 944076 42261 944077
rect 42195 944012 42196 944076
rect 42260 944012 42261 944076
rect 42195 944011 42261 944012
rect 40723 943804 40789 943805
rect 40723 943740 40724 943804
rect 40788 943740 40789 943804
rect 40723 943739 40789 943740
rect 42011 943804 42077 943805
rect 42011 943740 42012 943804
rect 42076 943740 42077 943804
rect 42011 943739 42077 943740
rect 41827 939452 41893 939453
rect 41827 939450 41828 939452
rect 40542 939390 41828 939450
rect 40542 935670 40602 939390
rect 41827 939388 41828 939390
rect 41892 939388 41893 939452
rect 41827 939387 41893 939388
rect 42014 937050 42074 943739
rect 41830 936990 42074 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 41827 935780 41893 935781
rect 41827 935716 41828 935780
rect 41892 935778 41893 935780
rect 42198 935778 42258 944011
rect 41892 935718 42258 935778
rect 41892 935716 41893 935718
rect 41827 935715 41893 935716
rect 39990 935610 40602 935670
rect 39990 814299 40050 935610
rect 676814 931565 676874 957747
rect 676995 956452 677061 956453
rect 676995 956388 676996 956452
rect 677060 956388 677061 956452
rect 676995 956387 677061 956388
rect 676998 931973 677058 956387
rect 676995 931972 677061 931973
rect 676995 931908 676996 931972
rect 677060 931908 677061 931972
rect 676995 931907 677061 931908
rect 676811 931564 676877 931565
rect 676811 931500 676812 931564
rect 676876 931500 676877 931564
rect 676811 931499 676877 931500
rect 42011 911980 42077 911981
rect 42011 911916 42012 911980
rect 42076 911916 42077 911980
rect 42011 911915 42077 911916
rect 42014 885461 42074 911915
rect 42195 911708 42261 911709
rect 42195 911644 42196 911708
rect 42260 911644 42261 911708
rect 42195 911643 42261 911644
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911643
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 673867 873220 673933 873221
rect 673867 873156 673868 873220
rect 673932 873156 673933 873220
rect 673867 873155 673933 873156
rect 39987 814298 40053 814299
rect 39987 814234 39988 814298
rect 40052 814234 40053 814298
rect 39987 814233 40053 814234
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40723 805492 40789 805493
rect 40723 805428 40724 805492
rect 40788 805428 40789 805492
rect 40723 805427 40789 805428
rect 40539 804812 40605 804813
rect 40539 804748 40540 804812
rect 40604 804748 40605 804812
rect 40539 804747 40605 804748
rect 40542 792573 40602 804747
rect 40726 794205 40786 805427
rect 40907 805084 40973 805085
rect 40907 805020 40908 805084
rect 40972 805020 40973 805084
rect 40907 805019 40973 805020
rect 40910 795429 40970 805019
rect 40907 795428 40973 795429
rect 40907 795364 40908 795428
rect 40972 795364 40973 795428
rect 40907 795363 40973 795364
rect 40723 794204 40789 794205
rect 40723 794140 40724 794204
rect 40788 794140 40789 794204
rect 40723 794139 40789 794140
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 786861 41522 812910
rect 42195 808756 42261 808757
rect 42195 808692 42196 808756
rect 42260 808692 42261 808756
rect 42195 808691 42261 808692
rect 42011 805628 42077 805629
rect 42011 805564 42012 805628
rect 42076 805564 42077 805628
rect 42011 805563 42077 805564
rect 41643 805356 41709 805357
rect 41643 805292 41644 805356
rect 41708 805292 41709 805356
rect 41643 805291 41709 805292
rect 41646 789037 41706 805291
rect 42014 794910 42074 805563
rect 42198 804813 42258 808691
rect 42195 804812 42261 804813
rect 42195 804748 42196 804812
rect 42260 804748 42261 804812
rect 42195 804747 42261 804748
rect 41830 794850 42074 794910
rect 41643 789036 41709 789037
rect 41643 788972 41644 789036
rect 41708 788972 41709 789036
rect 41643 788971 41709 788972
rect 41830 788629 41890 794850
rect 41827 788628 41893 788629
rect 41827 788564 41828 788628
rect 41892 788564 41893 788628
rect 41827 788563 41893 788564
rect 41459 786860 41525 786861
rect 41459 786796 41460 786860
rect 41524 786796 41525 786860
rect 41459 786795 41525 786796
rect 673870 770949 673930 873155
rect 675342 863157 675402 873971
rect 675339 863156 675405 863157
rect 675339 863092 675340 863156
rect 675404 863092 675405 863156
rect 675339 863091 675405 863092
rect 675523 777068 675589 777069
rect 675523 777004 675524 777068
rect 675588 777004 675589 777068
rect 675523 777003 675589 777004
rect 675526 775709 675586 777003
rect 675523 775708 675589 775709
rect 675523 775644 675524 775708
rect 675588 775644 675589 775708
rect 675523 775643 675589 775644
rect 675707 775572 675773 775573
rect 675707 775508 675708 775572
rect 675772 775508 675773 775572
rect 675707 775507 675773 775508
rect 675710 774349 675770 775507
rect 675707 774348 675773 774349
rect 675707 774284 675708 774348
rect 675772 774284 675773 774348
rect 675707 774283 675773 774284
rect 676078 772717 676138 875875
rect 676811 870908 676877 870909
rect 676811 870844 676812 870908
rect 676876 870844 676877 870908
rect 676811 870843 676877 870844
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 673867 770948 673933 770949
rect 673867 770884 673868 770948
rect 673932 770884 673933 770948
rect 673867 770883 673933 770884
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40542 747421 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750413 40786 764899
rect 40910 754901 40970 765715
rect 40907 754900 40973 754901
rect 40907 754836 40908 754900
rect 40972 754836 40973 754900
rect 40907 754835 40973 754836
rect 40723 750412 40789 750413
rect 40723 750348 40724 750412
rect 40788 750348 40789 750412
rect 40723 750347 40789 750348
rect 40539 747420 40605 747421
rect 40539 747356 40540 747420
rect 40604 747356 40605 747420
rect 40539 747355 40605 747356
rect 41462 743749 41522 769795
rect 675155 768228 675221 768229
rect 675155 768164 675156 768228
rect 675220 768164 675221 768228
rect 675155 768163 675221 768164
rect 675158 765930 675218 768163
rect 676075 766596 676141 766597
rect 676075 766532 676076 766596
rect 676140 766532 676141 766596
rect 676075 766531 676141 766532
rect 675158 765870 675954 765930
rect 41643 764556 41709 764557
rect 41643 764492 41644 764556
rect 41708 764492 41709 764556
rect 41643 764491 41709 764492
rect 41646 745109 41706 764491
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41643 745108 41709 745109
rect 41643 745044 41644 745108
rect 41708 745044 41709 745108
rect 41643 745043 41709 745044
rect 41830 744837 41890 757691
rect 42011 756396 42077 756397
rect 42011 756332 42012 756396
rect 42076 756332 42077 756396
rect 42011 756331 42077 756332
rect 42014 754085 42074 756331
rect 42011 754084 42077 754085
rect 42011 754020 42012 754084
rect 42076 754020 42077 754084
rect 42011 754019 42077 754020
rect 42195 753268 42261 753269
rect 42195 753204 42196 753268
rect 42260 753204 42261 753268
rect 42195 753203 42261 753204
rect 42198 751773 42258 753203
rect 42195 751772 42261 751773
rect 42195 751708 42196 751772
rect 42260 751708 42261 751772
rect 42195 751707 42261 751708
rect 41827 744836 41893 744837
rect 41827 744772 41828 744836
rect 41892 744772 41893 744836
rect 41827 744771 41893 744772
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674419 742524 674485 742525
rect 674419 742460 674420 742524
rect 674484 742460 674485 742524
rect 674419 742459 674485 742460
rect 674235 741572 674301 741573
rect 674235 741508 674236 741572
rect 674300 741508 674301 741572
rect 674235 741507 674301 741508
rect 672027 732868 672093 732869
rect 672027 732804 672028 732868
rect 672092 732804 672093 732868
rect 672027 732803 672093 732804
rect 673315 732868 673381 732869
rect 673315 732804 673316 732868
rect 673380 732804 673381 732868
rect 673315 732803 673381 732804
rect 672030 728245 672090 732803
rect 673318 728517 673378 732803
rect 673315 728516 673381 728517
rect 673315 728452 673316 728516
rect 673380 728452 673381 728516
rect 673315 728451 673381 728452
rect 672027 728244 672093 728245
rect 672027 728180 672028 728244
rect 672092 728180 672093 728244
rect 672027 728179 672093 728180
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 706485 40602 718523
rect 40726 707437 40786 721707
rect 41275 714236 41341 714237
rect 41275 714172 41276 714236
rect 41340 714172 41341 714236
rect 41275 714171 41341 714172
rect 41278 712197 41338 714171
rect 41275 712196 41341 712197
rect 41275 712132 41276 712196
rect 41340 712132 41341 712196
rect 41275 712131 41341 712132
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 40539 706484 40605 706485
rect 40539 706420 40540 706484
rect 40604 706420 40605 706484
rect 40539 706419 40605 706420
rect 41462 700501 41522 726550
rect 41827 722396 41893 722397
rect 41827 722332 41828 722396
rect 41892 722332 41893 722396
rect 41827 722331 41893 722332
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41646 702405 41706 721707
rect 41830 718589 41890 722331
rect 41827 718588 41893 718589
rect 41827 718524 41828 718588
rect 41892 718524 41893 718588
rect 41827 718523 41893 718524
rect 42011 714780 42077 714781
rect 42011 714716 42012 714780
rect 42076 714716 42077 714780
rect 42011 714715 42077 714716
rect 41827 714508 41893 714509
rect 41827 714444 41828 714508
rect 41892 714444 41893 714508
rect 41827 714443 41893 714444
rect 41830 709885 41890 714443
rect 41827 709884 41893 709885
rect 41827 709820 41828 709884
rect 41892 709820 41893 709884
rect 41827 709819 41893 709820
rect 42014 707970 42074 714715
rect 42379 713284 42445 713285
rect 42379 713220 42380 713284
rect 42444 713220 42445 713284
rect 42379 713219 42445 713220
rect 42014 707910 42258 707970
rect 41643 702404 41709 702405
rect 41643 702340 41644 702404
rect 41708 702340 41709 702404
rect 41643 702339 41709 702340
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 42198 699957 42258 707910
rect 42382 707437 42442 713219
rect 42379 707436 42445 707437
rect 42379 707372 42380 707436
rect 42444 707372 42445 707436
rect 42379 707371 42445 707372
rect 42195 699956 42261 699957
rect 42195 699892 42196 699956
rect 42260 699892 42261 699956
rect 42195 699891 42261 699892
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683090 41890 683571
rect 41462 683030 41890 683090
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40542 664053 40602 678927
rect 40726 668269 40786 678927
rect 40723 668268 40789 668269
rect 40723 668204 40724 668268
rect 40788 668204 40789 668268
rect 40723 668203 40789 668204
rect 40539 664052 40605 664053
rect 40539 663988 40540 664052
rect 40604 663988 40605 664052
rect 40539 663987 40605 663988
rect 41462 659701 41522 683030
rect 674238 682413 674298 741507
rect 674422 682685 674482 742459
rect 674603 739668 674669 739669
rect 674603 739604 674604 739668
rect 674668 739604 674669 739668
rect 674603 739603 674669 739604
rect 674419 682684 674485 682685
rect 674419 682620 674420 682684
rect 674484 682620 674485 682684
rect 674419 682619 674485 682620
rect 674235 682412 674301 682413
rect 674235 682348 674236 682412
rect 674300 682348 674301 682412
rect 674235 682347 674301 682348
rect 41827 681052 41893 681053
rect 41827 680988 41828 681052
rect 41892 680988 41893 681052
rect 41827 680987 41893 680988
rect 41830 678990 41890 680987
rect 41646 678930 41890 678990
rect 41459 659700 41525 659701
rect 41459 659636 41460 659700
rect 41524 659636 41525 659700
rect 41459 659635 41525 659636
rect 41646 658613 41706 678930
rect 674606 673470 674666 739603
rect 675894 730013 675954 765870
rect 675891 730012 675957 730013
rect 675891 729948 675892 730012
rect 675956 729948 675957 730012
rect 675891 729947 675957 729948
rect 676078 725797 676138 766531
rect 676814 761837 676874 870843
rect 676995 774484 677061 774485
rect 676995 774420 676996 774484
rect 677060 774420 677061 774484
rect 676995 774419 677061 774420
rect 676998 761973 677058 774419
rect 676995 761972 677061 761973
rect 676995 761908 676996 761972
rect 677060 761908 677061 761972
rect 676995 761907 677061 761908
rect 676811 761836 676877 761837
rect 676811 761772 676812 761836
rect 676876 761772 676877 761836
rect 676811 761771 676877 761772
rect 676811 730012 676877 730013
rect 676811 729948 676812 730012
rect 676876 729948 676877 730012
rect 676811 729947 676877 729948
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712110 676874 729947
rect 675894 712061 676874 712110
rect 675891 712060 676874 712061
rect 675891 711996 675892 712060
rect 675956 712050 676874 712060
rect 675956 711996 675957 712050
rect 675891 711995 675957 711996
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 686493 675402 696763
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 675339 686492 675405 686493
rect 675339 686428 675340 686492
rect 675404 686428 675405 686492
rect 675339 686427 675405 686428
rect 674422 673410 674666 673470
rect 42563 673164 42629 673165
rect 42563 673100 42564 673164
rect 42628 673100 42629 673164
rect 42563 673099 42629 673100
rect 42379 672892 42445 672893
rect 42379 672828 42380 672892
rect 42444 672828 42445 672892
rect 42379 672827 42445 672828
rect 41827 671260 41893 671261
rect 41827 671196 41828 671260
rect 41892 671196 41893 671260
rect 41827 671195 41893 671196
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 671195
rect 42195 669356 42261 669357
rect 42195 669330 42196 669356
rect 42014 669292 42196 669330
rect 42260 669292 42261 669356
rect 42014 669291 42261 669292
rect 42014 669270 42258 669291
rect 42014 667725 42074 669270
rect 42011 667724 42077 667725
rect 42011 667660 42012 667724
rect 42076 667660 42077 667724
rect 42011 667659 42077 667660
rect 42382 666637 42442 672827
rect 42566 668541 42626 673099
rect 42563 668540 42629 668541
rect 42563 668476 42564 668540
rect 42628 668476 42629 668540
rect 42563 668475 42629 668476
rect 42379 666636 42445 666637
rect 42379 666572 42380 666636
rect 42444 666572 42445 666636
rect 42379 666571 42445 666572
rect 674422 664053 674482 673410
rect 674603 670172 674669 670173
rect 674603 670108 674604 670172
rect 674668 670170 674669 670172
rect 674668 670110 675034 670170
rect 674668 670108 674669 670110
rect 674603 670107 674669 670108
rect 674974 669357 675034 670110
rect 674971 669356 675037 669357
rect 674971 669292 674972 669356
rect 675036 669292 675037 669356
rect 674971 669291 675037 669292
rect 674419 664052 674485 664053
rect 674419 663988 674420 664052
rect 674484 663988 674485 664052
rect 674419 663987 674485 663988
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 44219 653172 44285 653173
rect 44219 653108 44220 653172
rect 44284 653108 44285 653172
rect 44219 653107 44285 653108
rect 41643 640660 41709 640661
rect 41643 640596 41644 640660
rect 41708 640596 41709 640660
rect 41643 640595 41709 640596
rect 41459 639436 41525 639437
rect 41459 639372 41460 639436
rect 41524 639372 41525 639436
rect 41459 639371 41525 639372
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40539 634540 40605 634541
rect 40539 634476 40540 634540
rect 40604 634476 40605 634540
rect 40539 634475 40605 634476
rect 40542 619853 40602 634475
rect 40726 622165 40786 634883
rect 40723 622164 40789 622165
rect 40723 622100 40724 622164
rect 40788 622100 40789 622164
rect 40723 622099 40789 622100
rect 40539 619852 40605 619853
rect 40539 619788 40540 619852
rect 40604 619788 40605 619852
rect 40539 619787 40605 619788
rect 41462 615501 41522 639371
rect 41646 617130 41706 640595
rect 41827 637396 41893 637397
rect 41827 637332 41828 637396
rect 41892 637332 41893 637396
rect 41827 637331 41893 637332
rect 41830 630690 41890 637331
rect 41830 630630 42074 630690
rect 41646 617070 41890 617130
rect 41459 615500 41525 615501
rect 41459 615436 41460 615500
rect 41524 615436 41525 615500
rect 41459 615435 41525 615436
rect 41830 614141 41890 617070
rect 42014 615909 42074 630630
rect 42563 626652 42629 626653
rect 42563 626588 42564 626652
rect 42628 626588 42629 626652
rect 42563 626587 42629 626588
rect 42195 625292 42261 625293
rect 42195 625228 42196 625292
rect 42260 625228 42261 625292
rect 42195 625227 42261 625228
rect 42198 623389 42258 625227
rect 42566 625021 42626 626587
rect 42563 625020 42629 625021
rect 42563 624956 42564 625020
rect 42628 624956 42629 625020
rect 42563 624955 42629 624956
rect 42195 623388 42261 623389
rect 42195 623324 42196 623388
rect 42260 623324 42261 623388
rect 42195 623323 42261 623324
rect 42011 615908 42077 615909
rect 42011 615844 42012 615908
rect 42076 615844 42077 615908
rect 42011 615843 42077 615844
rect 44222 614141 44282 653107
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674971 651540 675037 651541
rect 674971 651476 674972 651540
rect 675036 651476 675037 651540
rect 674971 651475 675037 651476
rect 674419 648956 674485 648957
rect 674419 648892 674420 648956
rect 674484 648892 674485 648956
rect 674419 648891 674485 648892
rect 674422 647597 674482 648891
rect 674419 647596 674485 647597
rect 674419 647532 674420 647596
rect 674484 647532 674485 647596
rect 674419 647531 674485 647532
rect 674974 647325 675034 651475
rect 675155 649772 675221 649773
rect 675155 649708 675156 649772
rect 675220 649708 675221 649772
rect 675155 649707 675221 649708
rect 675158 647597 675218 649707
rect 675155 647596 675221 647597
rect 675155 647532 675156 647596
rect 675220 647532 675221 647596
rect 675155 647531 675221 647532
rect 674971 647324 675037 647325
rect 674971 647260 674972 647324
rect 675036 647260 675037 647324
rect 674971 647259 675037 647260
rect 674051 645148 674117 645149
rect 674051 645084 674052 645148
rect 674116 645084 674117 645148
rect 674051 645083 674117 645084
rect 671475 643516 671541 643517
rect 671475 643452 671476 643516
rect 671540 643452 671541 643516
rect 671475 643451 671541 643452
rect 41827 614140 41893 614141
rect 41827 614076 41828 614140
rect 41892 614076 41893 614140
rect 41827 614075 41893 614076
rect 44219 614140 44285 614141
rect 44219 614076 44220 614140
rect 44284 614076 44285 614140
rect 44219 614075 44285 614076
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 596460 41893 596461
rect 41827 596396 41828 596460
rect 41892 596396 41893 596460
rect 41827 596395 41893 596396
rect 41830 596050 41890 596395
rect 41646 595990 41890 596050
rect 40539 589660 40605 589661
rect 40539 589596 40540 589660
rect 40604 589596 40605 589660
rect 40539 589595 40605 589596
rect 40723 589660 40789 589661
rect 40723 589596 40724 589660
rect 40788 589596 40789 589660
rect 40723 589595 40789 589596
rect 40542 576877 40602 589595
rect 40726 578237 40786 589595
rect 40907 589388 40973 589389
rect 40907 589324 40908 589388
rect 40972 589324 40973 589388
rect 40907 589323 40973 589324
rect 40723 578236 40789 578237
rect 40723 578172 40724 578236
rect 40788 578172 40789 578236
rect 40723 578171 40789 578172
rect 40910 577557 40970 589323
rect 41646 589290 41706 595990
rect 41827 593196 41893 593197
rect 41827 593132 41828 593196
rect 41892 593132 41893 593196
rect 41827 593131 41893 593132
rect 41830 589661 41890 593131
rect 41827 589660 41893 589661
rect 41827 589596 41828 589660
rect 41892 589596 41893 589660
rect 41827 589595 41893 589596
rect 42014 589290 42074 597211
rect 42195 592380 42261 592381
rect 42195 592316 42196 592380
rect 42260 592316 42261 592380
rect 42195 592315 42261 592316
rect 42198 589389 42258 592315
rect 43851 591564 43917 591565
rect 43851 591500 43852 591564
rect 43916 591500 43917 591564
rect 43851 591499 43917 591500
rect 42195 589388 42261 589389
rect 42195 589324 42196 589388
rect 42260 589324 42261 589388
rect 42195 589323 42261 589324
rect 41462 589230 41706 589290
rect 41830 589230 42074 589290
rect 41091 584628 41157 584629
rect 41091 584564 41092 584628
rect 41156 584564 41157 584628
rect 41091 584563 41157 584564
rect 41094 580277 41154 584563
rect 41091 580276 41157 580277
rect 41091 580212 41092 580276
rect 41156 580212 41157 580276
rect 41091 580211 41157 580212
rect 40907 577556 40973 577557
rect 40907 577492 40908 577556
rect 40972 577492 40973 577556
rect 40907 577491 40973 577492
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 571981 41522 589230
rect 41830 587210 41890 589230
rect 41646 587150 41890 587210
rect 41459 571980 41525 571981
rect 41459 571916 41460 571980
rect 41524 571916 41525 571980
rect 41459 571915 41525 571916
rect 41646 571029 41706 587150
rect 42011 585444 42077 585445
rect 42011 585380 42012 585444
rect 42076 585380 42077 585444
rect 42011 585379 42077 585380
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41830 572253 41890 585107
rect 42014 580549 42074 585379
rect 42011 580548 42077 580549
rect 42011 580484 42012 580548
rect 42076 580484 42077 580548
rect 42011 580483 42077 580484
rect 42379 577420 42445 577421
rect 42379 577356 42380 577420
rect 42444 577356 42445 577420
rect 42379 577355 42445 577356
rect 42382 572661 42442 577355
rect 42379 572660 42445 572661
rect 42379 572596 42380 572660
rect 42444 572596 42445 572660
rect 42379 572595 42445 572596
rect 41827 572252 41893 572253
rect 41827 572188 41828 572252
rect 41892 572188 41893 572252
rect 41827 572187 41893 572188
rect 41643 571028 41709 571029
rect 41643 570964 41644 571028
rect 41708 570964 41709 571028
rect 41643 570963 41709 570964
rect 42011 553076 42077 553077
rect 42011 553012 42012 553076
rect 42076 553012 42077 553076
rect 42011 553011 42077 553012
rect 42014 549130 42074 553011
rect 42195 551852 42261 551853
rect 42195 551788 42196 551852
rect 42260 551788 42261 551852
rect 42195 551787 42261 551788
rect 41462 549070 42074 549130
rect 40539 545732 40605 545733
rect 40539 545668 40540 545732
rect 40604 545668 40605 545732
rect 40539 545667 40605 545668
rect 40542 537029 40602 545667
rect 40723 545460 40789 545461
rect 40723 545396 40724 545460
rect 40788 545396 40789 545460
rect 40723 545395 40789 545396
rect 40539 537028 40605 537029
rect 40539 536964 40540 537028
rect 40604 536964 40605 537028
rect 40539 536963 40605 536964
rect 40726 535261 40786 545395
rect 40723 535260 40789 535261
rect 40723 535196 40724 535260
rect 40788 535196 40789 535260
rect 40723 535195 40789 535196
rect 41462 530637 41522 549070
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 530636 41525 530637
rect 41459 530572 41460 530636
rect 41524 530572 41525 530636
rect 41459 530571 41525 530572
rect 41646 529141 41706 546347
rect 42198 543750 42258 551787
rect 41830 543690 42258 543750
rect 41830 529413 41890 543690
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 41643 529140 41709 529141
rect 41643 529076 41644 529140
rect 41708 529076 41709 529140
rect 41643 529075 41709 529076
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41646 424630 41890 424690
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40723 418572 40789 418573
rect 40723 418508 40724 418572
rect 40788 418508 40789 418572
rect 40723 418507 40789 418508
rect 40539 418300 40605 418301
rect 40539 418236 40540 418300
rect 40604 418236 40605 418300
rect 40539 418235 40605 418236
rect 40542 403885 40602 418235
rect 40726 409461 40786 418507
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 398853 41522 418779
rect 41646 402990 41706 424630
rect 42014 415410 42074 424763
rect 41830 415350 42074 415410
rect 41830 406333 41890 415350
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401845 41890 402930
rect 41827 401844 41893 401845
rect 41827 401780 41828 401844
rect 41892 401780 41893 401844
rect 41827 401779 41893 401780
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363629 40786 378115
rect 41275 373284 41341 373285
rect 41275 373220 41276 373284
rect 41340 373220 41341 373284
rect 41275 373219 41341 373220
rect 41278 368525 41338 373219
rect 41275 368524 41341 368525
rect 41275 368460 41276 368524
rect 41340 368460 41341 368524
rect 41275 368459 41341 368460
rect 40723 363628 40789 363629
rect 40723 363564 40724 363628
rect 40788 363564 40789 363628
rect 40723 363563 40789 363564
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 358733 41522 381787
rect 41643 376956 41709 376957
rect 41643 376892 41644 376956
rect 41708 376892 41709 376956
rect 41643 376891 41709 376892
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 41646 358050 41706 376891
rect 41827 371924 41893 371925
rect 41827 371860 41828 371924
rect 41892 371860 41893 371924
rect 41827 371859 41893 371860
rect 41830 359413 41890 371859
rect 41827 359412 41893 359413
rect 41827 359348 41828 359412
rect 41892 359348 41893 359412
rect 41827 359347 41893 359348
rect 41646 357990 41890 358050
rect 41830 355741 41890 357990
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43854 354245 43914 591499
rect 671478 571165 671538 643451
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 671475 571164 671541 571165
rect 671475 571100 671476 571164
rect 671540 571100 671541 571164
rect 671475 571099 671541 571100
rect 673683 475420 673749 475421
rect 673683 475356 673684 475420
rect 673748 475356 673749 475420
rect 673683 475355 673749 475356
rect 673686 464813 673746 475355
rect 673683 464812 673749 464813
rect 673683 464748 673684 464812
rect 673748 464748 673749 464812
rect 673683 464747 673749 464748
rect 673870 455157 673930 616115
rect 674054 475421 674114 645083
rect 675155 644060 675221 644061
rect 675155 643996 675156 644060
rect 675220 643996 675221 644060
rect 675155 643995 675221 643996
rect 675158 638077 675218 643995
rect 675155 638076 675221 638077
rect 675155 638012 675156 638076
rect 675220 638012 675221 638076
rect 675155 638011 675221 638012
rect 675342 637669 675402 652835
rect 676811 644332 676877 644333
rect 676811 644268 676812 644332
rect 676876 644268 676877 644332
rect 676811 644267 676877 644268
rect 676627 640252 676693 640253
rect 676627 640188 676628 640252
rect 676692 640188 676693 640252
rect 676627 640187 676693 640188
rect 676630 637941 676690 640187
rect 676627 637940 676693 637941
rect 676627 637876 676628 637940
rect 676692 637876 676693 637940
rect 676627 637875 676693 637876
rect 675339 637668 675405 637669
rect 675339 637604 675340 637668
rect 675404 637604 675405 637668
rect 675339 637603 675405 637604
rect 675339 631412 675405 631413
rect 675339 631348 675340 631412
rect 675404 631348 675405 631412
rect 675339 631347 675405 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674422 527101 674482 602923
rect 675342 592381 675402 631347
rect 675523 607748 675589 607749
rect 675523 607684 675524 607748
rect 675588 607684 675589 607748
rect 675523 607683 675589 607684
rect 675339 592380 675405 592381
rect 675339 592316 675340 592380
rect 675404 592316 675405 592380
rect 675339 592315 675405 592316
rect 675526 592109 675586 607683
rect 676078 593469 676138 631347
rect 676075 593468 676141 593469
rect 676075 593404 676076 593468
rect 676140 593404 676141 593468
rect 676075 593403 676141 593404
rect 675523 592108 675589 592109
rect 675523 592044 675524 592108
rect 675588 592044 675589 592108
rect 675523 592043 675589 592044
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 563140 675405 563141
rect 675339 563076 675340 563140
rect 675404 563076 675405 563140
rect 675339 563075 675405 563076
rect 675342 546005 675402 563075
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 675526 546549 675586 561171
rect 676078 546549 676138 586195
rect 676814 572797 676874 644267
rect 676998 619173 677058 694043
rect 676995 619172 677061 619173
rect 676995 619108 676996 619172
rect 677060 619108 677061 619172
rect 676995 619107 677061 619108
rect 676995 593468 677061 593469
rect 676995 593404 676996 593468
rect 677060 593404 677061 593468
rect 676995 593403 677061 593404
rect 676998 576061 677058 593403
rect 676995 576060 677061 576061
rect 676995 575996 676996 576060
rect 677060 575996 677061 576060
rect 676995 575995 677061 575996
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 676811 557564 676877 557565
rect 676811 557500 676812 557564
rect 676876 557500 676877 557564
rect 676811 557499 676877 557500
rect 675523 546548 675589 546549
rect 675523 546484 675524 546548
rect 675588 546484 675589 546548
rect 675523 546483 675589 546484
rect 676075 546548 676141 546549
rect 676075 546484 676076 546548
rect 676140 546484 676141 546548
rect 676075 546483 676141 546484
rect 675339 546004 675405 546005
rect 675339 545940 675340 546004
rect 675404 545940 675405 546004
rect 675339 545939 675405 545940
rect 674419 527100 674485 527101
rect 674419 527036 674420 527100
rect 674484 527036 674485 527100
rect 674419 527035 674485 527036
rect 676814 503709 676874 557499
rect 677179 550764 677245 550765
rect 677179 550700 677180 550764
rect 677244 550700 677245 550764
rect 677179 550699 677245 550700
rect 676811 503708 676877 503709
rect 676811 503644 676812 503708
rect 676876 503644 676877 503708
rect 676811 503643 676877 503644
rect 677182 495450 677242 550699
rect 677182 495390 677426 495450
rect 677366 492421 677426 495390
rect 677363 492420 677429 492421
rect 677363 492356 677364 492420
rect 677428 492356 677429 492420
rect 677363 492355 677429 492356
rect 675891 490516 675957 490517
rect 675891 490452 675892 490516
rect 675956 490452 675957 490516
rect 675891 490451 675957 490452
rect 675894 489970 675954 490451
rect 675894 489910 677058 489970
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 675894 488610 675954 488819
rect 675894 488550 676874 488610
rect 674051 475420 674117 475421
rect 674051 475356 674052 475420
rect 674116 475356 674117 475420
rect 674051 475355 674117 475356
rect 673867 455156 673933 455157
rect 673867 455092 673868 455156
rect 673932 455092 673933 455156
rect 673867 455091 673933 455092
rect 676814 401301 676874 488550
rect 676998 402933 677058 489910
rect 676995 402932 677061 402933
rect 676995 402868 676996 402932
rect 677060 402868 677061 402932
rect 676995 402867 677061 402868
rect 676811 401300 676877 401301
rect 676811 401236 676812 401300
rect 676876 401236 676877 401300
rect 676811 401235 676877 401236
rect 675891 398852 675957 398853
rect 675891 398788 675892 398852
rect 675956 398788 675957 398852
rect 675891 398787 675957 398788
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 674790 372605 674850 377979
rect 675894 377501 675954 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676075 393140 676141 393141
rect 676075 393076 676076 393140
rect 676140 393076 676141 393140
rect 676075 393075 676141 393076
rect 675891 377500 675957 377501
rect 675891 377436 675892 377500
rect 675956 377436 675957 377500
rect 675891 377435 675957 377436
rect 676078 373013 676138 393075
rect 676262 384981 676322 396747
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676259 384980 676325 384981
rect 676259 384916 676260 384980
rect 676324 384916 676325 384980
rect 676259 384915 676325 384916
rect 676446 380629 676506 394707
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676630 377229 676690 395115
rect 676627 377228 676693 377229
rect 676627 377164 676628 377228
rect 676692 377164 676693 377228
rect 676627 377163 676693 377164
rect 676075 373012 676141 373013
rect 676075 372948 676076 373012
rect 676140 372948 676141 373012
rect 676075 372947 676141 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 43851 354244 43917 354245
rect 43851 354180 43852 354244
rect 43916 354180 43917 354244
rect 43851 354179 43917 354180
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 44219 353836 44285 353837
rect 44219 353772 44220 353836
rect 44284 353772 44285 353836
rect 44219 353771 44285 353772
rect 44222 342549 44282 353771
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 342548 44285 342549
rect 44219 342484 44220 342548
rect 44284 342484 44285 342548
rect 44219 342483 44285 342484
rect 44406 341730 44466 342891
rect 44587 342140 44653 342141
rect 44587 342076 44588 342140
rect 44652 342076 44653 342140
rect 44587 342075 44653 342076
rect 44222 341670 44466 341730
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 40723 337788 40789 337789
rect 40723 337724 40724 337788
rect 40788 337724 40789 337788
rect 40723 337723 40789 337724
rect 40539 335748 40605 335749
rect 40539 335684 40540 335748
rect 40604 335684 40605 335748
rect 40539 335683 40605 335684
rect 40542 321197 40602 335683
rect 40726 326773 40786 337723
rect 42747 337652 42813 337653
rect 42747 337588 42748 337652
rect 42812 337588 42813 337652
rect 42747 337587 42813 337588
rect 42563 335476 42629 335477
rect 42563 335412 42564 335476
rect 42628 335412 42629 335476
rect 42563 335411 42629 335412
rect 41278 335341 41522 335370
rect 41275 335340 41522 335341
rect 41275 335276 41276 335340
rect 41340 335310 41522 335340
rect 41340 335276 41341 335310
rect 41275 335275 41341 335276
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40723 326772 40789 326773
rect 40723 326708 40724 326772
rect 40788 326708 40789 326772
rect 40723 326707 40789 326708
rect 40910 325413 40970 333643
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41462 324733 41522 335310
rect 42566 334661 42626 335411
rect 42563 334660 42629 334661
rect 42563 334596 42564 334660
rect 42628 334596 42629 334660
rect 42563 334595 42629 334596
rect 41643 329084 41709 329085
rect 41643 329020 41644 329084
rect 41708 329020 41709 329084
rect 41643 329019 41709 329020
rect 41459 324732 41525 324733
rect 41459 324668 41460 324732
rect 41524 324668 41525 324732
rect 41459 324667 41525 324668
rect 40539 321196 40605 321197
rect 40539 321132 40540 321196
rect 40604 321132 40605 321196
rect 40539 321131 40605 321132
rect 41646 315890 41706 329019
rect 42011 328404 42077 328405
rect 42011 328340 42012 328404
rect 42076 328340 42077 328404
rect 42011 328339 42077 328340
rect 41646 315830 41890 315890
rect 41830 315621 41890 315830
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 42014 312629 42074 328339
rect 42750 321570 42810 337587
rect 42931 336836 42997 336837
rect 42931 336772 42932 336836
rect 42996 336772 42997 336836
rect 42931 336771 42997 336772
rect 42934 331230 42994 336771
rect 43115 336156 43181 336157
rect 43115 336092 43116 336156
rect 43180 336092 43181 336156
rect 43115 336091 43181 336092
rect 43118 334661 43178 336091
rect 43115 334660 43181 334661
rect 43115 334596 43116 334660
rect 43180 334596 43181 334660
rect 43115 334595 43181 334596
rect 42934 331170 43178 331230
rect 42750 321510 42994 321570
rect 42934 312765 42994 321510
rect 43118 316437 43178 331170
rect 43115 316436 43181 316437
rect 43115 316372 43116 316436
rect 43180 316372 43181 316436
rect 43115 316371 43181 316372
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 42011 312628 42077 312629
rect 42011 312564 42012 312628
rect 42076 312564 42077 312628
rect 42011 312563 42077 312564
rect 43670 297669 43730 340443
rect 44222 311541 44282 341670
rect 44403 341324 44469 341325
rect 44403 341260 44404 341324
rect 44468 341260 44469 341324
rect 44403 341259 44469 341260
rect 44219 311540 44285 311541
rect 44219 311476 44220 311540
rect 44284 311476 44285 311540
rect 44219 311475 44285 311476
rect 44406 311269 44466 341259
rect 44403 311268 44469 311269
rect 44403 311204 44404 311268
rect 44468 311204 44469 311268
rect 44403 311203 44469 311204
rect 44590 311133 44650 342075
rect 675342 339013 675402 354179
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 350550 675770 352955
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 351250 675954 351731
rect 675894 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675526 350490 675770 350550
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675339 339012 675405 339013
rect 675339 338948 675340 339012
rect 675404 338948 675405 339012
rect 675339 338947 675405 338948
rect 675526 337789 675586 350490
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675891 349212 675957 349213
rect 675891 349148 675892 349212
rect 675956 349210 675957 349212
rect 675956 349150 676138 349210
rect 675956 349148 675957 349150
rect 675891 349147 675957 349148
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 676078 328405 676138 349150
rect 676262 332213 676322 349830
rect 676446 336701 676506 350510
rect 676630 340373 676690 351190
rect 676627 340372 676693 340373
rect 676627 340308 676628 340372
rect 676692 340308 676693 340372
rect 676627 340307 676693 340308
rect 676443 336700 676509 336701
rect 676443 336636 676444 336700
rect 676508 336636 676509 336700
rect 676443 336635 676509 336636
rect 676259 332212 676325 332213
rect 676259 332148 676260 332212
rect 676324 332148 676325 332212
rect 676259 332147 676325 332148
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 44587 311132 44653 311133
rect 44587 311068 44588 311132
rect 44652 311068 44653 311132
rect 44587 311067 44653 311068
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 303650 675770 308755
rect 675891 306780 675957 306781
rect 675891 306716 675892 306780
rect 675956 306716 675957 306780
rect 675891 306715 675957 306716
rect 675894 305010 675954 306715
rect 675894 304950 676322 305010
rect 675710 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 292770 41890 295563
rect 40726 292710 41890 292770
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 40726 278493 40786 292710
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 40907 292527 40973 292528
rect 40723 278492 40789 278493
rect 40723 278428 40724 278492
rect 40788 278428 40789 278492
rect 40723 278427 40789 278428
rect 40910 277949 40970 292527
rect 41827 292500 41893 292501
rect 41827 292436 41828 292500
rect 41892 292436 41893 292500
rect 41827 292435 41893 292436
rect 41830 292090 41890 292435
rect 41646 292030 41890 292090
rect 41646 289830 41706 292030
rect 41827 290460 41893 290461
rect 41827 290396 41828 290460
rect 41892 290396 41893 290460
rect 41827 290395 41893 290396
rect 41462 289770 41706 289830
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 289770
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 290395
rect 42014 281485 42074 296379
rect 675710 281621 675770 297331
rect 675894 282845 675954 302635
rect 676078 283661 676138 303590
rect 676262 295221 676322 304950
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676259 295220 676325 295221
rect 676259 295156 676260 295220
rect 676324 295156 676325 295220
rect 676259 295155 676325 295156
rect 676446 291549 676506 301547
rect 676627 301476 676693 301477
rect 676627 301412 676628 301476
rect 676692 301412 676693 301476
rect 676627 301411 676693 301412
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676630 287061 676690 301411
rect 676627 287060 676693 287061
rect 676627 286996 676628 287060
rect 676692 286996 676693 287060
rect 676627 286995 676693 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 674971 263668 675037 263669
rect 674971 263604 674972 263668
rect 675036 263604 675037 263668
rect 674971 263603 675037 263604
rect 674974 253950 675034 263603
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 674790 253890 675034 253950
rect 40723 251428 40789 251429
rect 40723 251364 40724 251428
rect 40788 251364 40789 251428
rect 40723 251363 40789 251364
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 235925 40602 249731
rect 40726 240141 40786 251363
rect 674790 249661 674850 253890
rect 676078 249661 676138 262379
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 676814 245309 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 245308 676877 245309
rect 676811 245244 676812 245308
rect 676876 245244 676877 245308
rect 676811 245243 676877 245244
rect 675155 245036 675221 245037
rect 675155 244972 675156 245036
rect 675220 244972 675221 245036
rect 675155 244971 675221 244972
rect 675158 240277 675218 244971
rect 675339 244764 675405 244765
rect 675339 244700 675340 244764
rect 675404 244700 675405 244764
rect 675339 244699 675405 244700
rect 675155 240276 675221 240277
rect 675155 240212 675156 240276
rect 675220 240212 675221 240276
rect 675155 240211 675221 240212
rect 40723 240140 40789 240141
rect 40723 240076 40724 240140
rect 40788 240076 40789 240140
rect 40723 240075 40789 240076
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40539 235924 40605 235925
rect 40539 235860 40540 235924
rect 40604 235860 40605 235924
rect 40539 235859 40605 235860
rect 42014 227357 42074 238035
rect 675342 236877 675402 244699
rect 675339 236876 675405 236877
rect 675339 236812 675340 236876
rect 675404 236812 675405 236876
rect 675339 236811 675405 236812
rect 674235 233204 674301 233205
rect 674235 233140 674236 233204
rect 674300 233140 674301 233204
rect 674235 233139 674301 233140
rect 673683 231436 673749 231437
rect 673683 231372 673684 231436
rect 673748 231372 673749 231436
rect 673683 231371 673749 231372
rect 673131 230348 673197 230349
rect 673131 230284 673132 230348
rect 673196 230284 673197 230348
rect 673131 230283 673197 230284
rect 673315 230348 673381 230349
rect 673315 230284 673316 230348
rect 673380 230284 673381 230348
rect 673315 230283 673381 230284
rect 667979 229804 668045 229805
rect 667979 229740 667980 229804
rect 668044 229740 668045 229804
rect 667979 229739 668045 229740
rect 668163 229804 668229 229805
rect 668163 229740 668164 229804
rect 668228 229740 668229 229804
rect 668163 229739 668229 229740
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 565675 222596 565741 222597
rect 565675 222532 565676 222596
rect 565740 222532 565741 222596
rect 565675 222531 565741 222532
rect 540099 220556 540165 220557
rect 540099 220492 540100 220556
rect 540164 220492 540165 220556
rect 540099 220491 540165 220492
rect 563651 220556 563717 220557
rect 563651 220492 563652 220556
rect 563716 220492 563717 220556
rect 563651 220491 563717 220492
rect 511027 220012 511093 220013
rect 511027 219948 511028 220012
rect 511092 219948 511093 220012
rect 511027 219947 511093 219948
rect 526483 220012 526549 220013
rect 526483 219948 526484 220012
rect 526548 219948 526549 220012
rect 526483 219947 526549 219948
rect 508267 217836 508333 217837
rect 508267 217772 508268 217836
rect 508332 217772 508333 217836
rect 508267 217771 508333 217772
rect 504403 217564 504469 217565
rect 504403 217500 504404 217564
rect 504468 217500 504469 217564
rect 504403 217499 504469 217500
rect 504406 216205 504466 217499
rect 508270 217021 508330 217771
rect 508267 217020 508333 217021
rect 508267 216956 508268 217020
rect 508332 216956 508333 217020
rect 508267 216955 508333 216956
rect 511030 216205 511090 219947
rect 519859 219740 519925 219741
rect 519859 219676 519860 219740
rect 519924 219676 519925 219740
rect 519859 219675 519925 219676
rect 522619 219740 522685 219741
rect 522619 219676 522620 219740
rect 522684 219676 522685 219740
rect 522619 219675 522685 219676
rect 519862 216477 519922 219675
rect 519307 216476 519373 216477
rect 519307 216412 519308 216476
rect 519372 216412 519373 216476
rect 519307 216411 519373 216412
rect 519859 216476 519925 216477
rect 519859 216412 519860 216476
rect 519924 216412 519925 216476
rect 519859 216411 519925 216412
rect 504403 216204 504469 216205
rect 504403 216140 504404 216204
rect 504468 216140 504469 216204
rect 504403 216139 504469 216140
rect 511027 216204 511093 216205
rect 511027 216140 511028 216204
rect 511092 216140 511093 216204
rect 511027 216139 511093 216140
rect 519310 215933 519370 216411
rect 519307 215932 519373 215933
rect 519307 215868 519308 215932
rect 519372 215868 519373 215932
rect 519307 215867 519373 215868
rect 522622 215661 522682 219675
rect 522619 215660 522685 215661
rect 522619 215596 522620 215660
rect 522684 215596 522685 215660
rect 522619 215595 522685 215596
rect 526486 215389 526546 219947
rect 538814 216550 539978 216610
rect 536051 215932 536117 215933
rect 536051 215868 536052 215932
rect 536116 215868 536117 215932
rect 536051 215867 536117 215868
rect 526483 215388 526549 215389
rect 526483 215324 526484 215388
rect 526548 215324 526549 215388
rect 526483 215323 526549 215324
rect 536054 215117 536114 215867
rect 538814 215525 538874 216550
rect 538811 215524 538877 215525
rect 538811 215460 538812 215524
rect 538876 215460 538877 215524
rect 538811 215459 538877 215460
rect 539179 215524 539245 215525
rect 539179 215460 539180 215524
rect 539244 215460 539245 215524
rect 539179 215459 539245 215460
rect 536051 215116 536117 215117
rect 536051 215052 536052 215116
rect 536116 215052 536117 215116
rect 536051 215051 536117 215052
rect 538995 215116 539061 215117
rect 538995 215052 538996 215116
rect 539060 215114 539061 215116
rect 539182 215114 539242 215459
rect 539918 215389 539978 216550
rect 539915 215388 539981 215389
rect 539915 215324 539916 215388
rect 539980 215324 539981 215388
rect 539915 215323 539981 215324
rect 540102 215117 540162 220491
rect 554083 220284 554149 220285
rect 554083 220220 554084 220284
rect 554148 220220 554149 220284
rect 554083 220219 554149 220220
rect 554086 219418 554146 220219
rect 562547 219740 562613 219741
rect 562547 219676 562548 219740
rect 562612 219676 562613 219740
rect 562547 219675 562613 219676
rect 562550 218650 562610 219675
rect 562915 218652 562981 218653
rect 562915 218650 562916 218652
rect 562550 218590 562916 218650
rect 562915 218588 562916 218590
rect 562980 218588 562981 218652
rect 562915 218587 562981 218588
rect 562182 218381 562242 218502
rect 562179 218380 562245 218381
rect 562179 218316 562180 218380
rect 562244 218316 562245 218380
rect 562179 218315 562245 218316
rect 562731 217772 562732 217822
rect 562796 217772 562797 217822
rect 562731 217771 562797 217772
rect 563099 217564 563165 217565
rect 563099 217500 563100 217564
rect 563164 217500 563165 217564
rect 563099 217499 563165 217500
rect 563102 217290 563162 217499
rect 563654 217290 563714 220491
rect 565678 218058 565738 222531
rect 572483 222052 572549 222053
rect 572483 221988 572484 222052
rect 572548 221988 572549 222052
rect 572483 221987 572549 221988
rect 572486 220693 572546 221987
rect 572483 220692 572549 220693
rect 572483 220628 572484 220692
rect 572548 220628 572549 220692
rect 572483 220627 572549 220628
rect 568619 219740 568685 219741
rect 568619 219676 568620 219740
rect 568684 219676 568685 219740
rect 568619 219675 568685 219676
rect 568622 218738 568682 219675
rect 572667 219196 572733 219197
rect 572667 219132 572668 219196
rect 572732 219132 572733 219196
rect 572667 219131 572733 219132
rect 572851 219196 572917 219197
rect 572851 219132 572852 219196
rect 572916 219132 572917 219196
rect 572851 219131 572917 219132
rect 572670 218650 572730 219131
rect 572854 218650 572914 219131
rect 572670 218590 572914 218650
rect 575062 218245 575122 219182
rect 575059 218244 575125 218245
rect 575059 218180 575060 218244
rect 575124 218180 575125 218244
rect 575059 218179 575125 218180
rect 565678 217429 565738 217822
rect 567699 217462 567765 217463
rect 565675 217428 565741 217429
rect 565675 217364 565676 217428
rect 565740 217364 565741 217428
rect 567699 217398 567700 217462
rect 567764 217398 567765 217462
rect 567699 217397 567765 217398
rect 565675 217363 565741 217364
rect 546726 217230 547890 217290
rect 563102 217230 563714 217290
rect 546726 215661 546786 217230
rect 546910 216550 547706 216610
rect 546723 215660 546789 215661
rect 546723 215596 546724 215660
rect 546788 215596 546789 215660
rect 546723 215595 546789 215596
rect 546910 215117 546970 216550
rect 547646 215661 547706 216550
rect 547830 215930 547890 217230
rect 564942 217094 566658 217154
rect 556478 216550 558930 216610
rect 547830 215870 548442 215930
rect 548382 215661 548442 215870
rect 556478 215661 556538 216550
rect 558870 215661 558930 216550
rect 564942 216477 565002 217094
rect 566598 216477 566658 217094
rect 564939 216476 565005 216477
rect 564939 216412 564940 216476
rect 565004 216412 565005 216476
rect 564939 216411 565005 216412
rect 566595 216476 566661 216477
rect 566595 216412 566596 216476
rect 566660 216412 566661 216476
rect 566595 216411 566661 216412
rect 566414 215870 567026 215930
rect 566414 215661 566474 215870
rect 547643 215660 547709 215661
rect 547643 215596 547644 215660
rect 547708 215596 547709 215660
rect 547643 215595 547709 215596
rect 548195 215660 548261 215661
rect 548195 215596 548196 215660
rect 548260 215596 548261 215660
rect 548195 215595 548261 215596
rect 548379 215660 548445 215661
rect 548379 215596 548380 215660
rect 548444 215596 548445 215660
rect 548379 215595 548445 215596
rect 556475 215660 556541 215661
rect 556475 215596 556476 215660
rect 556540 215596 556541 215660
rect 556475 215595 556541 215596
rect 558867 215660 558933 215661
rect 558867 215596 558868 215660
rect 558932 215596 558933 215660
rect 558867 215595 558933 215596
rect 566411 215660 566477 215661
rect 566411 215596 566412 215660
rect 566476 215596 566477 215660
rect 566411 215595 566477 215596
rect 548198 215117 548258 215595
rect 566966 215117 567026 215870
rect 539060 215054 539242 215114
rect 540099 215116 540165 215117
rect 539060 215052 539061 215054
rect 538995 215051 539061 215052
rect 540099 215052 540100 215116
rect 540164 215052 540165 215116
rect 540099 215051 540165 215052
rect 546907 215116 546973 215117
rect 546907 215052 546908 215116
rect 546972 215052 546973 215116
rect 546907 215051 546973 215052
rect 548195 215116 548261 215117
rect 548195 215052 548196 215116
rect 548260 215052 548261 215116
rect 548195 215051 548261 215052
rect 566963 215116 567029 215117
rect 566963 215052 566964 215116
rect 567028 215052 567029 215116
rect 567702 215114 567762 217397
rect 568438 216550 570154 216610
rect 567883 215388 567949 215389
rect 567883 215324 567884 215388
rect 567948 215386 567949 215388
rect 568438 215386 568498 216550
rect 570094 215930 570154 216550
rect 572851 215932 572917 215933
rect 572851 215930 572852 215932
rect 570094 215870 572852 215930
rect 572851 215868 572852 215870
rect 572916 215868 572917 215932
rect 572851 215867 572917 215868
rect 572483 215660 572549 215661
rect 572483 215596 572484 215660
rect 572548 215596 572549 215660
rect 572483 215595 572549 215596
rect 567948 215326 568498 215386
rect 572486 215386 572546 215595
rect 572486 215326 573466 215386
rect 567948 215324 567949 215326
rect 567883 215323 567949 215324
rect 568251 215116 568317 215117
rect 568251 215114 568252 215116
rect 567702 215054 568252 215114
rect 566963 215051 567029 215052
rect 568251 215052 568252 215054
rect 568316 215052 568317 215116
rect 568251 215051 568317 215052
rect 573406 214658 573466 215326
rect 575614 214981 575674 217142
rect 583710 215933 583770 217822
rect 583707 215932 583773 215933
rect 583707 215868 583708 215932
rect 583772 215868 583773 215932
rect 583707 215867 583773 215868
rect 576715 215388 576781 215389
rect 576715 215324 576716 215388
rect 576780 215324 576781 215388
rect 576715 215323 576781 215324
rect 575611 214980 575677 214981
rect 575611 214916 575612 214980
rect 575676 214916 575677 214980
rect 575611 214915 575677 214916
rect 576718 214658 576778 215323
rect 41459 209812 41525 209813
rect 41459 209748 41460 209812
rect 41524 209748 41525 209812
rect 41459 209747 41525 209748
rect 40723 208180 40789 208181
rect 40723 208116 40724 208180
rect 40788 208116 40789 208180
rect 40723 208115 40789 208116
rect 40539 206956 40605 206957
rect 40539 206892 40540 206956
rect 40604 206892 40605 206956
rect 40539 206891 40605 206892
rect 40542 194581 40602 206891
rect 40726 197165 40786 208115
rect 40907 207364 40973 207365
rect 40907 207300 40908 207364
rect 40972 207300 40973 207364
rect 40907 207299 40973 207300
rect 40723 197164 40789 197165
rect 40723 197100 40724 197164
rect 40788 197100 40789 197164
rect 40723 197099 40789 197100
rect 40910 195533 40970 207299
rect 40907 195532 40973 195533
rect 40907 195468 40908 195532
rect 40972 195468 40973 195532
rect 40907 195467 40973 195468
rect 41462 195261 41522 209747
rect 42011 207772 42077 207773
rect 42011 207708 42012 207772
rect 42076 207708 42077 207772
rect 42011 207707 42077 207708
rect 41827 197844 41893 197845
rect 41827 197780 41828 197844
rect 41892 197780 41893 197844
rect 41827 197779 41893 197780
rect 41830 195805 41890 197779
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 41459 195260 41525 195261
rect 41459 195196 41460 195260
rect 41524 195196 41525 195260
rect 41459 195195 41525 195196
rect 40539 194580 40605 194581
rect 40539 194516 40540 194580
rect 40604 194516 40605 194580
rect 40539 194515 40605 194516
rect 41643 194580 41709 194581
rect 41643 194516 41644 194580
rect 41708 194516 41709 194580
rect 41643 194515 41709 194516
rect 41646 190470 41706 194515
rect 41646 190410 41890 190470
rect 41830 187237 41890 190410
rect 41827 187236 41893 187237
rect 41827 187172 41828 187236
rect 41892 187172 41893 187236
rect 41827 187171 41893 187172
rect 42014 185877 42074 207707
rect 42379 192948 42445 192949
rect 42379 192884 42380 192948
rect 42444 192884 42445 192948
rect 42379 192883 42445 192884
rect 42382 186149 42442 192883
rect 42379 186148 42445 186149
rect 42379 186084 42380 186148
rect 42444 186084 42445 186148
rect 42379 186083 42445 186084
rect 42011 185876 42077 185877
rect 42011 185812 42012 185876
rect 42076 185812 42077 185876
rect 42011 185811 42077 185812
rect 667982 130525 668042 229739
rect 668166 229261 668226 229739
rect 668163 229260 668229 229261
rect 668163 229196 668164 229260
rect 668228 229196 668229 229260
rect 668163 229195 668229 229196
rect 672947 228716 673013 228717
rect 672947 228652 672948 228716
rect 673012 228652 673013 228716
rect 672947 228651 673013 228652
rect 671107 227220 671173 227221
rect 671107 227156 671108 227220
rect 671172 227156 671173 227220
rect 671107 227155 671173 227156
rect 671110 224093 671170 227155
rect 672027 226676 672093 226677
rect 672027 226612 672028 226676
rect 672092 226612 672093 226676
rect 672027 226611 672093 226612
rect 671659 226404 671725 226405
rect 671659 226340 671660 226404
rect 671724 226340 671725 226404
rect 671659 226339 671725 226340
rect 671662 225045 671722 226339
rect 672030 226133 672090 226611
rect 672027 226132 672093 226133
rect 672027 226068 672028 226132
rect 672092 226068 672093 226132
rect 672027 226067 672093 226068
rect 671659 225044 671725 225045
rect 671659 224980 671660 225044
rect 671724 224980 671725 225044
rect 671659 224979 671725 224980
rect 671107 224092 671173 224093
rect 671107 224028 671108 224092
rect 671172 224028 671173 224092
rect 671107 224027 671173 224028
rect 672027 221100 672093 221101
rect 672027 221036 672028 221100
rect 672092 221036 672093 221100
rect 672027 221035 672093 221036
rect 670739 220964 670805 220965
rect 670739 220900 670740 220964
rect 670804 220900 670805 220964
rect 670739 220899 670805 220900
rect 669451 211172 669517 211173
rect 669451 211108 669452 211172
rect 669516 211108 669517 211172
rect 669451 211107 669517 211108
rect 669454 195990 669514 211107
rect 669270 195930 669514 195990
rect 669270 176670 669330 195930
rect 669270 176610 669514 176670
rect 669454 147690 669514 176610
rect 669270 147630 669514 147690
rect 669270 143581 669330 147630
rect 669267 143580 669333 143581
rect 669267 143516 669268 143580
rect 669332 143516 669333 143580
rect 669267 143515 669333 143516
rect 670742 133789 670802 220899
rect 672030 219877 672090 221035
rect 672027 219876 672093 219877
rect 672027 219812 672028 219876
rect 672092 219812 672093 219876
rect 672027 219811 672093 219812
rect 672950 183565 673010 228651
rect 673134 224365 673194 230283
rect 673131 224364 673197 224365
rect 673131 224300 673132 224364
rect 673196 224300 673197 224364
rect 673131 224299 673197 224300
rect 673318 224093 673378 230283
rect 673499 226540 673565 226541
rect 673499 226476 673500 226540
rect 673564 226476 673565 226540
rect 673499 226475 673565 226476
rect 673502 224909 673562 226475
rect 673686 225181 673746 231371
rect 673683 225180 673749 225181
rect 673683 225116 673684 225180
rect 673748 225116 673749 225180
rect 673683 225115 673749 225116
rect 673499 224908 673565 224909
rect 673499 224844 673500 224908
rect 673564 224844 673565 224908
rect 673499 224843 673565 224844
rect 673315 224092 673381 224093
rect 673315 224028 673316 224092
rect 673380 224028 673381 224092
rect 673315 224027 673381 224028
rect 673499 223684 673565 223685
rect 673499 223620 673500 223684
rect 673564 223620 673565 223684
rect 673499 223619 673565 223620
rect 673131 214708 673197 214709
rect 673131 214644 673132 214708
rect 673196 214644 673197 214708
rect 673131 214643 673197 214644
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 673134 164253 673194 214643
rect 673131 164252 673197 164253
rect 673131 164188 673132 164252
rect 673196 164188 673197 164252
rect 673131 164187 673197 164188
rect 670739 133788 670805 133789
rect 670739 133724 670740 133788
rect 670804 133724 670805 133788
rect 670739 133723 670805 133724
rect 667979 130524 668045 130525
rect 667979 130460 667980 130524
rect 668044 130460 668045 130524
rect 667979 130459 668045 130460
rect 673502 128893 673562 223619
rect 674051 212124 674117 212125
rect 674051 212060 674052 212124
rect 674116 212060 674117 212124
rect 674051 212059 674117 212060
rect 673499 128892 673565 128893
rect 673499 128828 673500 128892
rect 673564 128828 673565 128892
rect 673499 128827 673565 128828
rect 674054 128349 674114 212059
rect 674238 154597 674298 233139
rect 675155 228580 675221 228581
rect 675155 228516 675156 228580
rect 675220 228516 675221 228580
rect 675155 228515 675221 228516
rect 674971 218652 675037 218653
rect 674971 218588 674972 218652
rect 675036 218588 675037 218652
rect 674971 218587 675037 218588
rect 674974 210493 675034 218587
rect 675158 217293 675218 228515
rect 675339 226812 675405 226813
rect 675339 226748 675340 226812
rect 675404 226748 675405 226812
rect 675339 226747 675405 226748
rect 675155 217292 675221 217293
rect 675155 217228 675156 217292
rect 675220 217228 675221 217292
rect 675155 217227 675221 217228
rect 675342 216885 675402 226747
rect 675523 220012 675589 220013
rect 675523 219948 675524 220012
rect 675588 219948 675589 220012
rect 675523 219947 675589 219948
rect 675526 218925 675586 219947
rect 675523 218924 675589 218925
rect 675523 218860 675524 218924
rect 675588 218860 675589 218924
rect 675523 218859 675589 218860
rect 675891 218244 675957 218245
rect 675891 218180 675892 218244
rect 675956 218180 675957 218244
rect 675891 218179 675957 218180
rect 675523 217428 675589 217429
rect 675523 217364 675524 217428
rect 675588 217364 675589 217428
rect 675523 217363 675589 217364
rect 675339 216884 675405 216885
rect 675339 216820 675340 216884
rect 675404 216820 675405 216884
rect 675339 216819 675405 216820
rect 674971 210492 675037 210493
rect 674971 210428 674972 210492
rect 675036 210428 675037 210492
rect 674971 210427 675037 210428
rect 675526 198253 675586 217363
rect 675707 217020 675773 217021
rect 675707 216956 675708 217020
rect 675772 216956 675773 217020
rect 675707 216955 675773 216956
rect 675710 211170 675770 216955
rect 675894 215310 675954 218179
rect 675894 215250 676690 215310
rect 676075 215150 676141 215151
rect 676075 215086 676076 215150
rect 676140 215086 676141 215150
rect 676075 215085 676141 215086
rect 675891 214572 675957 214573
rect 675891 214508 675892 214572
rect 675956 214508 675957 214572
rect 675891 214507 675957 214508
rect 675894 211445 675954 214507
rect 676078 213890 676138 215085
rect 676078 213830 676322 213890
rect 675891 211444 675957 211445
rect 675891 211380 675892 211444
rect 675956 211380 675957 211444
rect 675891 211379 675957 211380
rect 675710 211110 676138 211170
rect 675891 210492 675957 210493
rect 675891 210428 675892 210492
rect 675956 210428 675957 210492
rect 675891 210427 675957 210428
rect 675523 198252 675589 198253
rect 675523 198188 675524 198252
rect 675588 198188 675589 198252
rect 675523 198187 675589 198188
rect 675894 193221 675954 210427
rect 675891 193220 675957 193221
rect 675891 193156 675892 193220
rect 675956 193156 675957 193220
rect 675891 193155 675957 193156
rect 676078 191589 676138 211110
rect 676262 197165 676322 213830
rect 676443 211444 676509 211445
rect 676443 211380 676444 211444
rect 676508 211380 676509 211444
rect 676443 211379 676509 211380
rect 676446 200701 676506 211379
rect 676630 205597 676690 215250
rect 676627 205596 676693 205597
rect 676627 205532 676628 205596
rect 676692 205532 676693 205596
rect 676627 205531 676693 205532
rect 676443 200700 676509 200701
rect 676443 200636 676444 200700
rect 676508 200636 676509 200700
rect 676443 200635 676509 200636
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675523 167516 675589 167517
rect 675523 167452 675524 167516
rect 675588 167452 675589 167516
rect 675523 167451 675589 167452
rect 675339 161940 675405 161941
rect 675339 161876 675340 161940
rect 675404 161876 675405 161940
rect 675339 161875 675405 161876
rect 675342 157045 675402 161875
rect 675526 157350 675586 167451
rect 675710 162210 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675891 172004 675957 172005
rect 675891 171940 675892 172004
rect 675956 171940 675957 172004
rect 675891 171939 675957 171940
rect 675894 167010 675954 171939
rect 675894 166950 676138 167010
rect 675710 162150 675954 162210
rect 675526 157290 675770 157350
rect 675339 157044 675405 157045
rect 675339 156980 675340 157044
rect 675404 156980 675405 157044
rect 675339 156979 675405 156980
rect 674235 154596 674301 154597
rect 674235 154532 674236 154596
rect 674300 154532 674301 154596
rect 674235 154531 674301 154532
rect 675710 147661 675770 157290
rect 675894 148477 675954 162150
rect 675891 148476 675957 148477
rect 675891 148412 675892 148476
rect 675956 148412 675957 148476
rect 675891 148411 675957 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 676078 146029 676138 166950
rect 676262 153101 676322 172350
rect 676446 159357 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159356 676509 159357
rect 676443 159292 676444 159356
rect 676508 159292 676509 159356
rect 676443 159291 676509 159292
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 153100 676325 153101
rect 676259 153036 676260 153100
rect 676324 153036 676325 153100
rect 676259 153035 676325 153036
rect 676075 146028 676141 146029
rect 676075 145964 676076 146028
rect 676140 145964 676141 146028
rect 676075 145963 676141 145964
rect 676627 128620 676693 128621
rect 676627 128556 676628 128620
rect 676692 128556 676693 128620
rect 676627 128555 676693 128556
rect 674051 128348 674117 128349
rect 674051 128284 674052 128348
rect 674116 128284 674117 128348
rect 674051 128283 674117 128284
rect 676075 128212 676141 128213
rect 676075 128148 676076 128212
rect 676140 128148 676141 128212
rect 676075 128147 676141 128148
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 122364 675773 122365
rect 675707 122300 675708 122364
rect 675772 122300 675773 122364
rect 675707 122299 675773 122300
rect 675710 102645 675770 122299
rect 675894 108085 675954 127195
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 128147
rect 676259 126988 676325 126989
rect 676259 126924 676260 126988
rect 676324 126924 676325 126988
rect 676259 126923 676325 126924
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676262 101421 676322 126923
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 106181 676506 124475
rect 676630 113117 676690 128555
rect 676627 113116 676693 113117
rect 676627 113052 676628 113116
rect 676692 113052 676693 113116
rect 676627 113051 676693 113052
rect 676443 106180 676509 106181
rect 676443 106116 676444 106180
rect 676508 106116 676509 106180
rect 676443 106115 676509 106116
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 634859 96660 634925 96661
rect 634859 96596 634860 96660
rect 634924 96596 634925 96660
rect 634859 96595 634925 96596
rect 637251 96660 637317 96661
rect 637251 96596 637252 96660
rect 637316 96596 637317 96660
rect 637251 96595 637317 96596
rect 634862 80477 634922 96595
rect 637254 84210 637314 96595
rect 637070 84150 637314 84210
rect 634859 80476 634925 80477
rect 634859 80412 634860 80476
rect 634924 80412 634925 80476
rect 634859 80411 634925 80412
rect 637070 77893 637130 84150
rect 637067 77892 637133 77893
rect 637067 77828 637068 77892
rect 637132 77828 637133 77892
rect 637067 77827 637133 77828
rect 461715 55044 461781 55045
rect 461715 54980 461716 55044
rect 461780 54980 461781 55044
rect 461715 54979 461781 54980
rect 461718 53957 461778 54979
rect 462635 54500 462701 54501
rect 462635 54436 462636 54500
rect 462700 54436 462701 54500
rect 462635 54435 462701 54436
rect 462638 53957 462698 54435
rect 461715 53956 461781 53957
rect 461715 53892 461716 53956
rect 461780 53892 461781 53956
rect 461715 53891 461781 53892
rect 462635 53956 462701 53957
rect 462635 53892 462636 53956
rect 462700 53892 462701 53956
rect 462635 53891 462701 53892
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40493 141802 43963
rect 194366 42125 194426 50219
rect 308995 49740 309061 49741
rect 308995 49676 308996 49740
rect 309060 49676 309061 49740
rect 308995 49675 309061 49676
rect 308998 42805 309058 49675
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47564 515509 47565
rect 515443 47500 515444 47564
rect 515508 47500 515509 47564
rect 515443 47499 515509 47500
rect 461347 44436 461413 44437
rect 461347 44372 461348 44436
rect 461412 44372 461413 44436
rect 461347 44371 461413 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 440187 43892 440253 43893
rect 440187 43828 440188 43892
rect 440252 43890 440253 43892
rect 440923 43892 440989 43893
rect 440923 43890 440924 43892
rect 440252 43830 440924 43890
rect 440252 43828 440253 43830
rect 440187 43827 440253 43828
rect 440923 43828 440924 43830
rect 440988 43828 440989 43892
rect 440923 43827 440989 43828
rect 308995 42804 309061 42805
rect 308995 42740 308996 42804
rect 309060 42740 309061 42804
rect 308995 42739 309061 42740
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 421974 41850 422034 42059
rect 461350 41938 461410 44371
rect 462270 41938 462330 44371
rect 515446 42125 515506 47499
rect 518758 42805 518818 48859
rect 526483 48108 526549 48109
rect 526483 48044 526484 48108
rect 526548 48044 526549 48108
rect 526483 48043 526549 48044
rect 520963 47836 521029 47837
rect 520963 47772 520964 47836
rect 521028 47772 521029 47836
rect 520963 47771 521029 47772
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47771
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 48043
rect 529798 42125 529858 50219
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 421974 41790 422162 41850
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 141739 40492 141805 40493
rect 141739 40428 141740 40492
rect 141804 40428 141805 40492
rect 141739 40427 141805 40428
<< via4 >>
rect 510942 997252 511178 997338
rect 510942 997188 511028 997252
rect 511028 997188 511092 997252
rect 511092 997188 511178 997252
rect 510942 997102 511178 997188
rect 522718 997102 522954 997338
rect 524006 997102 524242 997338
rect 531918 997102 532154 997338
rect 553446 997252 553682 997338
rect 553446 997188 553532 997252
rect 553532 997188 553596 997252
rect 553596 997188 553682 997252
rect 553446 997102 553682 997188
rect 636614 997102 636850 997338
rect 364110 993022 364346 993258
rect 392998 993022 393234 993258
rect 493462 217292 493698 217378
rect 493462 217228 493548 217292
rect 493548 217228 493612 217292
rect 493612 217228 493698 217292
rect 493462 217142 493698 217228
rect 553998 219182 554234 219418
rect 562094 218502 562330 218738
rect 562646 217836 562882 218058
rect 562646 217822 562732 217836
rect 562732 217822 562796 217836
rect 562796 217822 562882 217836
rect 563198 217972 563434 218058
rect 563198 217908 563284 217972
rect 563284 217908 563348 217972
rect 563348 217908 563434 217972
rect 563198 217822 563434 217908
rect 574974 219182 575210 219418
rect 568534 218502 568770 218738
rect 565590 217822 565826 218058
rect 583622 217822 583858 218058
rect 575526 217142 575762 217378
rect 573318 214422 573554 214658
rect 576630 214422 576866 214658
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 510900 997338 522996 997380
rect 510900 997102 510942 997338
rect 511178 997102 522718 997338
rect 522954 997102 522996 997338
rect 510900 997060 522996 997102
rect 523964 997338 532196 997380
rect 523964 997102 524006 997338
rect 524242 997102 531918 997338
rect 532154 997102 532196 997338
rect 523964 997060 532196 997102
rect 553404 997338 636892 997380
rect 553404 997102 553446 997338
rect 553682 997102 636614 997338
rect 636850 997102 636892 997338
rect 553404 997060 636892 997102
rect 364068 993258 393276 993300
rect 364068 993022 364110 993258
rect 364346 993022 392998 993258
rect 393234 993022 393276 993258
rect 364068 992980 393276 993022
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 553956 219418 575252 219460
rect 553956 219182 553998 219418
rect 554234 219182 574974 219418
rect 575210 219182 575252 219418
rect 553956 219140 575252 219182
rect 562052 218738 568812 218780
rect 562052 218502 562094 218738
rect 562330 218502 568534 218738
rect 568770 218502 568812 218738
rect 562052 218460 568812 218502
rect 562604 218058 563476 218100
rect 562604 217822 562646 218058
rect 562882 217822 563198 218058
rect 563434 217822 563476 218058
rect 562604 217780 563476 217822
rect 565548 218058 583900 218100
rect 565548 217822 565590 218058
rect 565826 217822 583622 218058
rect 583858 217822 583900 218058
rect 565548 217780 583900 217822
rect 493420 217378 575804 217420
rect 493420 217142 493462 217378
rect 493698 217142 575526 217378
rect 575762 217142 575804 217378
rect 493420 217100 575804 217142
rect 573276 214658 576908 214700
rect 573276 214422 573318 214658
rect 573554 214422 576630 214658
rect 576866 214422 576908 214658
rect 573276 214380 576908 214422
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use xres_buf  rstb_level
timestamp 1665972027
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use caravel_clocking  clock_ctrl
timestamp 1665972027
transform 1 0 626764 0 1 63284
box 136 70 20000 12000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1665972027
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1665972027
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1665972027
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1665972027
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1665972027
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use simple_por  por
timestamp 1665972027
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1665972027
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1665972027
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1665972027
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1665972027
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1665972027
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1665972027
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1665972027
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1665972027
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1665972027
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1665972027
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1665972027
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1665972027
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1665972027
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1665972027
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1665972027
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1665972027
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1665972027
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1665972027
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1665972027
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1665972027
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1665972027
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1665972027
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1665972027
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1665972027
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1665972027
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1665972027
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1665972027
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1665972027
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1665972027
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1665972027
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1665972027
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1665972027
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1665972027
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1665972027
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1665972027
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1665972027
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1665972027
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1665972027
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1665972027
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1665972027
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1665972027
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1665972027
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1665972027
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1665972027
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1665972027
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1665972027
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1665972027
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1665972027
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1665972027
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1665972027
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1665972027
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1665972027
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1665972027
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1665972027
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1665972027
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1665972027
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1665972027
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1665972027
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1665972027
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1665972027
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1665972027
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1665972027
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1665972027
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1665972027
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1665972027
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1665972027
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1665972027
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1665972027
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1665972027
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1665972027
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1665972027
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1665972027
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1665972027
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1665972027
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1665972027
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1665972027
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1665972027
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1665972027
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1665972027
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1665972027
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1665972027
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1665972027
transform 1 0 0 0 1 0
box 6022 33900 711814 1031696
use user_project_wrapper  mprj
timestamp 1665972027
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1665972027
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering  sigbuf
timestamp 1665972027
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal3 s 418245 997803 418551 997897 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal3 s 417057 997799 417363 997893 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
