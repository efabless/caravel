magic
tech sky130A
magscale 1 2
timestamp 1636038212
<< obsli1 >>
rect 920 2159 10551 11441
<< obsm1 >>
rect 920 2128 22434 11824
<< obsm2 >>
rect 1032 167 22430 13841
<< metal3 >>
rect 14000 13744 34000 13864
rect 14000 13472 34000 13592
rect 14000 13064 34000 13184
rect 14000 12792 34000 12912
rect 14000 12520 34000 12640
rect 14000 12112 34000 12232
rect 14000 11840 34000 11960
rect 14000 11432 34000 11552
rect 14000 11160 34000 11280
rect 14000 10888 34000 11008
rect 14000 10480 34000 10600
rect 14000 10208 34000 10328
rect 14000 9800 34000 9920
rect 14000 9528 34000 9648
rect 14000 9256 34000 9376
rect 14000 8848 34000 8968
rect 14000 8576 34000 8696
rect 14000 8168 34000 8288
rect 14000 7896 34000 8016
rect 14000 7624 34000 7744
rect 14000 7216 34000 7336
rect 14000 6944 34000 7064
rect 14000 6536 34000 6656
rect 14000 6264 34000 6384
rect 14000 5992 34000 6112
rect 14000 5584 34000 5704
rect 14000 5312 34000 5432
rect 14000 4904 34000 5024
rect 14000 4632 34000 4752
rect 14000 4360 34000 4480
rect 14000 3952 34000 4072
rect 14000 3680 34000 3800
rect 14000 3272 34000 3392
rect 14000 3000 34000 3120
rect 14000 2728 34000 2848
rect 14000 2320 34000 2440
rect 14000 2048 34000 2168
rect 14000 1640 34000 1760
rect 14000 1368 34000 1488
rect 14000 1096 34000 1216
rect 14000 688 34000 808
rect 14000 416 34000 536
rect 14000 144 34000 264
<< obsm3 >>
rect 1117 13392 13920 13562
rect 1117 13264 14000 13392
rect 1117 12440 13920 13264
rect 1117 12312 14000 12440
rect 1117 11760 13920 12312
rect 1117 11632 14000 11760
rect 1117 10808 13920 11632
rect 1117 10680 14000 10808
rect 1117 10128 13920 10680
rect 1117 10000 14000 10128
rect 1117 9176 13920 10000
rect 1117 9048 14000 9176
rect 1117 8496 13920 9048
rect 1117 8368 14000 8496
rect 1117 7544 13920 8368
rect 1117 7416 14000 7544
rect 1117 6864 13920 7416
rect 1117 6736 14000 6864
rect 1117 5912 13920 6736
rect 1117 5784 14000 5912
rect 1117 5232 13920 5784
rect 1117 5104 14000 5232
rect 1117 4280 13920 5104
rect 1117 4152 14000 4280
rect 1117 3600 13920 4152
rect 1117 3472 14000 3600
rect 1117 2648 13920 3472
rect 1117 2520 14000 2648
rect 1117 1968 13920 2520
rect 1117 1840 14000 1968
rect 1117 1016 13920 1840
rect 1117 888 14000 1016
rect 1117 443 13920 888
<< metal4 >>
rect -1620 -364 -1300 13964
rect -960 296 -640 13304
rect -300 956 20 12644
rect 360 1616 680 11984
rect 2560 956 2880 12644
rect 4110 956 4430 12644
rect 5660 956 5980 12644
rect 7210 956 7530 12644
rect 8760 956 9080 12644
rect 10084 1616 10404 11984
rect 10744 956 11064 12644
rect 11404 296 11724 13304
rect 12064 -364 12384 13964
<< obsm4 >>
rect 1256 2632 2276 5448
<< metal5 >>
rect -1620 13644 12384 13964
rect -960 12984 11724 13304
rect -300 12324 11064 12644
rect 360 11664 10404 11984
rect -300 10166 11064 10486
rect -1620 9516 12384 9836
rect -300 8616 11064 8936
rect -1620 7966 12384 8286
rect -300 7066 11064 7386
rect -1620 6416 12384 6736
rect -300 5516 11064 5836
rect -1620 4866 12384 5186
rect -300 3966 11064 4286
rect -1620 3316 12384 3636
rect -300 2416 11064 2736
rect 360 1616 10404 1936
rect -300 956 11064 1276
rect -960 296 11724 616
rect -1620 -364 12384 -44
<< labels >>
rlabel metal3 s 14000 144 34000 264 6 gpio_defaults[0]
port 1 nsew signal input
rlabel metal3 s 14000 3272 34000 3392 6 gpio_defaults[10]
port 2 nsew signal input
rlabel metal3 s 14000 3680 34000 3800 6 gpio_defaults[11]
port 3 nsew signal input
rlabel metal3 s 14000 3952 34000 4072 6 gpio_defaults[12]
port 4 nsew signal input
rlabel metal3 s 14000 416 34000 536 6 gpio_defaults[1]
port 5 nsew signal input
rlabel metal3 s 14000 688 34000 808 6 gpio_defaults[2]
port 6 nsew signal input
rlabel metal3 s 14000 1096 34000 1216 6 gpio_defaults[3]
port 7 nsew signal input
rlabel metal3 s 14000 1368 34000 1488 6 gpio_defaults[4]
port 8 nsew signal input
rlabel metal3 s 14000 1640 34000 1760 6 gpio_defaults[5]
port 9 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 gpio_defaults[6]
port 10 nsew signal input
rlabel metal3 s 14000 2320 34000 2440 6 gpio_defaults[7]
port 11 nsew signal input
rlabel metal3 s 14000 2728 34000 2848 6 gpio_defaults[8]
port 12 nsew signal input
rlabel metal3 s 14000 3000 34000 3120 6 gpio_defaults[9]
port 13 nsew signal input
rlabel metal3 s 14000 4904 34000 5024 6 mgmt_gpio_in
port 14 nsew signal output
rlabel metal3 s 14000 5312 34000 5432 6 mgmt_gpio_oeb
port 15 nsew signal input
rlabel metal3 s 14000 5584 34000 5704 6 mgmt_gpio_out
port 16 nsew signal input
rlabel metal3 s 14000 4632 34000 4752 6 one
port 17 nsew signal output
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_ana_en
port 18 nsew signal output
rlabel metal3 s 14000 6264 34000 6384 6 pad_gpio_ana_pol
port 19 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ana_sel
port 20 nsew signal output
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_dm[0]
port 21 nsew signal output
rlabel metal3 s 14000 7216 34000 7336 6 pad_gpio_dm[1]
port 22 nsew signal output
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_dm[2]
port 23 nsew signal output
rlabel metal3 s 14000 7896 34000 8016 6 pad_gpio_holdover
port 24 nsew signal output
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_ib_mode_sel
port 25 nsew signal output
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_in
port 26 nsew signal input
rlabel metal3 s 14000 8848 34000 8968 6 pad_gpio_inenb
port 27 nsew signal output
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_out
port 28 nsew signal output
rlabel metal3 s 14000 9528 34000 9648 6 pad_gpio_outenb
port 29 nsew signal output
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_slow_sel
port 30 nsew signal output
rlabel metal3 s 14000 10208 34000 10328 6 pad_gpio_vtrip_sel
port 31 nsew signal output
rlabel metal3 s 14000 10480 34000 10600 6 resetn
port 32 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 resetn_out
port 33 nsew signal output
rlabel metal3 s 14000 11160 34000 11280 6 serial_clock
port 34 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_clock_out
port 35 nsew signal output
rlabel metal3 s 14000 11840 34000 11960 6 serial_data_in
port 36 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 37 nsew signal output
rlabel metal3 s 14000 12520 34000 12640 6 serial_load
port 38 nsew signal input
rlabel metal3 s 14000 12792 34000 12912 6 serial_load_out
port 39 nsew signal output
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_in
port 40 nsew signal output
rlabel metal3 s 14000 13472 34000 13592 6 user_gpio_oeb
port 41 nsew signal input
rlabel metal3 s 14000 13744 34000 13864 6 user_gpio_out
port 42 nsew signal input
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 43 nsew power input
rlabel metal5 s -300 2416 11064 2736 6 vccd
port 43 nsew power input
rlabel metal5 s -300 5516 11064 5836 6 vccd
port 43 nsew power input
rlabel metal5 s -300 8616 11064 8936 6 vccd
port 43 nsew power input
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 43 nsew power input
rlabel metal4 s 360 1616 680 11984 6 vccd
port 43 nsew power input
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 43 nsew power input
rlabel metal4 s 2560 956 2880 12644 6 vccd
port 43 nsew power input
rlabel metal4 s 5660 956 5980 12644 6 vccd
port 43 nsew power input
rlabel metal4 s 8760 956 9080 12644 6 vccd
port 43 nsew power input
rlabel metal5 s -960 296 11724 616 6 vccd1
port 44 nsew power input
rlabel metal5 s -1620 3316 12384 3636 6 vccd1
port 44 nsew power input
rlabel metal5 s -1620 6416 12384 6736 6 vccd1
port 44 nsew power input
rlabel metal5 s -1620 9516 12384 9836 6 vccd1
port 44 nsew power input
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 44 nsew power input
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 44 nsew power input
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 44 nsew power input
rlabel metal5 s -300 956 11064 1276 6 vssd
port 45 nsew ground input
rlabel metal5 s -300 3966 11064 4286 6 vssd
port 45 nsew ground input
rlabel metal5 s -300 7066 11064 7386 6 vssd
port 45 nsew ground input
rlabel metal5 s -300 10166 11064 10486 6 vssd
port 45 nsew ground input
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 45 nsew ground input
rlabel metal4 s -300 956 20 12644 4 vssd
port 45 nsew ground input
rlabel metal4 s 4110 956 4430 12644 6 vssd
port 45 nsew ground input
rlabel metal4 s 7210 956 7530 12644 6 vssd
port 45 nsew ground input
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 45 nsew ground input
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 46 nsew ground input
rlabel metal5 s -1620 4866 12384 5186 6 vssd1
port 46 nsew ground input
rlabel metal5 s -1620 7966 12384 8286 6 vssd1
port 46 nsew ground input
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 46 nsew ground input
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 46 nsew ground input
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 46 nsew ground input
rlabel metal3 s 14000 4360 34000 4480 6 zero
port 47 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 34000 14000
string LEFview TRUE
string GDS_FILE ../gds/gpio_control_block.gds
string GDS_END 601568
string GDS_START 153642
<< end >>

