module copyright_block_a ();
endmodule
