* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _386_/Y _460_/Q _432_/S VGND VGND VPWR VPWR _432_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_363_ _363_/A _363_/B VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__nor2_1
Xrebuffer7 _455_/Q VGND VGND VPWR VPWR _361_/C sky130_fd_sc_hd__clkbuf_2
X_294_ _296_/A _476_/Q _329_/B VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_415_ _366_/Y _455_/Q _417_/S VGND VGND VPWR VPWR _415_/X sky130_fd_sc_hd__mux2_1
X_277_ _434_/S _278_/B _278_/C VGND VGND VPWR VPWR _279_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _435_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ _335_/A _329_/B VGND VGND VPWR VPWR _338_/A sky130_fd_sc_hd__nand2_1
Xsplit8 split8/A VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__buf_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_431_ _430_/X _462_/Q _491_/Q VGND VGND VPWR VPWR _431_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _424_/X _291_/Y _292_/Y VGND VGND VPWR VPWR _477_/D sky130_fd_sc_hd__a21bo_1
X_362_ _361_/A _361_/C _456_/Q VGND VGND VPWR VPWR _363_/B sky130_fd_sc_hd__o21a_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_276_ _479_/Q VGND VGND VPWR VPWR _278_/C sky130_fd_sc_hd__clkinv_4
X_414_ _413_/X _454_/Q _467_/Q VGND VGND VPWR VPWR _414_/X sky130_fd_sc_hd__mux2_1
X_259_ _259_/A _480_/Q VGND VGND VPWR VPWR _259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_328_ _324_/Y _327_/Y _291_/Y VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__479__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput10 _399_/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__283__A2 _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_430_ _385_/X _462_/Q _430_/S VGND VGND VPWR VPWR _430_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_361_ _361_/A _456_/Q _361_/C VGND VGND VPWR VPWR _363_/A sky130_fd_sc_hd__nor3_1
Xrebuffer9 _454_/Q VGND VGND VPWR VPWR _341_/A sky130_fd_sc_hd__clkbuf_1
X_292_ _296_/A _477_/Q _335_/B VGND VGND VPWR VPWR _292_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ _460_/Q VGND VGND VPWR VPWR _278_/B sky130_fd_sc_hd__clkinv_4
X_413_ _337_/Y _454_/Q _417_/S VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_258_ _482_/Q _481_/Q VGND VGND VPWR VPWR _259_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_327_ _325_/Y _326_/X _284_/C VGND VGND VPWR VPWR _327_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput11 _393_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__485__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ _291_/A _329_/B VGND VGND VPWR VPWR _291_/Y sky130_fd_sc_hd__nand2_2
X_360_ _473_/Q _472_/Q VGND VGND VPWR VPWR _360_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_489_ _489_/CLK _489_/D _347_/S VGND VGND VPWR VPWR _489_/Q sky130_fd_sc_hd__dfrtp_1
X_274_ _493_/Q _494_/Q _492_/Q VGND VGND VPWR VPWR _434_/S sky130_fd_sc_hd__nor3b_2
X_343_ _463_/Q _343_/B VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__xnor2_1
X_412_ _365_/X _363_/B _467_/Q VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__mux2_1
XANTENNA__477__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_257_ _397_/S _257_/B _430_/S VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ _440_/D _440_/Q VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__and2_1
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _466_/Q _465_/Q _464_/Q VGND VGND VPWR VPWR _417_/S sky130_fd_sc_hd__nor3b_2
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__445__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput12 _400_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_488_ _489_/CLK _488_/D _347_/S VGND VGND VPWR VPWR _488_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__422__A1 _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ _290_/A _335_/B _290_/C VGND VGND VPWR VPWR _478_/D sky130_fd_sc_hd__nand3_1
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
X_273_ _271_/Y _272_/A _272_/Y VGND VGND VPWR VPWR _480_/D sky130_fd_sc_hd__o21ai_1
X_411_ _360_/Y _363_/Y _467_/Q VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__mux2_1
X_342_ _342_/A _342_/B _468_/Q VGND VGND VPWR VPWR _343_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_256_ _482_/Q _481_/Q _480_/Q VGND VGND VPWR VPWR _430_/S sky130_fd_sc_hd__nor3b_2
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_325_ _440_/D _440_/Q VGND VGND VPWR VPWR _325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_239_ _243_/A _269_/B _489_/Q VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__nand3_1
X_308_ _471_/Q VGND VGND VPWR VPWR _310_/B sky130_fd_sc_hd__inv_2
XANTENNA__468__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_487_ _437_/A1 _487_/D _347_/S VGND VGND VPWR VPWR _487_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_345__8 _399_/X VGND VGND VPWR VPWR _446_/CLK sky130_fd_sc_hd__inv_4
X_272_ _272_/A _402_/X VGND VGND VPWR VPWR _272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_410_ _358_/Y _359_/Y _467_/Q VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__mux2_1
X_341_ _341_/A VGND VGND VPWR VPWR _342_/B sky130_fd_sc_hd__clkinv_4
XANTENNA__486__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_255_ _483_/Q VGND VGND VPWR VPWR _257_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_324_ _324_/A _324_/B _438_/Q VGND VGND VPWR VPWR _324_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_238_ _238_/A _269_/B _238_/C VGND VGND VPWR VPWR _490_/D sky130_fd_sc_hd__nand3_1
X_307_ _456_/Q _455_/Q _454_/Q _306_/Y VGND VGND VPWR VPWR _398_/S sky130_fd_sc_hd__o211a_1
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_486_ _489_/CLK _486_/D _347_/S VGND VGND VPWR VPWR _486_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ _480_/Q VGND VGND VPWR VPWR _271_/Y sky130_fd_sc_hd__inv_2
X_340_ _470_/Q _469_/Q VGND VGND VPWR VPWR _342_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_469_ _478_/CLK _469_/D _347_/S VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_2
X_254_ _462_/Q _461_/Q _460_/Q _253_/Y VGND VGND VPWR VPWR _397_/S sky130_fd_sc_hd__o211a_1
X_323_ _439_/Q _439_/D VGND VGND VPWR VPWR _324_/B sky130_fd_sc_hd__or2b_1
X_237_ _243_/A _353_/A _234_/B VGND VGND VPWR VPWR _238_/C sky130_fd_sc_hd__o21bai_1
X_306_ _474_/Q _473_/Q VGND VGND VPWR VPWR _306_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__470__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__425__A1 _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_485_ _485_/CLK _485_/D _347_/S VGND VGND VPWR VPWR _485_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _270_/A _270_/B VGND VGND VPWR VPWR _481_/D sky130_fd_sc_hd__nand2_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_399_ _436_/X _355_/Y _449_/Q VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__mux2_1
X_468_ _478_/CLK _468_/D _347_/S VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ _439_/D _439_/Q VGND VGND VPWR VPWR _324_/A sky130_fd_sc_hd__or2b_1
X_253_ _486_/Q _485_/Q VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_236_ _236_/A VGND VGND VPWR VPWR _243_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _437_/A1 sky130_fd_sc_hd__clkbuf_2
X_219_ _219_/A VGND VGND VPWR VPWR _492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__449__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_484_ _489_/CLK _484_/D _347_/S VGND VGND VPWR VPWR _484_/Q sky130_fd_sc_hd__dfrtn_1
X_398_ _291_/Y _467_/Q _398_/S VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__mux2_2
XANTENNA__464__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_467_ _435_/A1 _467_/D _347_/S VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_321_ _321_/A VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _489_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__463__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_235_ _263_/B VGND VGND VPWR VPWR _269_/B sky130_fd_sc_hd__clkbuf_2
X_304_ _304_/A VGND VGND VPWR VPWR _472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ _409_/X _492_/Q _460_/Q VGND VGND VPWR VPWR _219_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _436_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_483_ _483_/CLK _483_/D _347_/S VGND VGND VPWR VPWR _483_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _478_/CLK sky130_fd_sc_hd__clkbuf_2
X_397_ _229_/Y _491_/Q _397_/S VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__mux2_1
X_466_ _435_/A1 _466_/D _347_/S VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfrtn_1
X_251_ _251_/A VGND VGND VPWR VPWR _484_/D sky130_fd_sc_hd__clkbuf_1
X_320_ _425_/X _468_/Q _320_/S VGND VGND VPWR VPWR _321_/A sky130_fd_sc_hd__mux2_1
X_449_ _435_/A1 _449_/D _347_/S VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfrtp_1
X_234_ _353_/A _234_/B _234_/C VGND VGND VPWR VPWR _238_/A sky130_fd_sc_hd__nand3b_1
X_303_ _472_/Q _410_/X _398_/X VGND VGND VPWR VPWR _304_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_217_ _217_/A VGND VGND VPWR VPWR _493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_482_ _489_/CLK _482_/D _347_/S VGND VGND VPWR VPWR _482_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__446__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_465_ _465_/CLK _465_/D _347_/S VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ _484_/Q _427_/X _397_/X VGND VGND VPWR VPWR _251_/A sky130_fd_sc_hd__mux2_1
X_305__5 _435_/A1 VGND VGND VPWR VPWR _471_/CLK sky130_fd_sc_hd__inv_4
X_379_ _460_/Q _461_/Q _462_/Q VGND VGND VPWR VPWR _380_/B sky130_fd_sc_hd__o21a_1
XANTENNA__492__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_448_ _435_/A1 _448_/D _347_/S VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__347__S _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_233_ _490_/Q VGND VGND VPWR VPWR _234_/B sky130_fd_sc_hd__inv_2
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_302_ _302_/A VGND VGND VPWR VPWR _473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ _434_/X _493_/Q _460_/Q VGND VGND VPWR VPWR _217_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_481_ _481_/CLK _481_/D _347_/S VGND VGND VPWR VPWR _481_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_464_ _435_/A1 _464_/D _347_/S VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfrtn_1
X_395_ _494_/Q _395_/B VGND VGND VPWR VPWR _494_/D sky130_fd_sc_hd__xor2_1
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__452__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_447_ _447_/CLK _447_/D _347_/S VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfstp_1
X_378_ _460_/Q _462_/Q _461_/Q VGND VGND VPWR VPWR _380_/A sky130_fd_sc_hd__nor3_1
X_232_ _232_/A _487_/Q VGND VGND VPWR VPWR _353_/A sky130_fd_sc_hd__nand2_1
X_301_ _473_/Q _411_/X _398_/X VGND VGND VPWR VPWR _302_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__467__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_480_ _489_/CLK _480_/D _347_/S VGND VGND VPWR VPWR _480_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_394_ _493_/Q _460_/Q _492_/Q VGND VGND VPWR VPWR _395_/B sky130_fd_sc_hd__nor3_1
XFILLER_4_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ _435_/A1 _463_/D _347_/S VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__482__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_446_ _446_/CLK hold2/X _347_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfstp_1
X_377_ _485_/Q _484_/Q VGND VGND VPWR VPWR _377_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
X_231_ _489_/Q _488_/Q VGND VGND VPWR VPWR _232_/A sky130_fd_sc_hd__nor2_1
X_429_ _382_/X _380_/B _491_/Q VGND VGND VPWR VPWR _429_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _392_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__481__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_393_ _393_/A _445_/Q VGND VGND VPWR VPWR _393_/Y sky130_fd_sc_hd__nor2_1
X_462_ _357_/Y _462_/D _347_/S VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__451__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_445_ _445_/CLK hold3/X _347_/S VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfstp_1
X_376_ _460_/Q _461_/Q VGND VGND VPWR VPWR _376_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _222_/Y _226_/Y _229_/Y VGND VGND VPWR VPWR _491_/D sky130_fd_sc_hd__o21a_1
X_428_ _377_/Y _380_/Y _491_/Q VGND VGND VPWR VPWR _428_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_359_ _361_/A _361_/C VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__xnor2_1
Xinput2 ext_reset VGND VGND VPWR VPWR _393_/A sky130_fd_sc_hd__clkbuf_1
X_267__3 _489_/CLK VGND VGND VPWR VPWR _481_/CLK sky130_fd_sc_hd__inv_4
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__458__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_461_ _357_/Y _461_/D _347_/S VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_392_ _392_/A VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__clkinv_4
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__491__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_444_ _478_/CLK _444_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
X_375_ _484_/Q VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__clkinv_2
X_427_ _375_/Y _376_/Y _491_/Q VGND VGND VPWR VPWR _427_/X sky130_fd_sc_hd__mux2_1
X_358_ _472_/Q VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__clkinv_2
Xinput3 resetb VGND VGND VPWR VPWR _347_/S sky130_fd_sc_hd__buf_12
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _296_/A _352_/A _284_/B VGND VGND VPWR VPWR _290_/C sky130_fd_sc_hd__o21bai_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__421__A1 _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_460_ _357_/Y _460_/D _347_/S VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtp_4
X_391_ _493_/Q _492_/Q VGND VGND VPWR VPWR _391_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__460__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_443_ _437_/A1 _462_/Q VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfxtp_1
X_374_ _469_/Q _468_/Q VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_357_ _278_/B _437_/X _243_/A _356_/Y VGND VGND VPWR VPWR _357_/Y sky130_fd_sc_hd__o2bb2ai_2
Xinput4 sel2[0] VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__clkbuf_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _291_/A VGND VGND VPWR VPWR _296_/A sky130_fd_sc_hd__clkbuf_2
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _374_/Y _440_/D _426_/S VGND VGND VPWR VPWR _426_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_409_ _390_/Y _461_/Q _434_/S VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_390_ _492_/Q VGND VGND VPWR VPWR _390_/Y sky130_fd_sc_hd__clkinv_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_346__7 _399_/X VGND VGND VPWR VPWR _445_/CLK sky130_fd_sc_hd__inv_4
X_442_ _489_/CLK _461_/Q VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_373_ _468_/Q VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__447__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 sel2[1] VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__clkbuf_1
X_356_ _490_/Q _483_/Q VGND VGND VPWR VPWR _356_/Y sky130_fd_sc_hd__xnor2_1
X_287_ _456_/Q _455_/Q _454_/Q VGND VGND VPWR VPWR _291_/A sky130_fd_sc_hd__o21ai_1
X_425_ _373_/Y _439_/D _426_/S VGND VGND VPWR VPWR _425_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_408_ _407_/X _462_/Q _491_/Q VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__mux2_1
X_339_ _337_/Y _338_/A _338_/Y VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__454__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_441_ _437_/A1 _460_/Q VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_372_ _477_/Q _372_/B VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__xor2_1
Xclkbuf_1_0_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _347_/A1 sky130_fd_sc_hd__clkbuf_2
X_286_ _329_/B VGND VGND VPWR VPWR _335_/B sky130_fd_sc_hd__clkbuf_2
X_424_ _423_/X _440_/D _467_/Q VGND VGND VPWR VPWR _424_/X sky130_fd_sc_hd__mux2_1
X_355_ _342_/B _435_/X _296_/A _354_/Y VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__o2bb2ai_2
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 sel2[2] VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__clkbuf_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _269_/A _269_/B _481_/Q VGND VGND VPWR VPWR _270_/B sky130_fd_sc_hd__nand3_1
X_407_ _389_/X _462_/Q _432_/S VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__mux2_1
X_338_ _338_/A _414_/X VGND VGND VPWR VPWR _338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__494__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__349__B _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ _476_/Q _475_/Q VGND VGND VPWR VPWR _372_/B sky130_fd_sc_hd__nor2_1
X_440_ _435_/A1 _440_/D VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__476__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_285_ _467_/Q VGND VGND VPWR VPWR _329_/B sky130_fd_sc_hd__clkinv_4
X_423_ _372_/X split8/A _423_/S VGND VGND VPWR VPWR _423_/X sky130_fd_sc_hd__mux2_1
X_354_ _478_/Q _471_/Q VGND VGND VPWR VPWR _354_/Y sky130_fd_sc_hd__xnor2_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _451_/D sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__448__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ _272_/A _404_/X VGND VGND VPWR VPWR _270_/A sky130_fd_sc_hd__nand2_1
X_406_ _405_/X _461_/Q _491_/Q VGND VGND VPWR VPWR _406_/X sky130_fd_sc_hd__mux2_1
X_337_ _464_/Q VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _476_/Q _475_/Q VGND VGND VPWR VPWR _370_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_353_ _353_/A VGND VGND VPWR VPWR _432_/S sky130_fd_sc_hd__clkinv_4
X_422_ _421_/X _439_/D _467_/Q VGND VGND VPWR VPWR _422_/X sky130_fd_sc_hd__mux2_1
X_284_ _352_/A _284_/B _284_/C VGND VGND VPWR VPWR _290_/A sky130_fd_sc_hd__nand3b_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 sel[1] VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_405_ _387_/Y _461_/Q _432_/S VGND VGND VPWR VPWR _405_/X sky130_fd_sc_hd__mux2_1
X_336_ _336_/A _336_/B VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__nand2_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__439__D _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_319_ _319_/A VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_300__4 _478_/CLK VGND VGND VPWR VPWR _473_/CLK sky130_fd_sc_hd__inv_4
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_421_ _370_/Y _439_/D _423_/S VGND VGND VPWR VPWR _421_/X sky130_fd_sc_hd__mux2_1
Xinput9 sel[2] VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__clkbuf_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _352_/A VGND VGND VPWR VPWR _423_/S sky130_fd_sc_hd__clkinv_4
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _440_/D _439_/D _454_/Q VGND VGND VPWR VPWR _284_/C sky130_fd_sc_hd__o21a_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_266_ _266_/A _266_/B VGND VGND VPWR VPWR _482_/D sky130_fd_sc_hd__nand2_1
X_404_ _403_/X _461_/Q _491_/Q VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__mux2_1
X_335_ _335_/A _335_/B _465_/Q VGND VGND VPWR VPWR _336_/B sky130_fd_sc_hd__nand3_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_249_ _249_/A VGND VGND VPWR VPWR _485_/D sky130_fd_sc_hd__clkbuf_1
X_318_ _426_/X _469_/Q _320_/S VGND VGND VPWR VPWR _319_/A sky130_fd_sc_hd__mux2_1
XANTENNA__472__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_396__13 VGND VGND VPWR VPWR _396__13/HI _447_/D sky130_fd_sc_hd__conb_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__465__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_420_ _419_/X _420_/A1 _467_/Q VGND VGND VPWR VPWR _420_/X sky130_fd_sc_hd__mux2_1
X_282_ _478_/Q VGND VGND VPWR VPWR _284_/B sky130_fd_sc_hd__inv_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ _470_/Q _469_/Q _468_/Q VGND VGND VPWR VPWR _426_/S sky130_fd_sc_hd__nor3b_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_403_ _383_/Y _461_/Q _430_/S VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__mux2_1
X_334_ _338_/A _416_/X VGND VGND VPWR VPWR _336_/A sky130_fd_sc_hd__nand2_1
XANTENNA__323__B_N _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_265_ _269_/A _269_/B _482_/Q VGND VGND VPWR VPWR _266_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_248_ _485_/Q _428_/X _397_/X VGND VGND VPWR VPWR _249_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_317_ _470_/Q _317_/B VGND VGND VPWR VPWR _470_/D sky130_fd_sc_hd__xor2_1
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__488__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__471__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_350_ _462_/Q _461_/Q VGND VGND VPWR VPWR _437_/S sky130_fd_sc_hd__nor2_1
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_281_ _281_/A _475_/Q VGND VGND VPWR VPWR _352_/A sky130_fd_sc_hd__nand2_1
X_479_ _437_/A1 _479_/D _347_/S VGND VGND VPWR VPWR _479_/Q sky130_fd_sc_hd__dfstp_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__466__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_264_ _272_/A _431_/X VGND VGND VPWR VPWR _266_/A sky130_fd_sc_hd__nand2_1
X_402_ _401_/X _460_/Q _491_/Q VGND VGND VPWR VPWR _402_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_316_ _454_/Q _469_/Q _468_/Q VGND VGND VPWR VPWR _317_/B sky130_fd_sc_hd__nor3_1
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ _477_/Q _476_/Q VGND VGND VPWR VPWR _281_/A sky130_fd_sc_hd__nor2_1
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_478_ _478_/CLK _478_/D _347_/S VGND VGND VPWR VPWR _478_/Q sky130_fd_sc_hd__dfstp_1
X_263_ _269_/A _263_/B VGND VGND VPWR VPWR _272_/A sky130_fd_sc_hd__nand2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_401_ _271_/Y _460_/Q _430_/S VGND VGND VPWR VPWR _401_/X sky130_fd_sc_hd__mux2_1
X_332_ _332_/A _332_/B VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__nand2_1
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_246_ _246_/A VGND VGND VPWR VPWR _486_/D sky130_fd_sc_hd__clkbuf_1
X_315_ _315_/A _315_/B _335_/B VGND VGND VPWR VPWR _471_/D sky130_fd_sc_hd__nand3_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__450__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_229_ _236_/A _263_/B VGND VGND VPWR VPWR _229_/Y sky130_fd_sc_hd__nand2_2
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_494_ _437_/A1 _494_/D _347_/S VGND VGND VPWR VPWR _494_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_477_ _478_/CLK _477_/D _347_/S VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfrtp_1
X_262_ _262_/A _262_/B _269_/B VGND VGND VPWR VPWR _483_/D sky130_fd_sc_hd__nand3_1
X_400_ _436_/X _357_/Y _449_/Q VGND VGND VPWR VPWR _400_/X sky130_fd_sc_hd__mux2_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _335_/A _335_/B _466_/Q VGND VGND VPWR VPWR _332_/B sky130_fd_sc_hd__nand3_1
XANTENNA__475__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_245_ _486_/Q _429_/X _397_/X VGND VGND VPWR VPWR _246_/A sky130_fd_sc_hd__mux2_1
X_314_ _312_/Y _335_/A _310_/B VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__o21bai_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_228_ _491_/Q VGND VGND VPWR VPWR _263_/B sky130_fd_sc_hd__clkinv_4
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_493_ _437_/A1 _493_/D _347_/S VGND VGND VPWR VPWR _493_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__322__A _439_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ _478_/CLK _476_/D _347_/S VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfstp_1
X_261_ _259_/Y _269_/A _257_/B VGND VGND VPWR VPWR _262_/B sky130_fd_sc_hd__o21bai_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _338_/A _418_/X VGND VGND VPWR VPWR _332_/A sky130_fd_sc_hd__nand2_1
X_333__6 _435_/A1 VGND VGND VPWR VPWR _465_/CLK sky130_fd_sc_hd__inv_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ _357_/Y _459_/D _347_/S VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__dfrtp_1
X_244_ _433_/X _229_/Y _243_/Y VGND VGND VPWR VPWR _487_/D sky130_fd_sc_hd__a21bo_1
X_313_ _313_/A1 _313_/A2 _313_/B1 _306_/Y VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__483__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_227_ _462_/Q _461_/Q _460_/Q VGND VGND VPWR VPWR _236_/A sky130_fd_sc_hd__o21ai_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__469__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_492_ _437_/A1 _492_/D _347_/S VGND VGND VPWR VPWR _492_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_475_ _435_/A1 _475_/D _347_/S VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_260_ _462_/Q _461_/Q _460_/Q _253_/Y VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__o211ai_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_458_ _357_/Y _458_/D _347_/S VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__dfstp_1
X_389_ _489_/Q _389_/B VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__xor2_1
XANTENNA__484__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_243_ _243_/A _263_/B _487_/Q VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_312_ _312_/A _464_/Q VGND VGND VPWR VPWR _312_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_226_ _223_/Y _224_/X _234_/C VGND VGND VPWR VPWR _226_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_491_ _437_/A1 _491_/D _347_/S VGND VGND VPWR VPWR _491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_474_ _478_/CLK _474_/D _347_/S VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfrtn_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__453__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_388_ _488_/Q _487_/Q VGND VGND VPWR VPWR _389_/B sky130_fd_sc_hd__nor2_1
X_457_ _357_/Y _457_/D _347_/S VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__dfrtp_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ _406_/X _229_/Y _241_/Y VGND VGND VPWR VPWR _488_/D sky130_fd_sc_hd__a21bo_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ _466_/Q _465_/Q VGND VGND VPWR VPWR _312_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_225_ _462_/Q _461_/Q _460_/Q VGND VGND VPWR VPWR _234_/C sky130_fd_sc_hd__o21a_1
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_490_ _437_/A1 _490_/D _347_/S VGND VGND VPWR VPWR _490_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_473_ _473_/CLK _473_/D _347_/S VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfstp_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__493__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_387_ _488_/Q _487_/Q VGND VGND VPWR VPWR _387_/Y sky130_fd_sc_hd__xnor2_1
X_456_ _355_/Y _456_/D _347_/S VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _310_/A _310_/B _417_/S VGND VGND VPWR VPWR _315_/A sky130_fd_sc_hd__nand3_1
X_241_ _243_/A _263_/B _488_/Q VGND VGND VPWR VPWR _241_/Y sky130_fd_sc_hd__nand3_1
X_439_ _435_/A1 _439_/D VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfxtp_1
X_224_ _462_/Q _443_/Q VGND VGND VPWR VPWR _224_/X sky130_fd_sc_hd__and2_1
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_472_ _478_/CLK _472_/D _347_/S VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfrtn_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer10 _454_/Q VGND VGND VPWR VPWR _313_/B1 sky130_fd_sc_hd__clkbuf_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__462__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_386_ _487_/Q VGND VGND VPWR VPWR _386_/Y sky130_fd_sc_hd__clkinv_2
X_455_ _355_/Y _455_/D _347_/S VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfstp_4
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_344__9 _399_/X VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__inv_4
X_240_ _408_/X _229_/Y _239_/Y VGND VGND VPWR VPWR _489_/D sky130_fd_sc_hd__a21bo_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_369_ _475_/Q VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__clkinv_2
X_438_ _435_/A1 _454_/Q VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfxtp_1
X_223_ _462_/Q _443_/Q VGND VGND VPWR VPWR _223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__487__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsplit15 _456_/Q VGND VGND VPWR VPWR split8/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__455__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_471_ _471_/CLK _471_/D _347_/S VGND VGND VPWR VPWR _471_/Q sky130_fd_sc_hd__dfstp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 _454_/Q VGND VGND VPWR VPWR _361_/A sky130_fd_sc_hd__clkbuf_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ _482_/Q _385_/B VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__xor2_1
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_454_ _355_/Y _454_/D _347_/S VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ _479_/Q _437_/A1 _437_/S VGND VGND VPWR VPWR _437_/X sky130_fd_sc_hd__mux2_1
X_368_ _466_/Q _368_/B VGND VGND VPWR VPWR _368_/X sky130_fd_sc_hd__xor2_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_299_ _299_/A VGND VGND VPWR VPWR _474_/D sky130_fd_sc_hd__clkbuf_1
X_222_ _222_/A _222_/B _441_/Q VGND VGND VPWR VPWR _222_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__478__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__456__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__461__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_470_ _478_/CLK _470_/D _347_/S VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer12 _361_/A VGND VGND VPWR VPWR _320_/S sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _481_/Q _480_/Q VGND VGND VPWR VPWR _385_/B sky130_fd_sc_hd__nor2_1
X_453_ _355_/Y _453_/D _347_/S VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__dfrtp_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_436_ _436_/A0 _450_/Q _449_/D VGND VGND VPWR VPWR _436_/X sky130_fd_sc_hd__mux2_1
X_367_ _465_/Q _464_/Q VGND VGND VPWR VPWR _368_/B sky130_fd_sc_hd__nor2_1
X_298_ _474_/Q _412_/X _398_/X VGND VGND VPWR VPWR _299_/A sky130_fd_sc_hd__mux2_1
X_221_ _442_/Q _461_/Q VGND VGND VPWR VPWR _222_/B sky130_fd_sc_hd__or2b_1
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_419_ _369_/Y _419_/A1 _423_/S VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit4 _455_/Q VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__clkbuf_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer13 _454_/Q VGND VGND VPWR VPWR _419_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_383_ _481_/Q _480_/Q VGND VGND VPWR VPWR _383_/Y sky130_fd_sc_hd__xnor2_1
X_452_ _355_/Y _452_/D _347_/S VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__dfstp_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_366_ _465_/Q _464_/Q VGND VGND VPWR VPWR _366_/Y sky130_fd_sc_hd__xnor2_1
X_297_ _420_/X _291_/Y _296_/Y VGND VGND VPWR VPWR _475_/D sky130_fd_sc_hd__a21bo_1
X_435_ _463_/Q _435_/A1 _435_/S VGND VGND VPWR VPWR _435_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_220_ _461_/Q _442_/Q VGND VGND VPWR VPWR _222_/A sky130_fd_sc_hd__or2b_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_349_ _440_/D _439_/D VGND VGND VPWR VPWR _435_/S sky130_fd_sc_hd__nor2_1
X_418_ _417_/X split8/A _467_/Q VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__490__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247__1 _489_/CLK VGND VGND VPWR VPWR _485_/CLK sky130_fd_sc_hd__inv_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer14 _419_/A1 VGND VGND VPWR VPWR _420_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__480__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_382_ _486_/Q _382_/B VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__xor2_1
X_451_ _355_/Y _451_/D _347_/S VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__dfrtp_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ _391_/Y _462_/Q _434_/S VGND VGND VPWR VPWR _434_/X sky130_fd_sc_hd__mux2_1
X_296_ _296_/A _475_/Q _329_/B VGND VGND VPWR VPWR _296_/Y sky130_fd_sc_hd__nand3_1
X_365_ _474_/Q _365_/B VGND VGND VPWR VPWR _365_/X sky130_fd_sc_hd__xor2_1
Xrebuffer5 split8/A VGND VGND VPWR VPWR _313_/A1 sky130_fd_sc_hd__clkbuf_1
X_348_ _348_/A VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__buf_1
X_279_ _279_/A _279_/B VGND VGND VPWR VPWR _479_/D sky130_fd_sc_hd__nand2_1
X_417_ _368_/X _456_/Q _417_/S VGND VGND VPWR VPWR _417_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_252__2 _489_/CLK VGND VGND VPWR VPWR _483_/CLK sky130_fd_sc_hd__inv_4
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_450_ _435_/A1 hold1/X _347_/S VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfrtp_1
X_381_ _485_/Q _484_/Q VGND VGND VPWR VPWR _382_/B sky130_fd_sc_hd__nor2_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _432_/X _460_/Q _491_/Q VGND VGND VPWR VPWR _433_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ _422_/X _291_/Y _294_/Y VGND VGND VPWR VPWR _476_/D sky130_fd_sc_hd__a21bo_1
X_364_ _473_/Q _472_/Q VGND VGND VPWR VPWR _365_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer6 _455_/Q VGND VGND VPWR VPWR _313_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_347_ hold1/A _347_/A1 _347_/S VGND VGND VPWR VPWR _348_/A sky130_fd_sc_hd__mux2_2
XANTENNA__459__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ _434_/S _278_/B _278_/C VGND VGND VPWR VPWR _279_/B sky130_fd_sc_hd__nand3_1
X_416_ _415_/X _455_/Q _467_/Q VGND VGND VPWR VPWR _416_/X sky130_fd_sc_hd__mux2_1
XANTENNA__473__SET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__474__RESET_B _347_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer16 _398_/S VGND VGND VPWR VPWR _310_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_380_ _380_/A _380_/B VGND VGND VPWR VPWR _380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

