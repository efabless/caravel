magic
tech sky130A
magscale 1 2
timestamp 1686252151
<< obsm1 >>
rect 4 953326 633378 953378
rect 4 0 56 953326
rect 633326 0 633378 953326
rect 4 -52 633378 0
<< metal2 >>
rect 27497 953270 27558 953726
rect 29498 953270 29559 953726
rect 34054 953689 34102 953726
rect 34046 953637 34110 953689
rect 34360 953270 34416 953750
rect 34912 953270 34968 953750
rect 35556 953270 35612 953750
rect 36200 953270 36256 953750
rect 36752 953603 36808 953726
rect 36692 953539 36864 953603
rect 36752 953270 36808 953539
rect 37396 953507 37452 953726
rect 37396 953443 37570 953507
rect 37396 953270 37452 953443
rect 38040 953270 38096 953750
rect 38592 953270 38648 953750
rect 39236 953270 39292 953750
rect 39880 953270 39936 953750
rect 40432 953411 40488 953726
rect 41076 953603 41132 953726
rect 41013 953539 41197 953603
rect 40432 953347 40605 953411
rect 40432 953270 40488 953347
rect 41076 953270 41132 953539
rect 41720 953507 41776 953726
rect 41720 953443 41894 953507
rect 41720 953270 41776 953443
rect 42364 953270 42420 953750
rect 42916 953270 42972 953750
rect 43560 953270 43616 953750
rect 44204 953270 44260 953750
rect 44756 953270 44812 953750
rect 45400 953270 45456 953750
rect 46044 953270 46100 953726
rect 46596 953270 46652 953750
rect 47240 953270 47296 953750
rect 47884 953270 47940 953726
rect 48436 953270 48492 953726
rect 49080 953270 49136 953750
rect 49724 953507 49780 953726
rect 49607 953443 49780 953507
rect 49724 953270 49780 953443
rect 78697 953270 78758 953726
rect 80698 953270 80759 953726
rect 85454 953689 85502 953726
rect 85446 953637 85510 953689
rect 85760 953270 85816 953750
rect 86312 953270 86368 953750
rect 86956 953270 87012 953750
rect 87600 953270 87656 953750
rect 88152 953603 88208 953726
rect 88092 953539 88264 953603
rect 88152 953270 88208 953539
rect 88796 953507 88852 953726
rect 88796 953443 88970 953507
rect 88796 953270 88852 953443
rect 89440 953270 89496 953750
rect 89992 953270 90048 953750
rect 90636 953270 90692 953750
rect 91280 953270 91336 953750
rect 91832 953411 91888 953726
rect 92476 953603 92532 953726
rect 92413 953539 92597 953603
rect 91832 953347 92005 953411
rect 91832 953270 91888 953347
rect 92476 953270 92532 953539
rect 93120 953507 93176 953726
rect 93120 953443 93294 953507
rect 93120 953270 93176 953443
rect 93764 953270 93820 953750
rect 94316 953270 94372 953750
rect 94960 953270 95016 953750
rect 95604 953270 95660 953750
rect 96156 953270 96212 953750
rect 96800 953270 96856 953750
rect 97444 953270 97500 953726
rect 97996 953270 98052 953750
rect 98640 953270 98696 953750
rect 99284 953270 99340 953726
rect 99836 953270 99892 953726
rect 100480 953270 100536 953750
rect 101124 953507 101180 953726
rect 101007 953443 101180 953507
rect 101124 953270 101180 953443
rect 129897 953270 129958 953726
rect 131898 953270 131959 953726
rect 136854 953689 136902 953726
rect 136846 953637 136910 953689
rect 137160 953270 137216 953750
rect 137712 953270 137768 953750
rect 138356 953270 138412 953750
rect 139000 953270 139056 953750
rect 139552 953603 139608 953726
rect 139492 953539 139664 953603
rect 139552 953270 139608 953539
rect 140196 953507 140252 953726
rect 140196 953443 140370 953507
rect 140196 953270 140252 953443
rect 140840 953270 140896 953750
rect 141392 953270 141448 953750
rect 142036 953270 142092 953750
rect 142680 953270 142736 953750
rect 143232 953411 143288 953726
rect 143876 953603 143932 953726
rect 143813 953539 143997 953603
rect 143232 953347 143405 953411
rect 143232 953270 143288 953347
rect 143876 953270 143932 953539
rect 144520 953507 144576 953726
rect 144520 953443 144694 953507
rect 144520 953270 144576 953443
rect 145164 953270 145220 953750
rect 145716 953270 145772 953750
rect 146360 953270 146416 953750
rect 147004 953270 147060 953750
rect 147556 953270 147612 953750
rect 148200 953270 148256 953750
rect 148844 953270 148900 953726
rect 149396 953270 149452 953750
rect 150040 953270 150096 953750
rect 150684 953270 150740 953726
rect 151236 953270 151292 953726
rect 151880 953270 151936 953750
rect 152524 953507 152580 953726
rect 152407 953443 152580 953507
rect 152524 953270 152580 953443
rect 181097 953270 181158 953726
rect 183098 953270 183159 953726
rect 188254 953689 188302 953726
rect 188246 953637 188310 953689
rect 188560 953270 188616 953750
rect 189112 953270 189168 953750
rect 189756 953270 189812 953750
rect 190400 953270 190456 953750
rect 190952 953603 191008 953726
rect 190892 953539 191064 953603
rect 190952 953270 191008 953539
rect 191596 953507 191652 953726
rect 191596 953443 191770 953507
rect 191596 953270 191652 953443
rect 192240 953270 192296 953750
rect 192792 953270 192848 953750
rect 193436 953270 193492 953750
rect 194080 953270 194136 953750
rect 194632 953411 194688 953726
rect 195276 953603 195332 953726
rect 195213 953539 195397 953603
rect 194632 953347 194805 953411
rect 194632 953270 194688 953347
rect 195276 953270 195332 953539
rect 195920 953507 195976 953726
rect 195920 953443 196094 953507
rect 195920 953270 195976 953443
rect 196564 953270 196620 953750
rect 197116 953270 197172 953750
rect 197760 953270 197816 953750
rect 198404 953270 198460 953750
rect 198956 953270 199012 953750
rect 199600 953270 199656 953750
rect 200244 953270 200300 953726
rect 200796 953270 200852 953750
rect 201440 953270 201496 953750
rect 202084 953270 202140 953726
rect 202636 953270 202692 953726
rect 203280 953270 203336 953750
rect 203924 953507 203980 953726
rect 203807 953443 203980 953507
rect 203924 953270 203980 953443
rect 232297 953270 232358 953726
rect 234298 953270 234359 953726
rect 239854 953689 239902 953726
rect 239846 953637 239910 953689
rect 240160 953270 240216 953750
rect 240712 953270 240768 953750
rect 241356 953270 241412 953750
rect 242000 953270 242056 953750
rect 242552 953603 242608 953726
rect 242492 953539 242664 953603
rect 242552 953270 242608 953539
rect 243196 953507 243252 953726
rect 243196 953443 243370 953507
rect 243196 953270 243252 953443
rect 243840 953270 243896 953750
rect 244392 953270 244448 953750
rect 245036 953270 245092 953750
rect 245680 953270 245736 953750
rect 246232 953411 246288 953726
rect 246876 953603 246932 953726
rect 246813 953539 246997 953603
rect 246232 953347 246405 953411
rect 246232 953270 246288 953347
rect 246876 953270 246932 953539
rect 247520 953507 247576 953726
rect 247520 953443 247694 953507
rect 247520 953270 247576 953443
rect 248164 953270 248220 953750
rect 248716 953270 248772 953750
rect 249360 953270 249416 953750
rect 250004 953270 250060 953750
rect 250556 953270 250612 953750
rect 251200 953270 251256 953750
rect 251844 953270 251900 953726
rect 252396 953270 252452 953750
rect 253040 953270 253096 953750
rect 253684 953270 253740 953726
rect 254236 953270 254292 953726
rect 254880 953270 254936 953750
rect 255524 953507 255580 953726
rect 255407 953443 255580 953507
rect 255524 953270 255580 953443
rect 336697 953270 336758 953726
rect 338698 953270 338759 953726
rect 341654 953689 341702 953726
rect 341646 953637 341710 953689
rect 341960 953270 342016 953750
rect 342512 953270 342568 953750
rect 343156 953270 343212 953750
rect 343800 953270 343856 953750
rect 344352 953603 344408 953726
rect 344292 953539 344464 953603
rect 344352 953270 344408 953539
rect 344996 953507 345052 953726
rect 344996 953443 345170 953507
rect 344996 953270 345052 953443
rect 345640 953270 345696 953750
rect 346192 953270 346248 953750
rect 346836 953270 346892 953750
rect 347480 953270 347536 953750
rect 348032 953411 348088 953726
rect 348676 953603 348732 953726
rect 348613 953539 348797 953603
rect 348032 953347 348205 953411
rect 348032 953270 348088 953347
rect 348676 953270 348732 953539
rect 349320 953507 349376 953726
rect 349320 953443 349494 953507
rect 349320 953270 349376 953443
rect 349964 953270 350020 953750
rect 350516 953270 350572 953750
rect 351160 953270 351216 953750
rect 351804 953270 351860 953750
rect 352356 953270 352412 953750
rect 353000 953270 353056 953750
rect 353644 953270 353700 953726
rect 354196 953270 354252 953750
rect 354840 953270 354896 953750
rect 355484 953270 355540 953726
rect 356036 953270 356092 953726
rect 356680 953270 356736 953750
rect 357324 953507 357380 953726
rect 357207 953443 357380 953507
rect 357324 953270 357380 953443
rect 425697 953270 425758 953726
rect 427698 953270 427759 953726
rect 430654 953689 430702 953726
rect 430646 953637 430710 953689
rect 430960 953270 431016 953750
rect 431512 953270 431568 953750
rect 432156 953270 432212 953750
rect 432800 953270 432856 953750
rect 433352 953603 433408 953726
rect 433292 953539 433464 953603
rect 433352 953270 433408 953539
rect 433996 953507 434052 953726
rect 433996 953443 434170 953507
rect 433996 953270 434052 953443
rect 434640 953270 434696 953750
rect 435192 953270 435248 953750
rect 435836 953270 435892 953750
rect 436480 953270 436536 953750
rect 437032 953411 437088 953726
rect 437676 953603 437732 953726
rect 437613 953539 437797 953603
rect 437032 953347 437205 953411
rect 437032 953270 437088 953347
rect 437676 953270 437732 953539
rect 438320 953507 438376 953726
rect 438320 953443 438494 953507
rect 438320 953270 438376 953443
rect 438964 953270 439020 953750
rect 439516 953270 439572 953750
rect 440160 953270 440216 953750
rect 440804 953270 440860 953750
rect 441356 953270 441412 953750
rect 442000 953270 442056 953750
rect 442644 953270 442700 953726
rect 443196 953270 443252 953750
rect 443840 953270 443896 953750
rect 444484 953270 444540 953726
rect 445036 953270 445092 953726
rect 445680 953270 445736 953750
rect 446324 953507 446380 953726
rect 446207 953443 446380 953507
rect 446324 953270 446380 953443
rect 476897 953270 476958 953726
rect 478898 953270 478959 953726
rect 482054 953689 482102 953726
rect 482046 953637 482110 953689
rect 482360 953270 482416 953750
rect 482912 953270 482968 953750
rect 483556 953270 483612 953750
rect 484200 953270 484256 953750
rect 484752 953603 484808 953726
rect 484692 953539 484864 953603
rect 484752 953270 484808 953539
rect 485396 953507 485452 953726
rect 485396 953443 485570 953507
rect 485396 953270 485452 953443
rect 486040 953270 486096 953750
rect 486592 953270 486648 953750
rect 487236 953270 487292 953750
rect 487880 953270 487936 953750
rect 488432 953411 488488 953726
rect 489076 953603 489132 953726
rect 489013 953539 489197 953603
rect 488432 953347 488605 953411
rect 488432 953270 488488 953347
rect 489076 953270 489132 953539
rect 489720 953507 489776 953726
rect 489720 953443 489894 953507
rect 489720 953270 489776 953443
rect 490364 953270 490420 953750
rect 490916 953270 490972 953750
rect 491560 953270 491616 953750
rect 492204 953270 492260 953750
rect 492756 953270 492812 953750
rect 493400 953270 493456 953750
rect 494044 953270 494100 953726
rect 494596 953270 494652 953750
rect 495240 953270 495296 953750
rect 495884 953270 495940 953726
rect 496436 953270 496492 953726
rect 497080 953270 497136 953750
rect 497724 953507 497780 953726
rect 497607 953443 497780 953507
rect 497724 953270 497780 953443
rect 576297 953270 576358 953726
rect 578298 953270 578359 953726
rect 583854 953689 583902 953726
rect 583846 953637 583910 953689
rect 584160 953270 584216 953750
rect 584712 953270 584768 953750
rect 585356 953270 585412 953750
rect 586000 953270 586056 953750
rect 586552 953603 586608 953726
rect 586492 953539 586664 953603
rect 586552 953270 586608 953539
rect 587196 953507 587252 953726
rect 587196 953443 587370 953507
rect 587196 953270 587252 953443
rect 587840 953270 587896 953750
rect 588392 953270 588448 953750
rect 589036 953270 589092 953750
rect 589680 953270 589736 953750
rect 590232 953411 590288 953726
rect 590876 953603 590932 953726
rect 590813 953539 590997 953603
rect 590232 953347 590405 953411
rect 590232 953270 590288 953347
rect 590876 953270 590932 953539
rect 591520 953507 591576 953726
rect 591520 953443 591694 953507
rect 591520 953270 591576 953443
rect 592164 953270 592220 953750
rect 592716 953270 592772 953750
rect 593360 953270 593416 953750
rect 594004 953270 594060 953750
rect 594556 953270 594612 953750
rect 595200 953270 595256 953750
rect 595844 953270 595900 953726
rect 596396 953270 596452 953750
rect 597040 953270 597096 953750
rect 597684 953270 597740 953726
rect 598236 953270 598292 953726
rect 598880 953270 598936 953750
rect 599524 953507 599580 953726
rect 599407 953443 599580 953507
rect 599524 953270 599580 953443
rect -400 927724 56 927780
rect -181 927607 -117 927724
rect -274 927136 56 927143
rect -400 927080 56 927136
rect -274 927073 56 927080
rect -400 926436 56 926492
rect -400 925884 56 925940
rect -274 925296 56 925303
rect -400 925240 56 925296
rect -274 925233 56 925240
rect 633270 925110 633726 925166
rect -274 924652 56 924659
rect -400 924596 56 924652
rect -274 924589 56 924596
rect 633270 924614 633600 924621
rect 633270 924558 633726 924614
rect 633270 924551 633600 924558
rect -400 924044 56 924100
rect 633270 923970 633600 923977
rect 633270 923914 633726 923970
rect 633270 923907 633600 923914
rect -274 923456 56 923463
rect -400 923400 56 923456
rect -274 923393 56 923400
rect 633270 923326 633600 923333
rect 633270 923270 633726 923326
rect 633270 923263 633600 923270
rect -400 922756 56 922812
rect 633539 922774 633603 922834
rect 633270 922718 633726 922774
rect 633539 922662 633603 922718
rect -274 922260 56 922267
rect -400 922204 56 922260
rect -274 922197 56 922204
rect 633270 922074 633726 922130
rect 633443 921956 633507 922074
rect -274 921616 56 921623
rect -400 921560 56 921616
rect -274 921553 56 921560
rect 633270 921486 633600 921493
rect 633270 921430 633726 921486
rect 633270 921423 633600 921430
rect -274 920972 56 920979
rect -400 920916 56 920972
rect -274 920909 56 920916
rect 633270 920934 633600 920941
rect 633270 920878 633726 920934
rect 633270 920871 633600 920878
rect -274 920420 56 920427
rect -400 920364 56 920420
rect -274 920357 56 920364
rect 633270 920290 633600 920297
rect 633270 920234 633726 920290
rect 633270 920227 633600 920234
rect -181 919776 -117 919894
rect -400 919720 56 919776
rect 633270 919646 633600 919653
rect 633270 919590 633726 919646
rect 633270 919583 633600 919590
rect -277 919132 -213 919197
rect -400 919076 56 919132
rect -277 919013 -213 919076
rect 633270 919038 633726 919094
rect 633347 918921 633411 919038
rect -85 918488 -21 918605
rect -400 918432 56 918488
rect 633539 918450 633603 918513
rect 633270 918394 633726 918450
rect 633539 918329 633603 918394
rect -274 917936 56 917943
rect -400 917880 56 917936
rect -274 917873 56 917880
rect 633270 917750 633726 917806
rect 633443 917632 633507 917750
rect -274 917292 56 917299
rect -400 917236 56 917292
rect -274 917229 56 917236
rect 633270 917162 633600 917169
rect 633270 917106 633726 917162
rect 633270 917099 633600 917106
rect -274 916648 56 916655
rect -400 916592 56 916648
rect -274 916585 56 916592
rect 633270 916610 633600 916617
rect 633270 916554 633726 916610
rect 633270 916547 633600 916554
rect -274 916096 56 916103
rect -400 916040 56 916096
rect -274 916033 56 916040
rect 633270 915966 633600 915973
rect 633270 915910 633726 915966
rect 633270 915903 633600 915910
rect -181 915452 -117 915570
rect -400 915396 56 915452
rect 633270 915322 633600 915329
rect 633270 915266 633726 915322
rect 633270 915259 633600 915266
rect -277 914808 -213 914864
rect -400 914752 56 914808
rect -277 914692 -213 914752
rect 633270 914714 633726 914770
rect -274 914256 56 914263
rect -400 914200 56 914256
rect -274 914193 56 914200
rect 633270 914126 633600 914133
rect 633270 914070 633726 914126
rect 633270 914063 633600 914070
rect -274 913612 56 913619
rect -400 913556 56 913612
rect -274 913549 56 913556
rect 633270 913426 633726 913482
rect -274 912968 56 912975
rect -400 912912 56 912968
rect -274 912905 56 912912
rect 633270 912930 633600 912937
rect 633270 912874 633726 912930
rect 633270 912867 633600 912874
rect -400 912360 56 912416
rect 633270 912286 633600 912293
rect 633270 912230 633726 912286
rect 633270 912223 633600 912230
rect 633270 911586 633726 911642
rect 633270 911034 633726 911090
rect 633270 910446 633600 910453
rect 633270 910390 633726 910446
rect 633270 910383 633600 910390
rect 633443 909802 633507 909919
rect 633270 909746 633726 909802
rect 633270 835910 633726 835966
rect 633270 835414 633600 835421
rect 633270 835358 633726 835414
rect 633270 835351 633600 835358
rect 633270 834770 633600 834777
rect 633270 834714 633726 834770
rect 633270 834707 633600 834714
rect 633270 834126 633600 834133
rect 633270 834070 633726 834126
rect 633270 834063 633600 834070
rect 633539 833574 633603 833634
rect 633270 833518 633726 833574
rect 633539 833462 633603 833518
rect 633270 832874 633726 832930
rect 633443 832756 633507 832874
rect 633270 832286 633600 832293
rect 633270 832230 633726 832286
rect 633270 832223 633600 832230
rect 633270 831734 633600 831741
rect 633270 831678 633726 831734
rect 633270 831671 633600 831678
rect 633270 831090 633600 831097
rect 633270 831034 633726 831090
rect 633270 831027 633600 831034
rect 633270 830446 633600 830453
rect 633270 830390 633726 830446
rect 633270 830383 633600 830390
rect 633270 829838 633726 829894
rect 633347 829721 633411 829838
rect 633539 829250 633603 829313
rect 633270 829194 633726 829250
rect 633539 829129 633603 829194
rect 633270 828550 633726 828606
rect 633443 828432 633507 828550
rect 633270 827962 633600 827969
rect 633270 827906 633726 827962
rect 633270 827899 633600 827906
rect 633270 827410 633600 827417
rect 633270 827354 633726 827410
rect 633270 827347 633600 827354
rect 633270 826766 633600 826773
rect 633270 826710 633726 826766
rect 633270 826703 633600 826710
rect 633270 826122 633600 826129
rect 633270 826066 633726 826122
rect 633270 826059 633600 826066
rect 633270 825514 633726 825570
rect 633270 824926 633600 824933
rect 633270 824870 633726 824926
rect 633270 824863 633600 824870
rect 633270 824226 633726 824282
rect 633270 823730 633600 823737
rect 633270 823674 633726 823730
rect 633270 823667 633600 823674
rect 633270 823086 633600 823093
rect 633270 823030 633726 823086
rect 633270 823023 633600 823030
rect 633270 822386 633726 822442
rect 633270 821834 633726 821890
rect 633270 821246 633600 821253
rect 633270 821190 633726 821246
rect 633270 821183 633600 821190
rect 633443 820602 633507 820719
rect 633270 820546 633726 820602
rect -400 757924 56 757980
rect -181 757807 -117 757924
rect -274 757336 56 757343
rect -400 757280 56 757336
rect -274 757273 56 757280
rect -400 756636 56 756692
rect -400 756084 56 756140
rect -274 755496 56 755503
rect -400 755440 56 755496
rect -274 755433 56 755440
rect -274 754852 56 754859
rect -400 754796 56 754852
rect -274 754789 56 754796
rect -400 754244 56 754300
rect -274 753656 56 753663
rect -400 753600 56 753656
rect -274 753593 56 753600
rect -400 752956 56 753012
rect -274 752460 56 752467
rect -400 752404 56 752460
rect -274 752397 56 752404
rect -274 751816 56 751823
rect -400 751760 56 751816
rect -274 751753 56 751760
rect -274 751172 56 751179
rect -400 751116 56 751172
rect -274 751109 56 751116
rect -274 750620 56 750627
rect -400 750564 56 750620
rect -274 750557 56 750564
rect -181 749976 -117 750094
rect -400 749920 56 749976
rect -277 749332 -213 749397
rect -400 749276 56 749332
rect -277 749213 -213 749276
rect -85 748688 -21 748805
rect -400 748632 56 748688
rect -274 748136 56 748143
rect -400 748080 56 748136
rect -274 748073 56 748080
rect -274 747492 56 747499
rect -400 747436 56 747492
rect -274 747429 56 747436
rect -274 746848 56 746855
rect -400 746792 56 746848
rect -274 746785 56 746792
rect 633270 746710 633726 746766
rect -274 746296 56 746303
rect -400 746240 56 746296
rect -274 746233 56 746240
rect 633270 746214 633600 746221
rect 633270 746158 633726 746214
rect 633270 746151 633600 746158
rect -181 745652 -117 745770
rect -400 745596 56 745652
rect 633270 745570 633600 745577
rect 633270 745514 633726 745570
rect 633270 745507 633600 745514
rect -277 745008 -213 745064
rect -400 744952 56 745008
rect -277 744892 -213 744952
rect 633270 744926 633600 744933
rect 633270 744870 633726 744926
rect 633270 744863 633600 744870
rect -274 744456 56 744463
rect -400 744400 56 744456
rect -274 744393 56 744400
rect 633539 744374 633603 744434
rect 633270 744318 633726 744374
rect 633539 744262 633603 744318
rect -274 743812 56 743819
rect -400 743756 56 743812
rect -274 743749 56 743756
rect 633270 743674 633726 743730
rect 633443 743556 633507 743674
rect -274 743168 56 743175
rect -400 743112 56 743168
rect -274 743105 56 743112
rect 633270 743086 633600 743093
rect 633270 743030 633726 743086
rect 633270 743023 633600 743030
rect -400 742560 56 742616
rect 633270 742534 633600 742541
rect 633270 742478 633726 742534
rect 633270 742471 633600 742478
rect 633270 741890 633600 741897
rect 633270 741834 633726 741890
rect 633270 741827 633600 741834
rect 633270 741246 633600 741253
rect 633270 741190 633726 741246
rect 633270 741183 633600 741190
rect 633270 740638 633726 740694
rect 633347 740521 633411 740638
rect 633539 740050 633603 740113
rect 633270 739994 633726 740050
rect 633539 739929 633603 739994
rect 633270 739350 633726 739406
rect 633443 739232 633507 739350
rect 633270 738762 633600 738769
rect 633270 738706 633726 738762
rect 633270 738699 633600 738706
rect 633270 738210 633600 738217
rect 633270 738154 633726 738210
rect 633270 738147 633600 738154
rect 633270 737566 633600 737573
rect 633270 737510 633726 737566
rect 633270 737503 633600 737510
rect 633270 736922 633600 736929
rect 633270 736866 633726 736922
rect 633270 736859 633600 736866
rect 633270 736314 633726 736370
rect 633270 735726 633600 735733
rect 633270 735670 633726 735726
rect 633270 735663 633600 735670
rect 633270 735026 633726 735082
rect 633270 734530 633600 734537
rect 633270 734474 633726 734530
rect 633270 734467 633600 734474
rect 633270 733886 633600 733893
rect 633270 733830 633726 733886
rect 633270 733823 633600 733830
rect 633270 733186 633726 733242
rect 633270 732634 633726 732690
rect 633270 732046 633600 732053
rect 633270 731990 633726 732046
rect 633270 731983 633600 731990
rect 633443 731402 633507 731519
rect 633270 731346 633726 731402
rect -400 714724 56 714780
rect -181 714607 -117 714724
rect -274 714136 56 714143
rect -400 714080 56 714136
rect -274 714073 56 714080
rect -400 713436 56 713492
rect -400 712884 56 712940
rect -274 712296 56 712303
rect -400 712240 56 712296
rect -274 712233 56 712240
rect -274 711652 56 711659
rect -400 711596 56 711652
rect -274 711589 56 711596
rect -400 711044 56 711100
rect -274 710456 56 710463
rect -400 710400 56 710456
rect -274 710393 56 710400
rect -400 709756 56 709812
rect -274 709260 56 709267
rect -400 709204 56 709260
rect -274 709197 56 709204
rect -274 708616 56 708623
rect -400 708560 56 708616
rect -274 708553 56 708560
rect -274 707972 56 707979
rect -400 707916 56 707972
rect -274 707909 56 707916
rect -274 707420 56 707427
rect -400 707364 56 707420
rect -274 707357 56 707364
rect -181 706776 -117 706894
rect -400 706720 56 706776
rect -277 706132 -213 706197
rect -400 706076 56 706132
rect -277 706013 -213 706076
rect -85 705488 -21 705605
rect -400 705432 56 705488
rect -274 704936 56 704943
rect -400 704880 56 704936
rect -274 704873 56 704880
rect -274 704292 56 704299
rect -400 704236 56 704292
rect -274 704229 56 704236
rect -274 703648 56 703655
rect -400 703592 56 703648
rect -274 703585 56 703592
rect -274 703096 56 703103
rect -400 703040 56 703096
rect -274 703033 56 703040
rect -181 702452 -117 702570
rect -400 702396 56 702452
rect -277 701808 -213 701864
rect -400 701752 56 701808
rect -277 701692 -213 701752
rect 633270 701710 633726 701766
rect -274 701256 56 701263
rect -400 701200 56 701256
rect -274 701193 56 701200
rect 633270 701214 633600 701221
rect 633270 701158 633726 701214
rect 633270 701151 633600 701158
rect -274 700612 56 700619
rect -400 700556 56 700612
rect -274 700549 56 700556
rect 633270 700570 633600 700577
rect 633270 700514 633726 700570
rect 633270 700507 633600 700514
rect -274 699968 56 699975
rect -400 699912 56 699968
rect -274 699905 56 699912
rect 633270 699926 633600 699933
rect 633270 699870 633726 699926
rect 633270 699863 633600 699870
rect -400 699360 56 699416
rect 633539 699374 633603 699434
rect 633270 699318 633726 699374
rect 633539 699262 633603 699318
rect 633270 698674 633726 698730
rect 633443 698556 633507 698674
rect 633270 698086 633600 698093
rect 633270 698030 633726 698086
rect 633270 698023 633600 698030
rect 633270 697534 633600 697541
rect 633270 697478 633726 697534
rect 633270 697471 633600 697478
rect 633270 696890 633600 696897
rect 633270 696834 633726 696890
rect 633270 696827 633600 696834
rect 633270 696246 633600 696253
rect 633270 696190 633726 696246
rect 633270 696183 633600 696190
rect 633270 695638 633726 695694
rect 633347 695521 633411 695638
rect 633539 695050 633603 695113
rect 633270 694994 633726 695050
rect 633539 694929 633603 694994
rect 633270 694350 633726 694406
rect 633443 694232 633507 694350
rect 633270 693762 633600 693769
rect 633270 693706 633726 693762
rect 633270 693699 633600 693706
rect 633270 693210 633600 693217
rect 633270 693154 633726 693210
rect 633270 693147 633600 693154
rect 633270 692566 633600 692573
rect 633270 692510 633726 692566
rect 633270 692503 633600 692510
rect 633270 691922 633600 691929
rect 633270 691866 633726 691922
rect 633270 691859 633600 691866
rect 633270 691314 633726 691370
rect 633270 690726 633600 690733
rect 633270 690670 633726 690726
rect 633270 690663 633600 690670
rect 633270 690026 633726 690082
rect 633270 689530 633600 689537
rect 633270 689474 633726 689530
rect 633270 689467 633600 689474
rect 633270 688886 633600 688893
rect 633270 688830 633726 688886
rect 633270 688823 633600 688830
rect 633270 688186 633726 688242
rect 633270 687634 633726 687690
rect 633270 687046 633600 687053
rect 633270 686990 633726 687046
rect 633270 686983 633600 686990
rect 633443 686402 633507 686519
rect 633270 686346 633726 686402
rect -400 671524 56 671580
rect -181 671407 -117 671524
rect -274 670936 56 670943
rect -400 670880 56 670936
rect -274 670873 56 670880
rect -400 670236 56 670292
rect -400 669684 56 669740
rect -274 669096 56 669103
rect -400 669040 56 669096
rect -274 669033 56 669040
rect -274 668452 56 668459
rect -400 668396 56 668452
rect -274 668389 56 668396
rect -400 667844 56 667900
rect -274 667256 56 667263
rect -400 667200 56 667256
rect -274 667193 56 667200
rect -400 666556 56 666612
rect -274 666060 56 666067
rect -400 666004 56 666060
rect -274 665997 56 666004
rect -274 665416 56 665423
rect -400 665360 56 665416
rect -274 665353 56 665360
rect -274 664772 56 664779
rect -400 664716 56 664772
rect -274 664709 56 664716
rect -274 664220 56 664227
rect -400 664164 56 664220
rect -274 664157 56 664164
rect -181 663576 -117 663694
rect -400 663520 56 663576
rect -277 662932 -213 662997
rect -400 662876 56 662932
rect -277 662813 -213 662876
rect -85 662288 -21 662405
rect -400 662232 56 662288
rect -274 661736 56 661743
rect -400 661680 56 661736
rect -274 661673 56 661680
rect -274 661092 56 661099
rect -400 661036 56 661092
rect -274 661029 56 661036
rect -274 660448 56 660455
rect -400 660392 56 660448
rect -274 660385 56 660392
rect -274 659896 56 659903
rect -400 659840 56 659896
rect -274 659833 56 659840
rect -181 659252 -117 659370
rect -400 659196 56 659252
rect -277 658608 -213 658664
rect -400 658552 56 658608
rect -277 658492 -213 658552
rect -274 658056 56 658063
rect -400 658000 56 658056
rect -274 657993 56 658000
rect -274 657412 56 657419
rect -400 657356 56 657412
rect -274 657349 56 657356
rect -274 656768 56 656775
rect -400 656712 56 656768
rect -274 656705 56 656712
rect 633270 656710 633726 656766
rect -400 656160 56 656216
rect 633270 656214 633600 656221
rect 633270 656158 633726 656214
rect 633270 656151 633600 656158
rect 633270 655570 633600 655577
rect 633270 655514 633726 655570
rect 633270 655507 633600 655514
rect 633270 654926 633600 654933
rect 633270 654870 633726 654926
rect 633270 654863 633600 654870
rect 633539 654374 633603 654434
rect 633270 654318 633726 654374
rect 633539 654262 633603 654318
rect 633270 653674 633726 653730
rect 633443 653556 633507 653674
rect 633270 653086 633600 653093
rect 633270 653030 633726 653086
rect 633270 653023 633600 653030
rect 633270 652534 633600 652541
rect 633270 652478 633726 652534
rect 633270 652471 633600 652478
rect 633270 651890 633600 651897
rect 633270 651834 633726 651890
rect 633270 651827 633600 651834
rect 633270 651246 633600 651253
rect 633270 651190 633726 651246
rect 633270 651183 633600 651190
rect 633270 650638 633726 650694
rect 633347 650521 633411 650638
rect 633539 650050 633603 650113
rect 633270 649994 633726 650050
rect 633539 649929 633603 649994
rect 633270 649350 633726 649406
rect 633443 649232 633507 649350
rect 633270 648762 633600 648769
rect 633270 648706 633726 648762
rect 633270 648699 633600 648706
rect 633270 648210 633600 648217
rect 633270 648154 633726 648210
rect 633270 648147 633600 648154
rect 633270 647566 633600 647573
rect 633270 647510 633726 647566
rect 633270 647503 633600 647510
rect 633270 646922 633600 646929
rect 633270 646866 633726 646922
rect 633270 646859 633600 646866
rect 633270 646314 633726 646370
rect 633270 645726 633600 645733
rect 633270 645670 633726 645726
rect 633270 645663 633600 645670
rect 633270 645026 633726 645082
rect 633270 644530 633600 644537
rect 633270 644474 633726 644530
rect 633270 644467 633600 644474
rect 633270 643886 633600 643893
rect 633270 643830 633726 643886
rect 633270 643823 633600 643830
rect 633270 643186 633726 643242
rect 633270 642634 633726 642690
rect 633270 642046 633600 642053
rect 633270 641990 633726 642046
rect 633270 641983 633600 641990
rect 633443 641402 633507 641519
rect 633270 641346 633726 641402
rect -400 628324 56 628380
rect -181 628207 -117 628324
rect -274 627736 56 627743
rect -400 627680 56 627736
rect -274 627673 56 627680
rect -400 627036 56 627092
rect -400 626484 56 626540
rect -274 625896 56 625903
rect -400 625840 56 625896
rect -274 625833 56 625840
rect -274 625252 56 625259
rect -400 625196 56 625252
rect -274 625189 56 625196
rect -400 624644 56 624700
rect -274 624056 56 624063
rect -400 624000 56 624056
rect -274 623993 56 624000
rect -400 623356 56 623412
rect -274 622860 56 622867
rect -400 622804 56 622860
rect -274 622797 56 622804
rect -274 622216 56 622223
rect -400 622160 56 622216
rect -274 622153 56 622160
rect -274 621572 56 621579
rect -400 621516 56 621572
rect -274 621509 56 621516
rect -274 621020 56 621027
rect -400 620964 56 621020
rect -274 620957 56 620964
rect -181 620376 -117 620494
rect -400 620320 56 620376
rect -277 619732 -213 619797
rect -400 619676 56 619732
rect -277 619613 -213 619676
rect -85 619088 -21 619205
rect -400 619032 56 619088
rect -274 618536 56 618543
rect -400 618480 56 618536
rect -274 618473 56 618480
rect -274 617892 56 617899
rect -400 617836 56 617892
rect -274 617829 56 617836
rect -274 617248 56 617255
rect -400 617192 56 617248
rect -274 617185 56 617192
rect -274 616696 56 616703
rect -400 616640 56 616696
rect -274 616633 56 616640
rect -181 616052 -117 616170
rect -400 615996 56 616052
rect -277 615408 -213 615464
rect -400 615352 56 615408
rect -277 615292 -213 615352
rect -274 614856 56 614863
rect -400 614800 56 614856
rect -274 614793 56 614800
rect -274 614212 56 614219
rect -400 614156 56 614212
rect -274 614149 56 614156
rect -274 613568 56 613575
rect -400 613512 56 613568
rect -274 613505 56 613512
rect -400 612960 56 613016
rect 633270 611510 633726 611566
rect 633270 611014 633600 611021
rect 633270 610958 633726 611014
rect 633270 610951 633600 610958
rect 633270 610370 633600 610377
rect 633270 610314 633726 610370
rect 633270 610307 633600 610314
rect 633270 609726 633600 609733
rect 633270 609670 633726 609726
rect 633270 609663 633600 609670
rect 633539 609174 633603 609234
rect 633270 609118 633726 609174
rect 633539 609062 633603 609118
rect 633270 608474 633726 608530
rect 633443 608356 633507 608474
rect 633270 607886 633600 607893
rect 633270 607830 633726 607886
rect 633270 607823 633600 607830
rect 633270 607334 633600 607341
rect 633270 607278 633726 607334
rect 633270 607271 633600 607278
rect 633270 606690 633600 606697
rect 633270 606634 633726 606690
rect 633270 606627 633600 606634
rect 633270 606046 633600 606053
rect 633270 605990 633726 606046
rect 633270 605983 633600 605990
rect 633270 605438 633726 605494
rect 633347 605321 633411 605438
rect 633539 604850 633603 604913
rect 633270 604794 633726 604850
rect 633539 604729 633603 604794
rect 633270 604150 633726 604206
rect 633443 604032 633507 604150
rect 633270 603562 633600 603569
rect 633270 603506 633726 603562
rect 633270 603499 633600 603506
rect 633270 603010 633600 603017
rect 633270 602954 633726 603010
rect 633270 602947 633600 602954
rect 633270 602366 633600 602373
rect 633270 602310 633726 602366
rect 633270 602303 633600 602310
rect 633270 601722 633600 601729
rect 633270 601666 633726 601722
rect 633270 601659 633600 601666
rect 633270 601114 633726 601170
rect 633270 600526 633600 600533
rect 633270 600470 633726 600526
rect 633270 600463 633600 600470
rect 633270 599826 633726 599882
rect 633270 599330 633600 599337
rect 633270 599274 633726 599330
rect 633270 599267 633600 599274
rect 633270 598686 633600 598693
rect 633270 598630 633726 598686
rect 633270 598623 633600 598630
rect 633270 597986 633726 598042
rect 633270 597434 633726 597490
rect 633270 596846 633600 596853
rect 633270 596790 633726 596846
rect 633270 596783 633600 596790
rect 633443 596202 633507 596319
rect 633270 596146 633726 596202
rect -400 585124 56 585180
rect -181 585007 -117 585124
rect -274 584536 56 584543
rect -400 584480 56 584536
rect -274 584473 56 584480
rect -400 583836 56 583892
rect -400 583284 56 583340
rect -274 582696 56 582703
rect -400 582640 56 582696
rect -274 582633 56 582640
rect -274 582052 56 582059
rect -400 581996 56 582052
rect -274 581989 56 581996
rect -400 581444 56 581500
rect -274 580856 56 580863
rect -400 580800 56 580856
rect -274 580793 56 580800
rect -400 580156 56 580212
rect -274 579660 56 579667
rect -400 579604 56 579660
rect -274 579597 56 579604
rect -274 579016 56 579023
rect -400 578960 56 579016
rect -274 578953 56 578960
rect -274 578372 56 578379
rect -400 578316 56 578372
rect -274 578309 56 578316
rect -274 577820 56 577827
rect -400 577764 56 577820
rect -274 577757 56 577764
rect -181 577176 -117 577294
rect -400 577120 56 577176
rect -277 576532 -213 576597
rect -400 576476 56 576532
rect -277 576413 -213 576476
rect -85 575888 -21 576005
rect -400 575832 56 575888
rect -274 575336 56 575343
rect -400 575280 56 575336
rect -274 575273 56 575280
rect -274 574692 56 574699
rect -400 574636 56 574692
rect -274 574629 56 574636
rect -274 574048 56 574055
rect -400 573992 56 574048
rect -274 573985 56 573992
rect -274 573496 56 573503
rect -400 573440 56 573496
rect -274 573433 56 573440
rect -181 572852 -117 572970
rect -400 572796 56 572852
rect -277 572208 -213 572264
rect -400 572152 56 572208
rect -277 572092 -213 572152
rect -274 571656 56 571663
rect -400 571600 56 571656
rect -274 571593 56 571600
rect -274 571012 56 571019
rect -400 570956 56 571012
rect -274 570949 56 570956
rect -274 570368 56 570375
rect -400 570312 56 570368
rect -274 570305 56 570312
rect -400 569760 56 569816
rect 633270 566510 633726 566566
rect 633270 566014 633600 566021
rect 633270 565958 633726 566014
rect 633270 565951 633600 565958
rect 633270 565370 633600 565377
rect 633270 565314 633726 565370
rect 633270 565307 633600 565314
rect 633270 564726 633600 564733
rect 633270 564670 633726 564726
rect 633270 564663 633600 564670
rect 633539 564174 633603 564234
rect 633270 564118 633726 564174
rect 633539 564062 633603 564118
rect 633270 563474 633726 563530
rect 633443 563356 633507 563474
rect 633270 562886 633600 562893
rect 633270 562830 633726 562886
rect 633270 562823 633600 562830
rect 633270 562334 633600 562341
rect 633270 562278 633726 562334
rect 633270 562271 633600 562278
rect 633270 561690 633600 561697
rect 633270 561634 633726 561690
rect 633270 561627 633600 561634
rect 633270 561046 633600 561053
rect 633270 560990 633726 561046
rect 633270 560983 633600 560990
rect 633270 560438 633726 560494
rect 633347 560321 633411 560438
rect 633539 559850 633603 559913
rect 633270 559794 633726 559850
rect 633539 559729 633603 559794
rect 633270 559150 633726 559206
rect 633443 559032 633507 559150
rect 633270 558562 633600 558569
rect 633270 558506 633726 558562
rect 633270 558499 633600 558506
rect 633270 558010 633600 558017
rect 633270 557954 633726 558010
rect 633270 557947 633600 557954
rect 633270 557366 633600 557373
rect 633270 557310 633726 557366
rect 633270 557303 633600 557310
rect 633270 556722 633600 556729
rect 633270 556666 633726 556722
rect 633270 556659 633600 556666
rect 633270 556114 633726 556170
rect 633270 555526 633600 555533
rect 633270 555470 633726 555526
rect 633270 555463 633600 555470
rect 633270 554826 633726 554882
rect 633270 554330 633600 554337
rect 633270 554274 633726 554330
rect 633270 554267 633600 554274
rect 633270 553686 633600 553693
rect 633270 553630 633726 553686
rect 633270 553623 633600 553630
rect 633270 552986 633726 553042
rect 633270 552434 633726 552490
rect 633270 551846 633600 551853
rect 633270 551790 633726 551846
rect 633270 551783 633600 551790
rect 633443 551202 633507 551319
rect 633270 551146 633726 551202
rect -400 541924 56 541980
rect -181 541807 -117 541924
rect -274 541336 56 541343
rect -400 541280 56 541336
rect -274 541273 56 541280
rect -400 540636 56 540692
rect -400 540084 56 540140
rect -274 539496 56 539503
rect -400 539440 56 539496
rect -274 539433 56 539440
rect -274 538852 56 538859
rect -400 538796 56 538852
rect -274 538789 56 538796
rect -400 538244 56 538300
rect -274 537656 56 537663
rect -400 537600 56 537656
rect -274 537593 56 537600
rect -400 536956 56 537012
rect -274 536460 56 536467
rect -400 536404 56 536460
rect -274 536397 56 536404
rect -274 535816 56 535823
rect -400 535760 56 535816
rect -274 535753 56 535760
rect -274 535172 56 535179
rect -400 535116 56 535172
rect -274 535109 56 535116
rect -274 534620 56 534627
rect -400 534564 56 534620
rect -274 534557 56 534564
rect -181 533976 -117 534094
rect -400 533920 56 533976
rect -277 533332 -213 533397
rect -400 533276 56 533332
rect -277 533213 -213 533276
rect -85 532688 -21 532805
rect -400 532632 56 532688
rect -274 532136 56 532143
rect -400 532080 56 532136
rect -274 532073 56 532080
rect -274 531492 56 531499
rect -400 531436 56 531492
rect -274 531429 56 531436
rect -274 530848 56 530855
rect -400 530792 56 530848
rect -274 530785 56 530792
rect -274 530296 56 530303
rect -400 530240 56 530296
rect -274 530233 56 530240
rect -181 529652 -117 529770
rect -400 529596 56 529652
rect -277 529008 -213 529064
rect -400 528952 56 529008
rect -277 528892 -213 528952
rect -274 528456 56 528463
rect -400 528400 56 528456
rect -274 528393 56 528400
rect -274 527812 56 527819
rect -400 527756 56 527812
rect -274 527749 56 527756
rect -274 527168 56 527175
rect -400 527112 56 527168
rect -274 527105 56 527112
rect -400 526560 56 526616
rect 633270 521310 633726 521366
rect 633270 520814 633600 520821
rect 633270 520758 633726 520814
rect 633270 520751 633600 520758
rect 633270 520170 633600 520177
rect 633270 520114 633726 520170
rect 633270 520107 633600 520114
rect 633270 519526 633600 519533
rect 633270 519470 633726 519526
rect 633270 519463 633600 519470
rect 633539 518974 633603 519034
rect 633270 518918 633726 518974
rect 633539 518862 633603 518918
rect 633270 518274 633726 518330
rect 633443 518156 633507 518274
rect 633270 517686 633600 517693
rect 633270 517630 633726 517686
rect 633270 517623 633600 517630
rect 633270 517134 633600 517141
rect 633270 517078 633726 517134
rect 633270 517071 633600 517078
rect 633270 516490 633600 516497
rect 633270 516434 633726 516490
rect 633270 516427 633600 516434
rect 633270 515846 633600 515853
rect 633270 515790 633726 515846
rect 633270 515783 633600 515790
rect 633270 515238 633726 515294
rect 633347 515121 633411 515238
rect 633539 514650 633603 514713
rect 633270 514594 633726 514650
rect 633539 514529 633603 514594
rect 633270 513950 633726 514006
rect 633443 513832 633507 513950
rect 633270 513362 633600 513369
rect 633270 513306 633726 513362
rect 633270 513299 633600 513306
rect 633270 512810 633600 512817
rect 633270 512754 633726 512810
rect 633270 512747 633600 512754
rect 633270 512166 633600 512173
rect 633270 512110 633726 512166
rect 633270 512103 633600 512110
rect 633270 511522 633600 511529
rect 633270 511466 633726 511522
rect 633270 511459 633600 511466
rect 633270 510914 633726 510970
rect 633270 510326 633600 510333
rect 633270 510270 633726 510326
rect 633270 510263 633600 510270
rect 633270 509626 633726 509682
rect 633270 509130 633600 509137
rect 633270 509074 633726 509130
rect 633270 509067 633600 509074
rect 633270 508486 633600 508493
rect 633270 508430 633726 508486
rect 633270 508423 633600 508430
rect 633270 507786 633726 507842
rect 633270 507234 633726 507290
rect 633270 506646 633600 506653
rect 633270 506590 633726 506646
rect 633270 506583 633600 506590
rect 633443 506002 633507 506119
rect 633270 505946 633726 506002
rect -400 498724 56 498780
rect -181 498607 -117 498724
rect -274 498136 56 498143
rect -400 498080 56 498136
rect -274 498073 56 498080
rect -400 497436 56 497492
rect -400 496884 56 496940
rect -274 496296 56 496303
rect -400 496240 56 496296
rect -274 496233 56 496240
rect -274 495652 56 495659
rect -400 495596 56 495652
rect -274 495589 56 495596
rect -400 495044 56 495100
rect -274 494456 56 494463
rect -400 494400 56 494456
rect -274 494393 56 494400
rect -400 493756 56 493812
rect -274 493260 56 493267
rect -400 493204 56 493260
rect -274 493197 56 493204
rect -274 492616 56 492623
rect -400 492560 56 492616
rect -274 492553 56 492560
rect -274 491972 56 491979
rect -400 491916 56 491972
rect -274 491909 56 491916
rect -274 491420 56 491427
rect -400 491364 56 491420
rect -274 491357 56 491364
rect -181 490776 -117 490894
rect -400 490720 56 490776
rect -277 490132 -213 490197
rect -400 490076 56 490132
rect -277 490013 -213 490076
rect -85 489488 -21 489605
rect -400 489432 56 489488
rect -274 488936 56 488943
rect -400 488880 56 488936
rect -274 488873 56 488880
rect -274 488292 56 488299
rect -400 488236 56 488292
rect -274 488229 56 488236
rect -274 487648 56 487655
rect -400 487592 56 487648
rect -274 487585 56 487592
rect -274 487096 56 487103
rect -400 487040 56 487096
rect -274 487033 56 487040
rect -181 486452 -117 486570
rect -400 486396 56 486452
rect -277 485808 -213 485864
rect -400 485752 56 485808
rect -277 485692 -213 485752
rect -274 485256 56 485263
rect -400 485200 56 485256
rect -274 485193 56 485200
rect -274 484612 56 484619
rect -400 484556 56 484612
rect -274 484549 56 484556
rect -274 483968 56 483975
rect -400 483912 56 483968
rect -274 483905 56 483912
rect -400 483360 56 483416
rect -400 371124 56 371180
rect -181 371007 -117 371124
rect -274 370536 56 370543
rect -400 370480 56 370536
rect -274 370473 56 370480
rect -400 369836 56 369892
rect -400 369284 56 369340
rect -274 368696 56 368703
rect -400 368640 56 368696
rect -274 368633 56 368640
rect -274 368052 56 368059
rect -400 367996 56 368052
rect -274 367989 56 367996
rect -400 367444 56 367500
rect -274 366856 56 366863
rect -400 366800 56 366856
rect -274 366793 56 366800
rect -400 366156 56 366212
rect -274 365660 56 365667
rect -400 365604 56 365660
rect -274 365597 56 365604
rect -274 365016 56 365023
rect -400 364960 56 365016
rect -274 364953 56 364960
rect -274 364372 56 364379
rect -400 364316 56 364372
rect -274 364309 56 364316
rect -274 363820 56 363827
rect -400 363764 56 363820
rect -274 363757 56 363764
rect -181 363176 -117 363294
rect -400 363120 56 363176
rect -277 362532 -213 362597
rect -400 362476 56 362532
rect -277 362413 -213 362476
rect -85 361888 -21 362005
rect -400 361832 56 361888
rect -274 361336 56 361343
rect -400 361280 56 361336
rect -274 361273 56 361280
rect -274 360692 56 360699
rect -400 360636 56 360692
rect -274 360629 56 360636
rect -274 360048 56 360055
rect -400 359992 56 360048
rect -274 359985 56 359992
rect -274 359496 56 359503
rect -400 359440 56 359496
rect -274 359433 56 359440
rect -181 358852 -117 358970
rect -400 358796 56 358852
rect -277 358208 -213 358264
rect -400 358152 56 358208
rect -277 358092 -213 358152
rect -274 357656 56 357663
rect -400 357600 56 357656
rect -274 357593 56 357600
rect -274 357012 56 357019
rect -400 356956 56 357012
rect -274 356949 56 356956
rect -274 356368 56 356375
rect -400 356312 56 356368
rect -274 356305 56 356312
rect -400 355760 56 355816
rect 633270 344110 633726 344166
rect 633270 343614 633600 343621
rect 633270 343558 633726 343614
rect 633270 343551 633600 343558
rect 633270 342970 633600 342977
rect 633270 342914 633726 342970
rect 633270 342907 633600 342914
rect 633270 342326 633600 342333
rect 633270 342270 633726 342326
rect 633270 342263 633600 342270
rect 633539 341774 633603 341834
rect 633270 341718 633726 341774
rect 633539 341662 633603 341718
rect 633270 341074 633726 341130
rect 633443 340956 633507 341074
rect 633270 340486 633600 340493
rect 633270 340430 633726 340486
rect 633270 340423 633600 340430
rect 633270 339934 633600 339941
rect 633270 339878 633726 339934
rect 633270 339871 633600 339878
rect 633270 339290 633600 339297
rect 633270 339234 633726 339290
rect 633270 339227 633600 339234
rect 633270 338646 633600 338653
rect 633270 338590 633726 338646
rect 633270 338583 633600 338590
rect 633270 338038 633726 338094
rect 633347 337921 633411 338038
rect 633539 337450 633603 337513
rect 633270 337394 633726 337450
rect 633539 337329 633603 337394
rect 633270 336750 633726 336806
rect 633443 336632 633507 336750
rect 633270 336162 633600 336169
rect 633270 336106 633726 336162
rect 633270 336099 633600 336106
rect 633270 335610 633600 335617
rect 633270 335554 633726 335610
rect 633270 335547 633600 335554
rect 633270 334966 633600 334973
rect 633270 334910 633726 334966
rect 633270 334903 633600 334910
rect 633270 334322 633600 334329
rect 633270 334266 633726 334322
rect 633270 334259 633600 334266
rect 633270 333714 633726 333770
rect 633270 333126 633600 333133
rect 633270 333070 633726 333126
rect 633270 333063 633600 333070
rect 633270 332426 633726 332482
rect 633270 331874 633726 331930
rect 633270 331286 633600 331293
rect 633270 331230 633726 331286
rect 633270 331223 633600 331230
rect 633270 330586 633726 330642
rect 633270 330034 633726 330090
rect 633270 329446 633600 329453
rect 633270 329390 633726 329446
rect 633270 329383 633600 329390
rect 633443 328802 633507 328919
rect 633270 328746 633726 328802
rect -400 327924 56 327980
rect -181 327807 -117 327924
rect -274 327336 56 327343
rect -400 327280 56 327336
rect -274 327273 56 327280
rect -400 326636 56 326692
rect -400 326084 56 326140
rect -274 325496 56 325503
rect -400 325440 56 325496
rect -274 325433 56 325440
rect -274 324852 56 324859
rect -400 324796 56 324852
rect -274 324789 56 324796
rect -400 324244 56 324300
rect -274 323656 56 323663
rect -400 323600 56 323656
rect -274 323593 56 323600
rect -400 322956 56 323012
rect -274 322460 56 322467
rect -400 322404 56 322460
rect -274 322397 56 322404
rect -274 321816 56 321823
rect -400 321760 56 321816
rect -274 321753 56 321760
rect -274 321172 56 321179
rect -400 321116 56 321172
rect -274 321109 56 321116
rect -274 320620 56 320627
rect -400 320564 56 320620
rect -274 320557 56 320564
rect -181 319976 -117 320094
rect -400 319920 56 319976
rect -277 319332 -213 319397
rect -400 319276 56 319332
rect -277 319213 -213 319276
rect -85 318688 -21 318805
rect -400 318632 56 318688
rect -274 318136 56 318143
rect -400 318080 56 318136
rect -274 318073 56 318080
rect -274 317492 56 317499
rect -400 317436 56 317492
rect -274 317429 56 317436
rect -274 316848 56 316855
rect -400 316792 56 316848
rect -274 316785 56 316792
rect -274 316296 56 316303
rect -400 316240 56 316296
rect -274 316233 56 316240
rect -181 315652 -117 315770
rect -400 315596 56 315652
rect -277 315008 -213 315064
rect -400 314952 56 315008
rect -277 314892 -213 314952
rect -274 314456 56 314463
rect -400 314400 56 314456
rect -274 314393 56 314400
rect -274 313812 56 313819
rect -400 313756 56 313812
rect -274 313749 56 313756
rect -274 313168 56 313175
rect -400 313112 56 313168
rect -274 313105 56 313112
rect -400 312560 56 312616
rect 633270 298910 633726 298966
rect 633270 298414 633600 298421
rect 633270 298358 633726 298414
rect 633270 298351 633600 298358
rect 633270 297770 633600 297777
rect 633270 297714 633726 297770
rect 633270 297707 633600 297714
rect 633270 297126 633600 297133
rect 633270 297070 633726 297126
rect 633270 297063 633600 297070
rect 633539 296574 633603 296634
rect 633270 296518 633726 296574
rect 633539 296462 633603 296518
rect 633270 295874 633726 295930
rect 633443 295756 633507 295874
rect 633270 295286 633600 295293
rect 633270 295230 633726 295286
rect 633270 295223 633600 295230
rect 633270 294734 633600 294741
rect 633270 294678 633726 294734
rect 633270 294671 633600 294678
rect 633270 294090 633600 294097
rect 633270 294034 633726 294090
rect 633270 294027 633600 294034
rect 633270 293446 633600 293453
rect 633270 293390 633726 293446
rect 633270 293383 633600 293390
rect 633270 292838 633726 292894
rect 633347 292721 633411 292838
rect 633539 292250 633603 292313
rect 633270 292194 633726 292250
rect 633539 292129 633603 292194
rect 633270 291550 633726 291606
rect 633443 291432 633507 291550
rect 633270 290962 633600 290969
rect 633270 290906 633726 290962
rect 633270 290899 633600 290906
rect 633270 290410 633600 290417
rect 633270 290354 633726 290410
rect 633270 290347 633600 290354
rect 633270 289766 633600 289773
rect 633270 289710 633726 289766
rect 633270 289703 633600 289710
rect 633270 289122 633600 289129
rect 633270 289066 633726 289122
rect 633270 289059 633600 289066
rect 633270 288514 633726 288570
rect 633270 287926 633600 287933
rect 633270 287870 633726 287926
rect 633270 287863 633600 287870
rect 633270 287226 633726 287282
rect 633270 286674 633726 286730
rect 633270 286086 633600 286093
rect 633270 286030 633726 286086
rect 633270 286023 633600 286030
rect 633270 285386 633726 285442
rect 633270 284834 633726 284890
rect -400 284724 56 284780
rect -181 284607 -117 284724
rect 633270 284246 633600 284253
rect 633270 284190 633726 284246
rect 633270 284183 633600 284190
rect -274 284136 56 284143
rect -400 284080 56 284136
rect -274 284073 56 284080
rect 633443 283602 633507 283719
rect 633270 283546 633726 283602
rect -400 283436 56 283492
rect -400 282884 56 282940
rect -274 282296 56 282303
rect -400 282240 56 282296
rect -274 282233 56 282240
rect -274 281652 56 281659
rect -400 281596 56 281652
rect -274 281589 56 281596
rect -400 281044 56 281100
rect -274 280456 56 280463
rect -400 280400 56 280456
rect -274 280393 56 280400
rect -400 279756 56 279812
rect -274 279260 56 279267
rect -400 279204 56 279260
rect -274 279197 56 279204
rect -274 278616 56 278623
rect -400 278560 56 278616
rect -274 278553 56 278560
rect -274 277972 56 277979
rect -400 277916 56 277972
rect -274 277909 56 277916
rect -274 277420 56 277427
rect -400 277364 56 277420
rect -274 277357 56 277364
rect -181 276776 -117 276894
rect -400 276720 56 276776
rect -277 276132 -213 276197
rect -400 276076 56 276132
rect -277 276013 -213 276076
rect -85 275488 -21 275605
rect -400 275432 56 275488
rect -274 274936 56 274943
rect -400 274880 56 274936
rect -274 274873 56 274880
rect -274 274292 56 274299
rect -400 274236 56 274292
rect -274 274229 56 274236
rect -274 273648 56 273655
rect -400 273592 56 273648
rect -274 273585 56 273592
rect -274 273096 56 273103
rect -400 273040 56 273096
rect -274 273033 56 273040
rect -181 272452 -117 272570
rect -400 272396 56 272452
rect -277 271808 -213 271864
rect -400 271752 56 271808
rect -277 271692 -213 271752
rect -274 271256 56 271263
rect -400 271200 56 271256
rect -274 271193 56 271200
rect -274 270612 56 270619
rect -400 270556 56 270612
rect -274 270549 56 270556
rect -274 269968 56 269975
rect -400 269912 56 269968
rect -274 269905 56 269912
rect -400 269360 56 269416
rect 633270 253910 633726 253966
rect 633270 253414 633600 253421
rect 633270 253358 633726 253414
rect 633270 253351 633600 253358
rect 633270 252770 633600 252777
rect 633270 252714 633726 252770
rect 633270 252707 633600 252714
rect 633270 252126 633600 252133
rect 633270 252070 633726 252126
rect 633270 252063 633600 252070
rect 633539 251574 633603 251634
rect 633270 251518 633726 251574
rect 633539 251462 633603 251518
rect 633270 250874 633726 250930
rect 633443 250756 633507 250874
rect 633270 250286 633600 250293
rect 633270 250230 633726 250286
rect 633270 250223 633600 250230
rect 633270 249734 633600 249741
rect 633270 249678 633726 249734
rect 633270 249671 633600 249678
rect 633270 249090 633600 249097
rect 633270 249034 633726 249090
rect 633270 249027 633600 249034
rect 633270 248446 633600 248453
rect 633270 248390 633726 248446
rect 633270 248383 633600 248390
rect 633270 247838 633726 247894
rect 633347 247721 633411 247838
rect 633539 247250 633603 247313
rect 633270 247194 633726 247250
rect 633539 247129 633603 247194
rect 633270 246550 633726 246606
rect 633443 246432 633507 246550
rect 633270 245962 633600 245969
rect 633270 245906 633726 245962
rect 633270 245899 633600 245906
rect 633270 245410 633600 245417
rect 633270 245354 633726 245410
rect 633270 245347 633600 245354
rect 633270 244766 633600 244773
rect 633270 244710 633726 244766
rect 633270 244703 633600 244710
rect 633270 244122 633600 244129
rect 633270 244066 633726 244122
rect 633270 244059 633600 244066
rect 633270 243514 633726 243570
rect 633270 242926 633600 242933
rect 633270 242870 633726 242926
rect 633270 242863 633600 242870
rect 633270 242226 633726 242282
rect 633270 241674 633726 241730
rect -400 241524 56 241580
rect -181 241407 -117 241524
rect 633270 241086 633600 241093
rect 633270 241030 633726 241086
rect 633270 241023 633600 241030
rect -274 240936 56 240943
rect -400 240880 56 240936
rect -274 240873 56 240880
rect 633270 240386 633726 240442
rect -400 240236 56 240292
rect 633270 239834 633726 239890
rect -400 239684 56 239740
rect 633270 239246 633600 239253
rect 633270 239190 633726 239246
rect 633270 239183 633600 239190
rect -274 239096 56 239103
rect -400 239040 56 239096
rect -274 239033 56 239040
rect 633443 238602 633507 238719
rect 633270 238546 633726 238602
rect -274 238452 56 238459
rect -400 238396 56 238452
rect -274 238389 56 238396
rect -400 237844 56 237900
rect -274 237256 56 237263
rect -400 237200 56 237256
rect -274 237193 56 237200
rect -400 236556 56 236612
rect -274 236060 56 236067
rect -400 236004 56 236060
rect -274 235997 56 236004
rect -274 235416 56 235423
rect -400 235360 56 235416
rect -274 235353 56 235360
rect -274 234772 56 234779
rect -400 234716 56 234772
rect -274 234709 56 234716
rect -274 234220 56 234227
rect -400 234164 56 234220
rect -274 234157 56 234164
rect -181 233576 -117 233694
rect -400 233520 56 233576
rect -277 232932 -213 232997
rect -400 232876 56 232932
rect -277 232813 -213 232876
rect -85 232288 -21 232405
rect -400 232232 56 232288
rect -274 231736 56 231743
rect -400 231680 56 231736
rect -274 231673 56 231680
rect -274 231092 56 231099
rect -400 231036 56 231092
rect -274 231029 56 231036
rect -274 230448 56 230455
rect -400 230392 56 230448
rect -274 230385 56 230392
rect -274 229896 56 229903
rect -400 229840 56 229896
rect -274 229833 56 229840
rect -181 229252 -117 229370
rect -400 229196 56 229252
rect -277 228608 -213 228664
rect -400 228552 56 228608
rect -277 228492 -213 228552
rect -274 228056 56 228063
rect -400 228000 56 228056
rect -274 227993 56 228000
rect -274 227412 56 227419
rect -400 227356 56 227412
rect -274 227349 56 227356
rect -274 226768 56 226775
rect -400 226712 56 226768
rect -274 226705 56 226712
rect -400 226160 56 226216
rect 633270 208910 633726 208966
rect 633270 208414 633600 208421
rect 633270 208358 633726 208414
rect 633270 208351 633600 208358
rect 633270 207770 633600 207777
rect 633270 207714 633726 207770
rect 633270 207707 633600 207714
rect 633270 207126 633600 207133
rect 633270 207070 633726 207126
rect 633270 207063 633600 207070
rect 633539 206574 633603 206634
rect 633270 206518 633726 206574
rect 633539 206462 633603 206518
rect 633270 205874 633726 205930
rect 633443 205756 633507 205874
rect 633270 205286 633600 205293
rect 633270 205230 633726 205286
rect 633270 205223 633600 205230
rect 633270 204734 633600 204741
rect 633270 204678 633726 204734
rect 633270 204671 633600 204678
rect 633270 204090 633600 204097
rect 633270 204034 633726 204090
rect 633270 204027 633600 204034
rect 633270 203446 633600 203453
rect 633270 203390 633726 203446
rect 633270 203383 633600 203390
rect 633270 202838 633726 202894
rect 633347 202721 633411 202838
rect 633539 202250 633603 202313
rect 633270 202194 633726 202250
rect 633539 202129 633603 202194
rect 633270 201550 633726 201606
rect 633443 201432 633507 201550
rect 633270 200962 633600 200969
rect 633270 200906 633726 200962
rect 633270 200899 633600 200906
rect 633270 200410 633600 200417
rect 633270 200354 633726 200410
rect 633270 200347 633600 200354
rect 633270 199766 633600 199773
rect 633270 199710 633726 199766
rect 633270 199703 633600 199710
rect 633270 199122 633600 199129
rect 633270 199066 633726 199122
rect 633270 199059 633600 199066
rect 633270 198514 633726 198570
rect -400 198324 56 198380
rect -181 198207 -117 198324
rect 633270 197926 633600 197933
rect 633270 197870 633726 197926
rect 633270 197863 633600 197870
rect -274 197736 56 197743
rect -400 197680 56 197736
rect -274 197673 56 197680
rect 633270 197226 633726 197282
rect -400 197036 56 197092
rect 633270 196674 633726 196730
rect -400 196484 56 196540
rect 633270 196086 633600 196093
rect 633270 196030 633726 196086
rect 633270 196023 633600 196030
rect -274 195896 56 195903
rect -400 195840 56 195896
rect -274 195833 56 195840
rect 633270 195386 633726 195442
rect -400 195196 56 195252
rect 633270 194834 633726 194890
rect -400 194644 56 194700
rect 633270 194246 633600 194253
rect 633270 194190 633726 194246
rect 633270 194183 633600 194190
rect -274 194056 56 194063
rect -400 194000 56 194056
rect -274 193993 56 194000
rect 633443 193602 633507 193719
rect 633270 193546 633726 193602
rect -400 193356 56 193412
rect -274 192860 56 192867
rect -400 192804 56 192860
rect -274 192797 56 192804
rect -274 192216 56 192223
rect -400 192160 56 192216
rect -274 192153 56 192160
rect -274 191572 56 191579
rect -400 191516 56 191572
rect -274 191509 56 191516
rect -274 191020 56 191027
rect -400 190964 56 191020
rect -274 190957 56 190964
rect -181 190376 -117 190494
rect -400 190320 56 190376
rect -277 189732 -213 189797
rect -400 189676 56 189732
rect -277 189613 -213 189676
rect -85 189088 -21 189205
rect -400 189032 56 189088
rect -274 188536 56 188543
rect -400 188480 56 188536
rect -274 188473 56 188480
rect -274 187892 56 187899
rect -400 187836 56 187892
rect -274 187829 56 187836
rect -274 187248 56 187255
rect -400 187192 56 187248
rect -274 187185 56 187192
rect -274 186696 56 186703
rect -400 186640 56 186696
rect -274 186633 56 186640
rect -181 186052 -117 186170
rect -400 185996 56 186052
rect -277 185408 -213 185464
rect -400 185352 56 185408
rect -277 185292 -213 185352
rect -274 184856 56 184863
rect -400 184800 56 184856
rect -274 184793 56 184800
rect -274 184212 56 184219
rect -400 184156 56 184212
rect -274 184149 56 184156
rect -274 183568 56 183575
rect -400 183512 56 183568
rect -274 183505 56 183512
rect -400 182960 56 183016
rect 633270 163710 633726 163766
rect 633270 163214 633600 163221
rect 633270 163158 633726 163214
rect 633270 163151 633600 163158
rect 633270 162570 633600 162577
rect 633270 162514 633726 162570
rect 633270 162507 633600 162514
rect 633270 161926 633600 161933
rect 633270 161870 633726 161926
rect 633270 161863 633600 161870
rect 633539 161374 633603 161434
rect 633270 161318 633726 161374
rect 633539 161262 633603 161318
rect 633270 160674 633726 160730
rect 633443 160556 633507 160674
rect 633270 160086 633600 160093
rect 633270 160030 633726 160086
rect 633270 160023 633600 160030
rect 633270 159534 633600 159541
rect 633270 159478 633726 159534
rect 633270 159471 633600 159478
rect 633270 158890 633600 158897
rect 633270 158834 633726 158890
rect 633270 158827 633600 158834
rect 633270 158246 633600 158253
rect 633270 158190 633726 158246
rect 633270 158183 633600 158190
rect 633270 157638 633726 157694
rect 633347 157521 633411 157638
rect 633539 157050 633603 157113
rect 633270 156994 633726 157050
rect 633539 156929 633603 156994
rect 633270 156350 633726 156406
rect 633443 156232 633507 156350
rect 633270 155762 633600 155769
rect 633270 155706 633726 155762
rect 633270 155699 633600 155706
rect 633270 155210 633600 155217
rect -400 155124 56 155180
rect 633270 155154 633726 155210
rect 633270 155147 633600 155154
rect -181 155007 -117 155124
rect 633270 154566 633600 154573
rect -274 154536 56 154543
rect -400 154480 56 154536
rect 633270 154510 633726 154566
rect 633270 154503 633600 154510
rect -274 154473 56 154480
rect 633270 153922 633600 153929
rect -400 153836 56 153892
rect 633270 153866 633726 153922
rect 633270 153859 633600 153866
rect -400 153284 56 153340
rect 633270 153314 633726 153370
rect 633270 152726 633600 152733
rect -274 152696 56 152703
rect -400 152640 56 152696
rect 633270 152670 633726 152726
rect 633270 152663 633600 152670
rect -274 152633 56 152640
rect -400 151996 56 152052
rect 633270 152026 633726 152082
rect -400 151444 56 151500
rect 633270 151474 633726 151530
rect 633270 150886 633600 150893
rect -274 150856 56 150863
rect -400 150800 56 150856
rect 633270 150830 633726 150886
rect 633270 150823 633600 150830
rect -274 150793 56 150800
rect -400 150156 56 150212
rect 633270 150186 633726 150242
rect -274 149660 56 149667
rect -400 149604 56 149660
rect 633270 149634 633726 149690
rect -274 149597 56 149604
rect 633270 149046 633600 149053
rect -274 149016 56 149023
rect -400 148960 56 149016
rect 633270 148990 633726 149046
rect 633270 148983 633600 148990
rect -274 148953 56 148960
rect 633443 148402 633507 148519
rect -274 148372 56 148379
rect -400 148316 56 148372
rect 633270 148346 633726 148402
rect -274 148309 56 148316
rect -274 147820 56 147827
rect -400 147764 56 147820
rect -274 147757 56 147764
rect -181 147176 -117 147294
rect -400 147120 56 147176
rect -277 146532 -213 146597
rect -400 146476 56 146532
rect -277 146413 -213 146476
rect -85 145888 -21 146005
rect -400 145832 56 145888
rect -274 145336 56 145343
rect -400 145280 56 145336
rect -274 145273 56 145280
rect -274 144692 56 144699
rect -400 144636 56 144692
rect -274 144629 56 144636
rect -274 144048 56 144055
rect -400 143992 56 144048
rect -274 143985 56 143992
rect -274 143496 56 143503
rect -400 143440 56 143496
rect -274 143433 56 143440
rect -181 142852 -117 142970
rect -400 142796 56 142852
rect -277 142208 -213 142264
rect -400 142152 56 142208
rect -277 142092 -213 142152
rect -274 141656 56 141663
rect -400 141600 56 141656
rect -274 141593 56 141600
rect -274 141012 56 141019
rect -400 140956 56 141012
rect -274 140949 56 140956
rect -274 140368 56 140375
rect -400 140312 56 140368
rect -274 140305 56 140312
rect -400 139760 56 139816
rect 633270 118710 633726 118766
rect 633270 118214 633600 118221
rect 633270 118158 633726 118214
rect 633270 118151 633600 118158
rect 633270 117570 633600 117577
rect 633270 117514 633726 117570
rect 633270 117507 633600 117514
rect 633270 116926 633600 116933
rect 633270 116870 633726 116926
rect 633270 116863 633600 116870
rect 633539 116374 633603 116434
rect 633270 116318 633726 116374
rect 633539 116262 633603 116318
rect 633270 115674 633726 115730
rect 633443 115556 633507 115674
rect 633270 115086 633600 115093
rect 633270 115030 633726 115086
rect 633270 115023 633600 115030
rect 633270 114534 633600 114541
rect 633270 114478 633726 114534
rect 633270 114471 633600 114478
rect 633270 113890 633600 113897
rect 633270 113834 633726 113890
rect 633270 113827 633600 113834
rect 633270 113246 633600 113253
rect 633270 113190 633726 113246
rect 633270 113183 633600 113190
rect 633270 112638 633726 112694
rect 633347 112521 633411 112638
rect 633539 112050 633603 112113
rect 633270 111994 633726 112050
rect 633539 111929 633603 111994
rect 633270 111350 633726 111406
rect 633443 111232 633507 111350
rect 633270 110762 633600 110769
rect 633270 110706 633726 110762
rect 633270 110699 633600 110706
rect 633270 110210 633600 110217
rect 633270 110154 633726 110210
rect 633270 110147 633600 110154
rect 633270 109566 633600 109573
rect 633270 109510 633726 109566
rect 633270 109503 633600 109510
rect 633270 108922 633600 108929
rect 633270 108866 633726 108922
rect 633270 108859 633600 108866
rect 633270 108314 633726 108370
rect 633270 107726 633600 107733
rect 633270 107670 633726 107726
rect 633270 107663 633600 107670
rect 633270 107026 633726 107082
rect 633270 106474 633726 106530
rect 633270 105886 633600 105893
rect 633270 105830 633726 105886
rect 633270 105823 633600 105830
rect 633270 105242 633600 105249
rect 633270 105186 633726 105242
rect 633270 105179 633600 105186
rect 633270 104634 633726 104690
rect 633270 104046 633600 104053
rect 633270 103990 633726 104046
rect 633270 103983 633600 103990
rect 633443 103402 633507 103519
rect 633270 103346 633726 103402
rect 633270 73510 633726 73566
rect 633270 73014 633600 73021
rect 633270 72958 633726 73014
rect 633270 72951 633600 72958
rect 633270 72370 633600 72377
rect 633270 72314 633726 72370
rect 633270 72307 633600 72314
rect 633270 71726 633600 71733
rect 633270 71670 633726 71726
rect 633270 71663 633600 71670
rect 633539 71174 633603 71234
rect 633270 71118 633726 71174
rect 633539 71062 633603 71118
rect 633270 70474 633726 70530
rect 633443 70356 633507 70474
rect 633270 69886 633600 69893
rect 633270 69830 633726 69886
rect 633270 69823 633600 69830
rect 633270 69334 633600 69341
rect 633270 69278 633726 69334
rect 633270 69271 633600 69278
rect 633270 68690 633600 68697
rect 633270 68634 633726 68690
rect 633270 68627 633600 68634
rect 633270 68046 633600 68053
rect 633270 67990 633726 68046
rect 633270 67983 633600 67990
rect 633270 67438 633726 67494
rect 633347 67321 633411 67438
rect 633539 66850 633603 66913
rect 633270 66794 633726 66850
rect 633539 66729 633603 66794
rect 633270 66150 633726 66206
rect 633443 66032 633507 66150
rect 633270 65562 633600 65569
rect 633270 65506 633726 65562
rect 633270 65499 633600 65506
rect 633270 65010 633600 65017
rect 633270 64954 633726 65010
rect 633270 64947 633600 64954
rect 633270 64366 633600 64373
rect 633270 64310 633726 64366
rect 633270 64303 633600 64310
rect 633270 63722 633600 63729
rect 633270 63666 633726 63722
rect 633270 63659 633600 63666
rect 633270 63114 633726 63170
rect 633270 62526 633600 62533
rect 633270 62470 633726 62526
rect 633270 62463 633600 62470
rect 633270 61826 633726 61882
rect 633270 61274 633726 61330
rect 633270 60686 633600 60693
rect 633270 60630 633726 60686
rect 633270 60623 633600 60630
rect 633270 59986 633726 60042
rect 633270 59434 633726 59490
rect 633270 58846 633600 58853
rect 633270 58790 633726 58846
rect 633270 58783 633600 58790
rect 633443 58202 633507 58319
rect 633270 58146 633726 58202
rect -400 53602 -292 53658
rect -400 53378 -292 53434
rect -400 53154 -292 53210
rect 99571 -90 99637 56
rect 99573 -400 99634 -90
rect 110164 -400 110220 56
rect 144546 -117 144602 56
rect 144546 -181 144719 -117
rect 144546 -400 144602 -181
rect 145190 -424 145246 56
rect 145834 -400 145890 56
rect 146386 -400 146442 56
rect 147030 -424 147086 56
rect 147674 -424 147730 56
rect 148226 -400 148282 56
rect 148870 -424 148926 56
rect 149514 -424 149570 56
rect 150066 -274 150123 56
rect 150066 -424 150122 -274
rect 150710 -424 150766 56
rect 151354 -424 151410 56
rect 151906 -424 151962 56
rect 152550 -117 152606 56
rect 152432 -181 152606 -117
rect 152550 -400 152606 -181
rect 153194 -213 153250 56
rect 153838 -21 153894 56
rect 153721 -85 153894 -21
rect 153129 -277 153313 -213
rect 153194 -400 153250 -277
rect 153838 -400 153894 -85
rect 154390 -424 154446 56
rect 155034 -424 155090 56
rect 155678 -424 155734 56
rect 156230 -424 156286 56
rect 156874 -117 156930 56
rect 156756 -181 156930 -117
rect 156874 -400 156930 -181
rect 157518 -213 157574 56
rect 157462 -277 157634 -213
rect 157518 -400 157574 -277
rect 158070 -424 158126 56
rect 158714 -424 158770 56
rect 159358 -424 159414 56
rect 159910 -424 159966 56
rect 160580 -400 160632 56
rect 163791 -400 163843 56
rect 253146 -117 253202 56
rect 253146 -181 253319 -117
rect 253146 -400 253202 -181
rect 253790 -424 253846 56
rect 254434 -400 254490 56
rect 254986 -400 255042 56
rect 255630 -424 255686 56
rect 256274 -424 256330 56
rect 256826 -400 256882 56
rect 257470 -424 257526 56
rect 258114 -424 258170 56
rect 258666 -424 258722 56
rect 259310 -424 259366 56
rect 259954 -424 260010 56
rect 260506 -424 260562 56
rect 261150 -117 261206 56
rect 261032 -181 261206 -117
rect 261150 -400 261206 -181
rect 261794 -213 261850 56
rect 262438 -21 262494 56
rect 262321 -85 262494 -21
rect 261729 -277 261913 -213
rect 261794 -400 261850 -277
rect 262438 -400 262494 -85
rect 262990 -424 263046 56
rect 263634 -424 263690 56
rect 264278 -424 264334 56
rect 264830 -424 264886 56
rect 265474 -117 265530 56
rect 265356 -181 265530 -117
rect 265474 -400 265530 -181
rect 266118 -213 266174 56
rect 266062 -277 266234 -213
rect 266118 -400 266174 -277
rect 266670 -424 266726 56
rect 267314 -424 267370 56
rect 267958 -424 268014 56
rect 268510 -424 268566 56
rect 268816 -363 268880 -311
rect 268824 -400 268872 -363
rect 269180 -400 269232 56
rect 273360 -400 273412 56
rect 307946 -117 308002 56
rect 307946 -181 308119 -117
rect 307946 -400 308002 -181
rect 308590 -424 308646 56
rect 309234 -400 309290 56
rect 309786 -400 309842 56
rect 310430 -424 310486 56
rect 311074 -424 311130 56
rect 311626 -400 311682 56
rect 312270 -424 312326 56
rect 312914 -424 312970 56
rect 313466 -424 313522 56
rect 314110 -424 314166 56
rect 314754 -424 314810 56
rect 315306 -424 315362 56
rect 315950 -117 316006 56
rect 315832 -181 316006 -117
rect 315950 -400 316006 -181
rect 316594 -213 316650 56
rect 317238 -21 317294 56
rect 317121 -85 317294 -21
rect 316529 -277 316713 -213
rect 316594 -400 316650 -277
rect 317238 -400 317294 -85
rect 317790 -424 317846 56
rect 318434 -424 318490 56
rect 319078 -424 319134 56
rect 319630 -424 319686 56
rect 320274 -117 320330 56
rect 320156 -181 320330 -117
rect 320274 -400 320330 -181
rect 320918 -213 320974 56
rect 320862 -277 321034 -213
rect 320918 -400 320974 -277
rect 321470 -424 321526 56
rect 322114 -424 322170 56
rect 322758 -424 322814 56
rect 323310 -424 323366 56
rect 323616 -363 323680 -311
rect 323624 -400 323672 -363
rect 323980 -400 324032 56
rect 328165 -400 328217 34
rect 362746 -117 362802 56
rect 362746 -181 362919 -117
rect 362746 -400 362802 -181
rect 363390 -424 363446 56
rect 364034 -400 364090 56
rect 364586 -400 364642 56
rect 365230 -424 365286 56
rect 365874 -424 365930 56
rect 366426 -400 366482 56
rect 367070 -424 367126 56
rect 367714 -424 367770 56
rect 368266 -424 368322 56
rect 368910 -424 368966 56
rect 369554 -424 369610 56
rect 370106 -424 370162 56
rect 370750 -117 370806 56
rect 370632 -181 370806 -117
rect 370750 -400 370806 -181
rect 371394 -213 371450 56
rect 372038 -21 372094 56
rect 371921 -85 372094 -21
rect 371329 -277 371513 -213
rect 371394 -400 371450 -277
rect 372038 -400 372094 -85
rect 372590 -424 372646 56
rect 373234 -424 373290 56
rect 373878 -424 373934 56
rect 374430 -424 374486 56
rect 375074 -117 375130 56
rect 374956 -181 375130 -117
rect 375074 -400 375130 -181
rect 375718 -213 375774 56
rect 375662 -277 375834 -213
rect 375718 -400 375774 -277
rect 376270 -424 376326 56
rect 376914 -424 376970 56
rect 377558 -424 377614 56
rect 378110 -424 378166 56
rect 378416 -363 378480 -311
rect 378424 -400 378472 -363
rect 378780 -400 378832 56
rect 382978 -400 383030 56
rect 417546 -117 417602 56
rect 417546 -181 417719 -117
rect 417546 -400 417602 -181
rect 418190 -424 418246 56
rect 418834 -400 418890 56
rect 419386 -400 419442 56
rect 420030 -424 420086 56
rect 420674 -424 420730 56
rect 421226 -400 421282 56
rect 421870 -424 421926 56
rect 422514 -424 422570 56
rect 423066 -424 423122 56
rect 423710 -424 423766 56
rect 424354 -424 424410 56
rect 424906 -424 424962 56
rect 425550 -117 425606 56
rect 425432 -181 425606 -117
rect 425550 -400 425606 -181
rect 426194 -213 426250 56
rect 426838 -21 426894 56
rect 426721 -85 426894 -21
rect 426129 -277 426313 -213
rect 426194 -400 426250 -277
rect 426838 -400 426894 -85
rect 427390 -424 427446 56
rect 428034 -424 428090 56
rect 428678 -424 428734 56
rect 429230 -424 429286 56
rect 429874 -117 429930 56
rect 429756 -181 429930 -117
rect 429874 -400 429930 -181
rect 430518 -213 430574 56
rect 430462 -277 430634 -213
rect 430518 -400 430574 -277
rect 431070 -424 431126 56
rect 431714 -424 431770 56
rect 432358 -424 432414 56
rect 432910 -424 432966 56
rect 433216 -363 433280 -311
rect 433224 -400 433272 -363
rect 433580 -400 433632 56
rect 437778 -400 437830 56
rect 472346 -117 472402 56
rect 472346 -181 472519 -117
rect 472346 -400 472402 -181
rect 472990 -424 473046 56
rect 473634 -400 473690 56
rect 474186 -400 474242 56
rect 474830 -424 474886 56
rect 475474 -424 475530 56
rect 476026 -400 476082 56
rect 476670 -424 476726 56
rect 477314 -424 477370 56
rect 477866 -424 477922 56
rect 478510 -424 478566 56
rect 479154 -424 479210 56
rect 479706 -424 479762 56
rect 480350 -117 480406 56
rect 480232 -181 480406 -117
rect 480350 -400 480406 -181
rect 480994 -213 481050 56
rect 481638 -21 481694 56
rect 481521 -85 481694 -21
rect 480929 -277 481113 -213
rect 480994 -400 481050 -277
rect 481638 -400 481694 -85
rect 482190 -424 482246 56
rect 482834 -424 482890 56
rect 483478 -424 483534 56
rect 484030 -424 484086 56
rect 484674 -117 484730 56
rect 484556 -181 484730 -117
rect 484674 -400 484730 -181
rect 485318 -213 485374 56
rect 485262 -277 485434 -213
rect 485318 -400 485374 -277
rect 485870 -424 485926 56
rect 486514 -424 486570 56
rect 487158 -424 487214 56
rect 487710 -424 487766 56
rect 488016 -363 488080 -311
rect 488024 -400 488072 -363
rect 488380 -400 488432 56
rect 492635 -400 492687 56
rect 605082 -260 605134 56
rect 605306 -260 605358 56
rect 605530 -260 605582 56
rect 605754 -260 605806 56
rect 605978 -260 606030 56
rect 606202 -260 606254 56
rect 606426 -260 606478 56
rect 606650 -260 606702 56
rect 606874 -260 606926 56
rect 607098 -260 607150 56
rect 607322 -260 607374 56
rect 607546 -260 607598 56
rect 607770 -260 607822 56
rect 607994 -260 608046 56
rect 608218 -260 608270 56
rect 608442 -260 608494 56
rect 608666 -260 608718 56
rect 608890 -260 608942 56
rect 609114 -260 609166 56
rect 609338 -260 609390 56
rect 609562 -260 609614 56
rect 609786 -260 609838 56
rect 610010 -260 610062 56
rect 610234 -260 610286 56
rect 610458 -260 610510 56
rect 610682 -260 610734 56
rect 610906 -260 610958 56
rect 611130 -260 611182 56
rect 611354 -260 611406 56
rect 611578 -260 611630 56
rect 611802 -260 611854 56
rect 612026 -260 612078 56
rect 605093 -400 605121 -260
rect 605317 -400 605345 -260
rect 605541 -400 605569 -260
rect 605765 -400 605793 -260
rect 605989 -400 606017 -260
rect 606213 -400 606241 -260
rect 606437 -400 606465 -260
rect 606661 -400 606689 -260
rect 606885 -400 606913 -260
rect 607109 -400 607137 -260
rect 607333 -400 607361 -260
rect 607557 -400 607585 -260
rect 607781 -400 607809 -260
rect 608005 -400 608033 -260
rect 608229 -400 608257 -260
rect 608453 -400 608481 -260
rect 608677 -400 608705 -260
rect 608901 -400 608929 -260
rect 609125 -400 609153 -260
rect 609349 -400 609377 -260
rect 609573 -400 609601 -260
rect 609797 -400 609825 -260
rect 610021 -400 610049 -260
rect 610245 -400 610273 -260
rect 610469 -400 610497 -260
rect 610693 -400 610721 -260
rect 610917 -400 610945 -260
rect 611141 -400 611169 -260
rect 611365 -400 611393 -260
rect 611589 -400 611617 -260
rect 611813 -400 611841 -260
rect 612037 -400 612065 -260
<< metal3 >>
rect 291362 953270 296142 953770
rect 301341 953270 306121 953770
rect 533562 953270 538342 953770
rect 543541 953270 548321 953770
rect 633270 929007 633726 929069
rect -424 927073 56 927143
rect 633270 927005 633726 927067
rect -424 925233 56 925303
rect 633270 925103 633750 925173
rect -424 924589 56 924659
rect 633270 924551 633750 924621
rect 633270 923907 633750 923977
rect -424 923393 56 923463
rect 633270 923263 633750 923333
rect -424 922749 57 922819
rect -424 922197 56 922267
rect -424 921553 56 921623
rect 633270 921423 633750 921493
rect -424 920909 56 920979
rect 633270 920871 633750 920941
rect -424 920357 56 920427
rect 633270 920227 633750 920297
rect 633270 919583 633750 919653
rect -424 917873 56 917943
rect -424 917229 56 917299
rect 633270 917099 633750 917169
rect -424 916585 56 916655
rect 633270 916547 633750 916617
rect -424 916033 56 916103
rect 633270 915903 633750 915973
rect 633270 915259 633750 915329
rect 633269 914707 633750 914777
rect -424 914193 56 914263
rect 633270 914063 633750 914133
rect -424 913549 56 913619
rect -424 912905 56 912975
rect 633270 912867 633750 912937
rect -424 912353 56 912423
rect 633270 912223 633750 912293
rect 633270 910383 633750 910453
rect -400 906644 56 906704
rect -400 904644 56 904704
rect -444 880014 56 884803
rect -444 875053 56 879715
rect 633270 875563 633770 880363
rect -444 869963 56 874763
rect 633270 870611 633770 875273
rect 633270 865523 633770 870312
rect -444 837741 56 842521
rect 633270 839007 633726 839069
rect 633270 837005 633726 837067
rect 633270 835903 633750 835973
rect 633270 835351 633750 835421
rect 633270 834707 633750 834777
rect 633270 834063 633750 834133
rect -444 827762 56 832542
rect 633270 832223 633750 832293
rect 633270 831671 633750 831741
rect 633270 831027 633750 831097
rect 633270 830383 633750 830453
rect 633270 827899 633750 827969
rect 633270 827347 633750 827417
rect 633270 826703 633750 826773
rect 633270 826059 633750 826129
rect 633269 825507 633750 825577
rect 633270 824863 633750 824933
rect 633270 823667 633750 823737
rect 633270 823023 633750 823093
rect 633270 821183 633750 821253
rect -444 795541 56 800321
rect -444 785562 56 790342
rect 633270 786384 633770 791164
rect 633270 776405 633770 781185
rect -424 757273 56 757343
rect -424 755433 56 755503
rect -424 754789 56 754859
rect -424 753593 56 753663
rect -424 752949 57 753019
rect -424 752397 56 752467
rect -424 751753 56 751823
rect -424 751109 56 751179
rect -424 750557 56 750627
rect 633270 750007 633726 750069
rect -424 748073 56 748143
rect 633270 748005 633726 748067
rect -424 747429 56 747499
rect -424 746785 56 746855
rect 633270 746703 633750 746773
rect -424 746233 56 746303
rect 633270 746151 633750 746221
rect 633270 745507 633750 745577
rect 633270 744863 633750 744933
rect -424 744393 56 744463
rect -424 743749 56 743819
rect -424 743105 56 743175
rect 633270 743023 633750 743093
rect -424 742553 56 742623
rect 633270 742471 633750 742541
rect 633270 741827 633750 741897
rect 633270 741183 633750 741253
rect 633270 738699 633750 738769
rect 633270 738147 633750 738217
rect 633270 737503 633750 737573
rect 633270 736859 633750 736929
rect -400 736644 56 736704
rect 633269 736307 633750 736377
rect 633270 735663 633750 735733
rect -400 734644 56 734704
rect 633270 734467 633750 734537
rect 633270 733823 633750 733893
rect 633270 731983 633750 732053
rect -424 714073 56 714143
rect -424 712233 56 712303
rect -424 711589 56 711659
rect -424 710393 56 710463
rect -424 709749 57 709819
rect -424 709197 56 709267
rect -424 708553 56 708623
rect -424 707909 56 707979
rect -424 707357 56 707427
rect 633270 705007 633726 705069
rect -424 704873 56 704943
rect -424 704229 56 704299
rect -424 703585 56 703655
rect -424 703033 56 703103
rect 633270 703005 633726 703067
rect 633270 701703 633750 701773
rect -424 701193 56 701263
rect 633270 701151 633750 701221
rect -424 700549 56 700619
rect 633270 700507 633750 700577
rect -424 699905 56 699975
rect 633270 699863 633750 699933
rect -424 699353 56 699423
rect 633270 698023 633750 698093
rect 633270 697471 633750 697541
rect 633270 696827 633750 696897
rect 633270 696183 633750 696253
rect -400 693644 56 693704
rect 633270 693699 633750 693769
rect 633270 693147 633750 693217
rect 633270 692503 633750 692573
rect 633270 691859 633750 691929
rect -400 691644 56 691704
rect 633269 691307 633750 691377
rect 633270 690663 633750 690733
rect 633270 689467 633750 689537
rect 633270 688823 633750 688893
rect 633270 686983 633750 687053
rect -424 670873 56 670943
rect -424 669033 56 669103
rect -424 668389 56 668459
rect -424 667193 56 667263
rect -424 666549 57 666619
rect -424 665997 56 666067
rect -424 665353 56 665423
rect -424 664709 56 664779
rect -424 664157 56 664227
rect -424 661673 56 661743
rect -424 661029 56 661099
rect -424 660385 56 660455
rect 633270 660007 633726 660069
rect -424 659833 56 659903
rect -424 657993 56 658063
rect 633270 658005 633726 658067
rect -424 657349 56 657419
rect -424 656705 56 656775
rect 633270 656703 633750 656773
rect -424 656153 56 656223
rect 633270 656151 633750 656221
rect 633270 655507 633750 655577
rect 633270 654863 633750 654933
rect 633270 653023 633750 653093
rect 633270 652471 633750 652541
rect 633270 651827 633750 651897
rect 633270 651183 633750 651253
rect -400 650644 56 650704
rect -400 648644 56 648704
rect 633270 648699 633750 648769
rect 633270 648147 633750 648217
rect 633270 647503 633750 647573
rect 633270 646859 633750 646929
rect 633269 646307 633750 646377
rect 633270 645663 633750 645733
rect 633270 644467 633750 644537
rect 633270 643823 633750 643893
rect 633270 641983 633750 642053
rect -424 627673 56 627743
rect -424 625833 56 625903
rect -424 625189 56 625259
rect -424 623993 56 624063
rect -424 623349 57 623419
rect -424 622797 56 622867
rect -424 622153 56 622223
rect -424 621509 56 621579
rect -424 620957 56 621027
rect -424 618473 56 618543
rect -424 617829 56 617899
rect -424 617185 56 617255
rect -424 616633 56 616703
rect 633270 615007 633726 615069
rect -424 614793 56 614863
rect -424 614149 56 614219
rect -424 613505 56 613575
rect -424 612953 56 613023
rect 633270 613005 633726 613067
rect 633270 611503 633750 611573
rect 633270 610951 633750 611021
rect 633270 610307 633750 610377
rect 633270 609663 633750 609733
rect 633270 607823 633750 607893
rect -400 607644 56 607704
rect 633270 607271 633750 607341
rect 633270 606627 633750 606697
rect 633270 605983 633750 606053
rect -400 605644 56 605704
rect 633270 603499 633750 603569
rect 633270 602947 633750 603017
rect 633270 602303 633750 602373
rect 633270 601659 633750 601729
rect 633269 601107 633750 601177
rect 633270 600463 633750 600533
rect 633270 599267 633750 599337
rect 633270 598623 633750 598693
rect 633270 596783 633750 596853
rect -424 584473 56 584543
rect -424 582633 56 582703
rect -424 581989 56 582059
rect -424 580793 56 580863
rect -424 580149 57 580219
rect -424 579597 56 579667
rect -424 578953 56 579023
rect -424 578309 56 578379
rect -424 577757 56 577827
rect -424 575273 56 575343
rect -424 574629 56 574699
rect -424 573985 56 574055
rect -424 573433 56 573503
rect -424 571593 56 571663
rect -424 570949 56 571019
rect -424 570305 56 570375
rect 633270 570007 633726 570069
rect -424 569753 56 569823
rect 633270 568005 633726 568067
rect 633270 566503 633750 566573
rect 633270 565951 633750 566021
rect 633270 565307 633750 565377
rect -400 564644 56 564704
rect 633270 564663 633750 564733
rect 633270 562823 633750 562893
rect -400 562644 56 562704
rect 633270 562271 633750 562341
rect 633270 561627 633750 561697
rect 633270 560983 633750 561053
rect 633270 558499 633750 558569
rect 633270 557947 633750 558017
rect 633270 557303 633750 557373
rect 633270 556659 633750 556729
rect 633269 556107 633750 556177
rect 633270 555463 633750 555533
rect 633270 554267 633750 554337
rect 633270 553623 633750 553693
rect 633270 551783 633750 551853
rect -424 541273 56 541343
rect -424 539433 56 539503
rect -424 538789 56 538859
rect -424 537593 56 537663
rect -424 536949 57 537019
rect -424 536397 56 536467
rect -424 535753 56 535823
rect -424 535109 56 535179
rect -424 534557 56 534627
rect -424 532073 56 532143
rect -424 531429 56 531499
rect -424 530785 56 530855
rect -424 530233 56 530303
rect -424 528393 56 528463
rect -424 527749 56 527819
rect -424 527105 56 527175
rect -424 526553 56 526623
rect 633270 525007 633726 525069
rect 633270 523005 633726 523067
rect -400 521644 56 521704
rect 633270 521303 633750 521373
rect 633270 520751 633750 520821
rect 633270 520107 633750 520177
rect -400 519644 56 519704
rect 633270 519463 633750 519533
rect 633270 517623 633750 517693
rect 633270 517071 633750 517141
rect 633270 516427 633750 516497
rect 633270 515783 633750 515853
rect 633270 513299 633750 513369
rect 633270 512747 633750 512817
rect 633270 512103 633750 512173
rect 633270 511459 633750 511529
rect 633269 510907 633750 510977
rect 633270 510263 633750 510333
rect 633270 509067 633750 509137
rect 633270 508423 633750 508493
rect 633270 506583 633750 506653
rect -424 498073 56 498143
rect -424 496233 56 496303
rect -424 495589 56 495659
rect -424 494393 56 494463
rect -424 493749 57 493819
rect -424 493197 56 493267
rect -424 492553 56 492623
rect -424 491909 56 491979
rect -424 491357 56 491427
rect -424 488873 56 488943
rect -424 488229 56 488299
rect -424 487585 56 487655
rect -424 487033 56 487103
rect -424 485193 56 485263
rect -424 484549 56 484619
rect -424 483905 56 483975
rect -424 483353 56 483423
rect -400 478644 56 478704
rect -400 476644 56 476704
rect 633270 471784 633770 476564
rect 633270 461805 633770 466585
rect -444 450941 56 455721
rect -444 440962 56 445742
rect 633270 427763 633770 432563
rect 633270 422812 633770 427463
rect 633270 417723 633770 422512
rect -444 408814 56 413603
rect -444 403863 56 408514
rect -444 398763 56 403563
rect 633270 383584 633770 388364
rect 633270 373605 633770 378385
rect -424 370473 56 370543
rect -424 368633 56 368703
rect -424 367989 56 368059
rect -424 366793 56 366863
rect -424 366149 57 366219
rect -424 365597 56 365667
rect -424 364953 56 365023
rect -424 364309 56 364379
rect -424 363757 56 363827
rect -424 361273 56 361343
rect -424 360629 56 360699
rect -424 359985 56 360055
rect -424 359433 56 359503
rect -424 357593 56 357663
rect -424 356949 56 357019
rect -424 356305 56 356375
rect -424 355753 56 355823
rect -400 349644 56 349704
rect 633270 348007 633726 348069
rect -400 347644 56 347704
rect 633270 346005 633726 346067
rect 633270 344103 633750 344173
rect 633270 343551 633750 343621
rect 633270 342907 633750 342977
rect 633270 342263 633750 342333
rect 633270 340423 633750 340493
rect 633270 339871 633750 339941
rect 633270 339227 633750 339297
rect 633270 338583 633750 338653
rect 633270 336099 633750 336169
rect 633270 335547 633750 335617
rect 633270 334903 633750 334973
rect 633270 334259 633750 334329
rect 633269 333707 633750 333777
rect 633270 333063 633750 333133
rect 633270 331867 633750 331937
rect 633270 331223 633750 331293
rect 633270 329383 633750 329453
rect -424 327273 56 327343
rect -424 325433 56 325503
rect -424 324789 56 324859
rect -424 323593 56 323663
rect -424 322949 57 323019
rect -424 322397 56 322467
rect -424 321753 56 321823
rect -424 321109 56 321179
rect -424 320557 56 320627
rect -424 318073 56 318143
rect -424 317429 56 317499
rect -424 316785 56 316855
rect -424 316233 56 316303
rect -424 314393 56 314463
rect -424 313749 56 313819
rect -424 313105 56 313175
rect -424 312553 56 312623
rect -400 306644 56 306704
rect -400 304644 56 304704
rect 633270 303007 633726 303069
rect 633270 301005 633726 301067
rect 633270 298903 633750 298973
rect 633270 298351 633750 298421
rect 633270 297707 633750 297777
rect 633270 297063 633750 297133
rect 633270 295223 633750 295293
rect 633270 294671 633750 294741
rect 633270 294027 633750 294097
rect 633270 293383 633750 293453
rect 633270 290899 633750 290969
rect 633270 290347 633750 290417
rect 633270 289703 633750 289773
rect 633270 289059 633750 289129
rect 633269 288507 633750 288577
rect 633270 287863 633750 287933
rect 633270 286667 633750 286737
rect 633270 286023 633750 286093
rect 633270 284183 633750 284253
rect -424 284073 56 284143
rect -424 282233 56 282303
rect -424 281589 56 281659
rect -424 280393 56 280463
rect -424 279749 57 279819
rect -424 279197 56 279267
rect -424 278553 56 278623
rect -424 277909 56 277979
rect -424 277357 56 277427
rect -424 274873 56 274943
rect -424 274229 56 274299
rect -424 273585 56 273655
rect -424 273033 56 273103
rect -424 271193 56 271263
rect -424 270549 56 270619
rect -424 269905 56 269975
rect -424 269353 56 269423
rect -400 263644 56 263704
rect -400 261644 56 261704
rect 633270 258007 633726 258069
rect 633270 256005 633726 256067
rect 633270 253903 633750 253973
rect 633270 253351 633750 253421
rect 633270 252707 633750 252777
rect 633270 252063 633750 252133
rect 633270 250223 633750 250293
rect 633270 249671 633750 249741
rect 633270 249027 633750 249097
rect 633270 248383 633750 248453
rect 633270 245899 633750 245969
rect 633270 245347 633750 245417
rect 633270 244703 633750 244773
rect 633270 244059 633750 244129
rect 633269 243507 633750 243577
rect 633270 242863 633750 242933
rect 633270 241667 633750 241737
rect 633270 241023 633750 241093
rect -424 240873 56 240943
rect 633270 239183 633750 239253
rect -424 239033 56 239103
rect -424 238389 56 238459
rect -424 237193 56 237263
rect -424 236549 57 236619
rect -424 235997 56 236067
rect -424 235353 56 235423
rect -424 234709 56 234779
rect -424 234157 56 234227
rect -424 231673 56 231743
rect -424 231029 56 231099
rect -424 230385 56 230455
rect -424 229833 56 229903
rect -424 227993 56 228063
rect -424 227349 56 227419
rect -424 226705 56 226775
rect -424 226153 56 226223
rect -400 220644 56 220704
rect -400 218644 56 218704
rect 633270 213007 633726 213069
rect 633270 211005 633726 211067
rect 633270 208903 633750 208973
rect 633270 208351 633750 208421
rect 633270 207707 633750 207777
rect 633270 207063 633750 207133
rect 633270 205223 633750 205293
rect 633270 204671 633750 204741
rect 633270 204027 633750 204097
rect 633270 203383 633750 203453
rect 633270 200899 633750 200969
rect 633270 200347 633750 200417
rect 633270 199703 633750 199773
rect 633270 199059 633750 199129
rect 633269 198507 633750 198577
rect 633270 197863 633750 197933
rect -424 197673 56 197744
rect 633270 196667 633750 196737
rect 633270 196023 633750 196093
rect -424 195833 56 195904
rect -424 195189 56 195260
rect 633270 194183 633750 194253
rect -424 193993 56 194064
rect -424 193419 56 193420
rect -424 193349 57 193419
rect -424 192797 56 192868
rect -424 192153 56 192224
rect -424 191509 56 191580
rect -424 190957 56 191028
rect -424 188473 56 188544
rect -424 187829 56 187900
rect -424 187185 56 187256
rect -424 186633 56 186704
rect -424 184793 56 184864
rect -424 184149 56 184220
rect -424 183505 56 183576
rect -424 182953 56 183024
rect -400 177644 56 177704
rect -400 175644 56 175704
rect 633270 168007 633726 168069
rect 633270 166005 633726 166067
rect 633270 163703 633750 163773
rect 633270 163151 633750 163221
rect 633270 162507 633750 162577
rect 633270 161863 633750 161933
rect 633270 160023 633750 160093
rect 633270 159471 633750 159541
rect 633270 158827 633750 158897
rect 633270 158183 633750 158253
rect 633270 155699 633750 155769
rect 633270 155147 633750 155217
rect -424 154473 56 154544
rect 633270 154503 633750 154573
rect 633270 153859 633750 153929
rect 633269 153307 633750 153377
rect -424 152633 56 152704
rect 633270 152663 633750 152733
rect -424 151989 56 152060
rect 633270 151467 633750 151537
rect -424 150793 56 150864
rect 633270 150823 633750 150893
rect -424 150219 56 150220
rect -424 150149 57 150219
rect -424 149597 56 149668
rect -424 148953 56 149024
rect 633270 148983 633750 149053
rect -424 148309 56 148380
rect -424 147757 56 147828
rect -424 145273 56 145344
rect -424 144629 56 144700
rect -424 143985 56 144056
rect -424 143433 56 143504
rect -424 141592 56 141663
rect -424 140949 56 141020
rect -424 140305 56 140376
rect -424 139753 56 139824
rect -400 134644 56 134704
rect -400 132644 56 132704
rect 633270 123007 633726 123069
rect 633270 121005 633726 121067
rect 633270 118703 633750 118773
rect 633270 118151 633750 118221
rect 633270 117507 633750 117577
rect 633270 116863 633750 116933
rect 633270 115023 633750 115093
rect 633270 114471 633750 114541
rect 633270 113827 633750 113897
rect 633270 113183 633750 113253
rect 633270 110699 633750 110769
rect 633270 110147 633750 110217
rect 633270 109503 633750 109573
rect 633270 108859 633750 108929
rect 633269 108307 633750 108377
rect 633270 107663 633750 107733
rect 633270 106467 633750 106537
rect 633270 105823 633750 105893
rect 633270 103983 633750 104053
rect -444 78141 56 82921
rect 633270 78007 633726 78069
rect 633270 76005 633726 76067
rect 633270 73503 633750 73573
rect 633270 72951 633750 73021
rect -444 68162 56 72942
rect 633270 72307 633750 72377
rect 633270 71663 633750 71733
rect 633270 69823 633750 69893
rect 633270 69271 633750 69341
rect 633270 68627 633750 68697
rect 633270 67983 633750 68053
rect 633270 65499 633750 65569
rect 633270 64947 633750 65017
rect 633270 64303 633750 64373
rect 633270 63659 633750 63729
rect 633269 63107 633750 63177
rect 633270 62463 633750 62533
rect 633270 61267 633750 61337
rect 633270 60623 633750 60693
rect 633270 58783 633750 58853
rect -400 53595 56 53665
rect -400 53372 56 53442
rect -400 53147 56 53217
rect -444 36014 56 40803
rect -444 25963 56 30763
rect 36805 -444 41585 56
rect 46784 -444 51564 57
rect 199283 -444 203912 56
rect 209163 -444 213963 56
rect 527005 -444 531785 56
rect 536984 -444 541764 56
rect 580805 -444 585585 56
rect 590784 -444 595564 56
<< comment >>
rect -400 953326 633726 953726
rect -400 0 0 953326
rect 633326 0 633726 953326
rect -400 -400 633726 0
<< labels >>
flabel metal2 485870 -424 485926 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[43]
port 290 nsew
flabel metal2 s 594004 953270 594060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[15]
port 450 nsew
flabel metal2 s 592716 953270 592772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[15]
port 538 nsew
flabel metal2 s 589680 953270 589736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[15]
port 494 nsew
flabel metal2 s 593360 953270 593416 953750 0 FreeSans 400 90 0 0 gpio_dm0[15]
port 582 nsew
flabel metal2 s 595200 953270 595256 953750 0 FreeSans 400 90 0 0 gpio_dm1[15]
port 626 nsew
flabel metal2 s 589036 953270 589092 953750 0 FreeSans 400 90 0 0 gpio_dm2[15]
port 670 nsew
flabel metal2 s 588392 953270 588448 953750 0 FreeSans 400 90 0 0 gpio_holdover[15]
port 406 nsew
flabel metal2 s 585356 953270 585412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[15]
port 274 nsew
flabel metal2 s 592164 953270 592220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[15]
port 230 nsew
flabel metal2 s 584712 953270 584768 953750 0 FreeSans 400 90 0 0 gpio_oeb[15]
port 186 nsew
flabel metal2 s 587840 953270 587896 953750 0 FreeSans 400 90 0 0 gpio_out[15]
port 142 nsew
flabel metal2 s 597040 953270 597096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[15]
port 362 nsew
flabel metal2 s 586000 953270 586056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[15]
port 318 nsew
flabel metal2 s 598880 953270 598936 953750 0 FreeSans 400 90 0 0 gpio_in[15]
port 714 nsew
flabel metal2 s 492204 953270 492260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[16]
port 449 nsew
flabel metal2 s 490916 953270 490972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[16]
port 537 nsew
flabel metal2 s 487880 953270 487936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[16]
port 493 nsew
flabel metal2 s 491560 953270 491616 953750 0 FreeSans 400 90 0 0 gpio_dm0[16]
port 581 nsew
flabel metal2 s 493400 953270 493456 953750 0 FreeSans 400 90 0 0 gpio_dm1[16]
port 625 nsew
flabel metal2 s 487236 953270 487292 953750 0 FreeSans 400 90 0 0 gpio_dm2[16]
port 669 nsew
flabel metal2 s 486592 953270 486648 953750 0 FreeSans 400 90 0 0 gpio_holdover[16]
port 405 nsew
flabel metal2 s 483556 953270 483612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[16]
port 273 nsew
flabel metal2 s 490364 953270 490420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[16]
port 229 nsew
flabel metal2 s 482912 953270 482968 953750 0 FreeSans 400 90 0 0 gpio_oeb[16]
port 185 nsew
flabel metal2 s 486040 953270 486096 953750 0 FreeSans 400 90 0 0 gpio_out[16]
port 141 nsew
flabel metal2 s 495240 953270 495296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[16]
port 361 nsew
flabel metal2 s 484200 953270 484256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[16]
port 317 nsew
flabel metal2 s 497080 953270 497136 953750 0 FreeSans 400 90 0 0 gpio_in[16]
port 713 nsew
flabel metal2 s 442000 953270 442056 953750 0 FreeSans 400 90 0 0 gpio_dm1[17]
port 624 nsew
flabel metal2 s 435836 953270 435892 953750 0 FreeSans 400 90 0 0 gpio_dm2[17]
port 668 nsew
flabel metal2 s 435192 953270 435248 953750 0 FreeSans 400 90 0 0 gpio_holdover[17]
port 404 nsew
flabel metal2 s 432156 953270 432212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[17]
port 272 nsew
flabel metal2 s 438964 953270 439020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[17]
port 228 nsew
flabel metal2 s 431512 953270 431568 953750 0 FreeSans 400 90 0 0 gpio_oeb[17]
port 184 nsew
flabel metal2 s 434640 953270 434696 953750 0 FreeSans 400 90 0 0 gpio_out[17]
port 140 nsew
flabel metal2 s 443840 953270 443896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[17]
port 360 nsew
flabel metal2 s 432800 953270 432856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[17]
port 316 nsew
flabel metal2 s 445680 953270 445736 953750 0 FreeSans 400 90 0 0 gpio_in[17]
port 712 nsew
flabel metal2 s 351804 953270 351860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[18]
port 447 nsew
flabel metal2 s 350516 953270 350572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[18]
port 535 nsew
flabel metal2 s 347480 953270 347536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[18]
port 491 nsew
flabel metal2 s 351160 953270 351216 953750 0 FreeSans 400 90 0 0 gpio_dm0[18]
port 579 nsew
flabel metal2 s 353000 953270 353056 953750 0 FreeSans 400 90 0 0 gpio_dm1[18]
port 623 nsew
flabel metal2 s 346836 953270 346892 953750 0 FreeSans 400 90 0 0 gpio_dm2[18]
port 667 nsew
flabel metal2 s 346192 953270 346248 953750 0 FreeSans 400 90 0 0 gpio_holdover[18]
port 403 nsew
flabel metal2 s 343156 953270 343212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[18]
port 271 nsew
flabel metal2 s 349964 953270 350020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[18]
port 227 nsew
flabel metal2 s 342512 953270 342568 953750 0 FreeSans 400 90 0 0 gpio_oeb[18]
port 183 nsew
flabel metal2 s 345640 953270 345696 953750 0 FreeSans 400 90 0 0 gpio_out[18]
port 139 nsew
flabel metal2 s 354840 953270 354896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[18]
port 359 nsew
flabel metal2 s 343800 953270 343856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[18]
port 315 nsew
flabel metal2 s 356680 953270 356736 953750 0 FreeSans 400 90 0 0 gpio_in[18]
port 711 nsew
flabel metal2 s 440804 953270 440860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[17]
port 448 nsew
flabel metal2 s 439516 953270 439572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[17]
port 536 nsew
flabel metal2 s 436480 953270 436536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[17]
port 492 nsew
flabel metal2 s 440160 953270 440216 953750 0 FreeSans 400 90 0 0 gpio_dm0[17]
port 580 nsew
flabel metal2 s 253040 953270 253096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[19]
port 358 nsew
flabel metal2 s 242000 953270 242056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[19]
port 314 nsew
flabel metal2 s 254880 953270 254936 953750 0 FreeSans 400 90 0 0 gpio_in[19]
port 710 nsew
flabel metal2 s 198404 953270 198460 953750 0 FreeSans 400 90 0 0 gpio_analog_en[20]
port 445 nsew
flabel metal2 s 197116 953270 197172 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[20]
port 533 nsew
flabel metal2 s 194080 953270 194136 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[20]
port 489 nsew
flabel metal2 s 197760 953270 197816 953750 0 FreeSans 400 90 0 0 gpio_dm0[20]
port 577 nsew
flabel metal2 s 199600 953270 199656 953750 0 FreeSans 400 90 0 0 gpio_dm1[20]
port 621 nsew
flabel metal2 s 193436 953270 193492 953750 0 FreeSans 400 90 0 0 gpio_dm2[20]
port 665 nsew
flabel metal2 s 192792 953270 192848 953750 0 FreeSans 400 90 0 0 gpio_holdover[20]
port 401 nsew
flabel metal2 s 189756 953270 189812 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[20]
port 269 nsew
flabel metal2 s 196564 953270 196620 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[20]
port 225 nsew
flabel metal2 s 189112 953270 189168 953750 0 FreeSans 400 90 0 0 gpio_oeb[20]
port 181 nsew
flabel metal2 s 192240 953270 192296 953750 0 FreeSans 400 90 0 0 gpio_out[20]
port 137 nsew
flabel metal2 s 201440 953270 201496 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[20]
port 357 nsew
flabel metal2 s 190400 953270 190456 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[20]
port 313 nsew
flabel metal2 s 203280 953270 203336 953750 0 FreeSans 400 90 0 0 gpio_in[20]
port 709 nsew
flabel metal2 s 250004 953270 250060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[19]
port 446 nsew
flabel metal2 s 248716 953270 248772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[19]
port 534 nsew
flabel metal2 s 245680 953270 245736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[19]
port 490 nsew
flabel metal2 s 249360 953270 249416 953750 0 FreeSans 400 90 0 0 gpio_dm0[19]
port 578 nsew
flabel metal2 s 251200 953270 251256 953750 0 FreeSans 400 90 0 0 gpio_dm1[19]
port 622 nsew
flabel metal2 s 245036 953270 245092 953750 0 FreeSans 400 90 0 0 gpio_dm2[19]
port 666 nsew
flabel metal2 s 244392 953270 244448 953750 0 FreeSans 400 90 0 0 gpio_holdover[19]
port 402 nsew
flabel metal2 s 241356 953270 241412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[19]
port 270 nsew
flabel metal2 s 248164 953270 248220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[19]
port 226 nsew
flabel metal2 s 240712 953270 240768 953750 0 FreeSans 400 90 0 0 gpio_oeb[19]
port 182 nsew
flabel metal2 s 243840 953270 243896 953750 0 FreeSans 400 90 0 0 gpio_out[19]
port 138 nsew
flabel metal2 s 151880 953270 151936 953750 0 FreeSans 400 90 0 0 gpio_in[21]
port 708 nsew
flabel metal2 s 95604 953270 95660 953750 0 FreeSans 400 90 0 0 gpio_analog_en[22]
port 443 nsew
flabel metal2 s 94316 953270 94372 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[22]
port 531 nsew
flabel metal2 s 91280 953270 91336 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[22]
port 487 nsew
flabel metal2 s 94960 953270 95016 953750 0 FreeSans 400 90 0 0 gpio_dm0[22]
port 575 nsew
flabel metal2 s 96800 953270 96856 953750 0 FreeSans 400 90 0 0 gpio_dm1[22]
port 619 nsew
flabel metal2 s 90636 953270 90692 953750 0 FreeSans 400 90 0 0 gpio_dm2[22]
port 663 nsew
flabel metal2 s 89992 953270 90048 953750 0 FreeSans 400 90 0 0 gpio_holdover[22]
port 399 nsew
flabel metal2 s 86956 953270 87012 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[22]
port 267 nsew
flabel metal2 s 93764 953270 93820 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[22]
port 223 nsew
flabel metal2 s 86312 953270 86368 953750 0 FreeSans 400 90 0 0 gpio_oeb[22]
port 179 nsew
flabel metal2 s 89440 953270 89496 953750 0 FreeSans 400 90 0 0 gpio_out[22]
port 135 nsew
flabel metal2 s 98640 953270 98696 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[22]
port 355 nsew
flabel metal2 s 87600 953270 87656 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[22]
port 311 nsew
flabel metal2 s 100480 953270 100536 953750 0 FreeSans 400 90 0 0 gpio_in[22]
port 707 nsew
flabel metal2 s 44204 953270 44260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[23]
port 442 nsew
flabel metal2 s 42916 953270 42972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[23]
port 530 nsew
flabel metal2 s 39880 953270 39936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[23]
port 486 nsew
flabel metal2 s 43560 953270 43616 953750 0 FreeSans 400 90 0 0 gpio_dm0[23]
port 574 nsew
flabel metal2 s 45400 953270 45456 953750 0 FreeSans 400 90 0 0 gpio_dm1[23]
port 618 nsew
flabel metal2 s 39236 953270 39292 953750 0 FreeSans 400 90 0 0 gpio_dm2[23]
port 662 nsew
flabel metal2 s 38592 953270 38648 953750 0 FreeSans 400 90 0 0 gpio_holdover[23]
port 398 nsew
flabel metal2 s 35556 953270 35612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[23]
port 266 nsew
flabel metal2 s 42364 953270 42420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[23]
port 222 nsew
flabel metal2 s 34912 953270 34968 953750 0 FreeSans 400 90 0 0 gpio_oeb[23]
port 178 nsew
flabel metal2 s 38040 953270 38096 953750 0 FreeSans 400 90 0 0 gpio_out[23]
port 134 nsew
flabel metal2 s 47240 953270 47296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[23]
port 354 nsew
flabel metal2 s 36200 953270 36256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[23]
port 310 nsew
flabel metal2 s 49080 953270 49136 953750 0 FreeSans 400 90 0 0 gpio_in[23]
port 706 nsew
flabel metal2 s 147004 953270 147060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[21]
port 444 nsew
flabel metal2 s 145716 953270 145772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[21]
port 532 nsew
flabel metal2 s 142680 953270 142736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[21]
port 488 nsew
flabel metal2 s 146360 953270 146416 953750 0 FreeSans 400 90 0 0 gpio_dm0[21]
port 576 nsew
flabel metal2 s 148200 953270 148256 953750 0 FreeSans 400 90 0 0 gpio_dm1[21]
port 620 nsew
flabel metal2 s 142036 953270 142092 953750 0 FreeSans 400 90 0 0 gpio_dm2[21]
port 664 nsew
flabel metal2 s 141392 953270 141448 953750 0 FreeSans 400 90 0 0 gpio_holdover[21]
port 400 nsew
flabel metal2 s 138356 953270 138412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[21]
port 268 nsew
flabel metal2 s 145164 953270 145220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[21]
port 224 nsew
flabel metal2 s 137712 953270 137768 953750 0 FreeSans 400 90 0 0 gpio_oeb[21]
port 180 nsew
flabel metal2 s 140840 953270 140896 953750 0 FreeSans 400 90 0 0 gpio_out[21]
port 136 nsew
flabel metal2 s 150040 953270 150096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[21]
port 356 nsew
flabel metal2 s 139000 953270 139056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[21]
port 312 nsew
flabel metal2 145190 -424 145246 56 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal2 147030 -424 147086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 148870 -424 148926 56 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 559 nsew
flabel metal2 150710 -424 150766 56 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 603 nsew
flabel metal2 151354 -424 151410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[38]
port 515 nsew
flabel metal2 150066 -424 150122 56 0 FreeSans 400 270 0 0 gpio_analog_en[38]
port 427 nsew
flabel metal2 151906 -424 151962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[38]
port 207 nsew
flabel metal2 154390 -424 154446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[38]
port 471 nsew
flabel metal2 155034 -424 155090 56 0 FreeSans 400 270 0 0 gpio_dm2[38]
port 647 nsew
flabel metal2 155678 -424 155734 56 0 FreeSans 400 270 0 0 gpio_holdover[38]
port 383 nsew
flabel metal2 156230 -424 156286 56 0 FreeSans 400 270 0 0 gpio_out[38]
port 119 nsew
flabel metal2 158070 -424 158126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[38]
port 295 nsew
flabel metal2 158714 -424 158770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[38]
port 251 nsew
flabel metal2 159358 -424 159414 56 0 FreeSans 400 270 0 0 gpio_oeb[38]
port 163 nsew
flabel metal2 253790 -424 253846 56 0 FreeSans 400 270 0 0 gpio_in[39]
port 690 nsew
flabel metal2 255630 -424 255686 56 0 FreeSans 400 270 0 0 gpio_slow_sel[39]
port 338 nsew
flabel metal2 257470 -424 257526 56 0 FreeSans 400 270 0 0 gpio_dm1[39]
port 602 nsew
flabel metal2 259310 -424 259366 56 0 FreeSans 400 270 0 0 gpio_dm0[39]
port 558 nsew
flabel metal2 259954 -424 260010 56 0 FreeSans 400 270 0 0 gpio_analog_pol[39]
port 514 nsew
flabel metal2 258666 -424 258722 56 0 FreeSans 400 270 0 0 gpio_analog_en[39]
port 426 nsew
flabel metal2 260506 -424 260562 56 0 FreeSans 400 270 0 0 gpio_inp_dis[39]
port 206 nsew
flabel metal2 262990 -424 263046 56 0 FreeSans 400 270 0 0 gpio_analog_sel[39]
port 470 nsew
flabel metal2 263634 -424 263690 56 0 FreeSans 400 270 0 0 gpio_dm2[39]
port 646 nsew
flabel metal2 264278 -424 264334 56 0 FreeSans 400 270 0 0 gpio_holdover[39]
port 382 nsew
flabel metal2 264830 -424 264886 56 0 FreeSans 400 270 0 0 gpio_out[39]
port 118 nsew
flabel metal2 266670 -424 266726 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[39]
port 294 nsew
flabel metal2 267314 -424 267370 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[39]
port 250 nsew
flabel metal2 267958 -424 268014 56 0 FreeSans 400 270 0 0 gpio_oeb[39]
port 162 nsew
flabel metal2 308590 -424 308646 56 0 FreeSans 400 270 0 0 gpio_in[40]
port 689 nsew
flabel metal2 310430 -424 310486 56 0 FreeSans 400 270 0 0 gpio_slow_sel[40]
port 337 nsew
flabel metal2 312270 -424 312326 56 0 FreeSans 400 270 0 0 gpio_dm1[40]
port 601 nsew
flabel metal2 314110 -424 314166 56 0 FreeSans 400 270 0 0 gpio_dm0[40]
port 557 nsew
flabel metal2 314754 -424 314810 56 0 FreeSans 400 270 0 0 gpio_analog_pol[40]
port 513 nsew
flabel metal2 313466 -424 313522 56 0 FreeSans 400 270 0 0 gpio_analog_en[40]
port 425 nsew
flabel metal2 315306 -424 315362 56 0 FreeSans 400 270 0 0 gpio_inp_dis[40]
port 205 nsew
flabel metal2 317790 -424 317846 56 0 FreeSans 400 270 0 0 gpio_analog_sel[40]
port 469 nsew
flabel metal2 318434 -424 318490 56 0 FreeSans 400 270 0 0 gpio_dm2[40]
port 645 nsew
flabel metal2 319078 -424 319134 56 0 FreeSans 400 270 0 0 gpio_holdover[40]
port 381 nsew
flabel metal2 319630 -424 319686 56 0 FreeSans 400 270 0 0 gpio_out[40]
port 117 nsew
flabel metal2 321470 -424 321526 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[40]
port 293 nsew
flabel metal2 322114 -424 322170 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[40]
port 249 nsew
flabel metal2 322758 -424 322814 56 0 FreeSans 400 270 0 0 gpio_oeb[40]
port 161 nsew
flabel metal2 363390 -424 363446 56 0 FreeSans 400 270 0 0 gpio_in[41]
port 688 nsew
flabel metal2 365230 -424 365286 56 0 FreeSans 400 270 0 0 gpio_slow_sel[41]
port 336 nsew
flabel metal2 367070 -424 367126 56 0 FreeSans 400 270 0 0 gpio_dm1[41]
port 600 nsew
flabel metal2 368910 -424 368966 56 0 FreeSans 400 270 0 0 gpio_dm0[41]
port 556 nsew
flabel metal2 369554 -424 369610 56 0 FreeSans 400 270 0 0 gpio_analog_pol[41]
port 512 nsew
flabel metal2 368266 -424 368322 56 0 FreeSans 400 270 0 0 gpio_analog_en[41]
port 424 nsew
flabel metal2 370106 -424 370162 56 0 FreeSans 400 270 0 0 gpio_inp_dis[41]
port 204 nsew
flabel metal2 372590 -424 372646 56 0 FreeSans 400 270 0 0 gpio_analog_sel[41]
port 468 nsew
flabel metal2 373234 -424 373290 56 0 FreeSans 400 270 0 0 gpio_dm2[41]
port 644 nsew
flabel metal2 373878 -424 373934 56 0 FreeSans 400 270 0 0 gpio_holdover[41]
port 380 nsew
flabel metal2 374430 -424 374486 56 0 FreeSans 400 270 0 0 gpio_out[41]
port 116 nsew
flabel metal2 376270 -424 376326 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[41]
port 292 nsew
flabel metal2 376914 -424 376970 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[41]
port 248 nsew
flabel metal2 377558 -424 377614 56 0 FreeSans 400 270 0 0 gpio_oeb[41]
port 160 nsew
flabel metal2 418190 -424 418246 56 0 FreeSans 400 270 0 0 gpio_in[42]
port 687 nsew
flabel metal2 420030 -424 420086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[42]
port 335 nsew
flabel metal2 421870 -424 421926 56 0 FreeSans 400 270 0 0 gpio_dm1[42]
port 599 nsew
flabel metal2 423710 -424 423766 56 0 FreeSans 400 270 0 0 gpio_dm0[42]
port 555 nsew
flabel metal2 424354 -424 424410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[42]
port 511 nsew
flabel metal2 423066 -424 423122 56 0 FreeSans 400 270 0 0 gpio_analog_en[42]
port 423 nsew
flabel metal2 424906 -424 424962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[42]
port 203 nsew
flabel metal2 427390 -424 427446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[42]
port 467 nsew
flabel metal2 428034 -424 428090 56 0 FreeSans 400 270 0 0 gpio_dm2[42]
port 643 nsew
flabel metal2 428678 -424 428734 56 0 FreeSans 400 270 0 0 gpio_holdover[42]
port 379 nsew
flabel metal2 429230 -424 429286 56 0 FreeSans 400 270 0 0 gpio_out[42]
port 115 nsew
flabel metal2 431070 -424 431126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[42]
port 291 nsew
flabel metal2 431714 -424 431770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[42]
port 247 nsew
flabel metal2 432358 -424 432414 56 0 FreeSans 400 270 0 0 gpio_oeb[42]
port 159 nsew
flabel metal2 472990 -424 473046 56 0 FreeSans 400 270 0 0 gpio_in[43]
port 686 nsew
flabel metal2 474830 -424 474886 56 0 FreeSans 400 270 0 0 gpio_slow_sel[43]
port 334 nsew
flabel metal2 476670 -424 476726 56 0 FreeSans 400 270 0 0 gpio_dm1[43]
port 598 nsew
flabel metal2 478510 -424 478566 56 0 FreeSans 400 270 0 0 gpio_dm0[43]
port 554 nsew
flabel metal2 479154 -424 479210 56 0 FreeSans 400 270 0 0 gpio_analog_pol[43]
port 510 nsew
flabel metal2 477866 -424 477922 56 0 FreeSans 400 270 0 0 gpio_analog_en[43]
port 422 nsew
flabel metal2 479706 -424 479762 56 0 FreeSans 400 270 0 0 gpio_inp_dis[43]
port 202 nsew
flabel metal2 482190 -424 482246 56 0 FreeSans 400 270 0 0 gpio_analog_sel[43]
port 466 nsew
flabel metal2 482834 -424 482890 56 0 FreeSans 400 270 0 0 gpio_dm2[43]
port 642 nsew
flabel metal2 483478 -424 483534 56 0 FreeSans 400 270 0 0 gpio_holdover[43]
port 378 nsew
flabel metal2 484030 -424 484086 56 0 FreeSans 400 270 0 0 gpio_out[43]
port 114 nsew
flabel metal2 486514 -424 486570 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[43]
port 246 nsew
flabel metal2 487158 -424 487214 56 0 FreeSans 400 270 0 0 gpio_oeb[43]
port 158 nsew
flabel metal2 s 584160 953270 584216 953750 0 FreeSans 400 90 0 0 gpio_in_h[15]
port 758 nsew
flabel metal2 s 482360 953270 482416 953750 0 FreeSans 400 90 0 0 gpio_in_h[16]
port 757 nsew
flabel metal2 s 430960 953270 431016 953750 0 FreeSans 400 90 0 0 gpio_in_h[17]
port 756 nsew
flabel metal2 s 341960 953270 342016 953750 0 FreeSans 400 90 0 0 gpio_in_h[18]
port 755 nsew
flabel metal2 s 240160 953270 240216 953750 0 FreeSans 400 90 0 0 gpio_in_h[19]
port 754 nsew
flabel metal2 s 188560 953270 188616 953750 0 FreeSans 400 90 0 0 gpio_in_h[20]
port 753 nsew
flabel metal2 s 137160 953270 137216 953750 0 FreeSans 400 90 0 0 gpio_in_h[21]
port 752 nsew
flabel metal2 s 85760 953270 85816 953750 0 FreeSans 400 90 0 0 gpio_in_h[22]
port 751 nsew
flabel metal2 s 34360 953270 34416 953750 0 FreeSans 400 90 0 0 gpio_in_h[23]
port 750 nsew
flabel metal2 s 159910 -424 159966 56 0 FreeSans 400 90 0 0 gpio_in_h[38]
port 735 nsew
flabel metal2 s 268510 -424 268566 56 0 FreeSans 400 90 0 0 gpio_in_h[39]
port 734 nsew
flabel metal2 s 323310 -424 323366 56 0 FreeSans 400 90 0 0 gpio_in_h[40]
port 733 nsew
flabel metal2 s 378110 -424 378166 56 0 FreeSans 400 90 0 0 gpio_in_h[41]
port 732 nsew
flabel metal2 s 432910 -424 432966 56 0 FreeSans 400 90 0 0 gpio_in_h[42]
port 731 nsew
flabel metal2 s 487710 -424 487766 56 0 FreeSans 400 90 0 0 gpio_in_h[43]
port 730 nsew
flabel metal2 s 596396 953270 596452 953750 0 FreeSans 400 90 0 0 analog_io[15]
port 890 nsew
flabel metal2 s 494596 953270 494652 953750 0 FreeSans 400 90 0 0 analog_io[16]
port 889 nsew
flabel metal2 s 443196 953270 443252 953750 0 FreeSans 400 90 0 0 analog_io[17]
port 888 nsew
flabel metal2 s 354196 953270 354252 953750 0 FreeSans 400 90 0 0 analog_io[18]
port 887 nsew
flabel metal2 s 252396 953270 252452 953750 0 FreeSans 400 90 0 0 analog_io[19]
port 886 nsew
flabel metal2 s 200796 953270 200852 953750 0 FreeSans 400 90 0 0 analog_io[20]
port 885 nsew
flabel metal2 s 149396 953270 149452 953750 0 FreeSans 400 90 0 0 analog_io[21]
port 884 nsew
flabel metal2 s 97996 953270 98052 953750 0 FreeSans 400 90 0 0 analog_io[22]
port 883 nsew
flabel metal2 s 46596 953270 46652 953750 0 FreeSans 400 90 0 0 analog_io[23]
port 882 nsew
flabel metal2 s 147674 -424 147730 56 0 FreeSans 400 90 0 0 analog_io[38]
port 867 nsew
flabel metal2 s 256274 -424 256330 56 0 FreeSans 400 90 0 0 analog_io[39]
port 866 nsew
flabel metal2 s 311074 -424 311130 56 0 FreeSans 400 90 0 0 analog_io[40]
port 865 nsew
flabel metal2 s 365874 -424 365930 56 0 FreeSans 400 90 0 0 analog_io[41]
port 864 nsew
flabel metal2 s 420674 -424 420730 56 0 FreeSans 400 90 0 0 analog_io[42]
port 863 nsew
flabel metal2 s 475474 -424 475530 56 0 FreeSans 400 90 0 0 analog_io[43]
port 862 nsew
flabel metal2 s 594556 953270 594612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[15]
port 934 nsew
flabel metal2 s 492756 953270 492812 953750 0 FreeSans 400 90 0 0 analog_noesd_io[16]
port 933 nsew
flabel metal2 s 441356 953270 441412 953750 0 FreeSans 400 90 0 0 analog_noesd_io[17]
port 932 nsew
flabel metal2 s 352356 953270 352412 953750 0 FreeSans 400 90 0 0 analog_noesd_io[18]
port 931 nsew
flabel metal2 s 250556 953270 250612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[19]
port 930 nsew
flabel metal2 s 198956 953270 199012 953750 0 FreeSans 400 90 0 0 analog_noesd_io[20]
port 929 nsew
flabel metal2 s 147556 953270 147612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[21]
port 928 nsew
flabel metal2 s 96156 953270 96212 953750 0 FreeSans 400 90 0 0 analog_noesd_io[22]
port 927 nsew
flabel metal2 s 44756 953270 44812 953750 0 FreeSans 400 90 0 0 analog_noesd_io[23]
port 926 nsew
flabel metal2 s 149514 -424 149570 56 0 FreeSans 400 90 0 0 analog_noesd_io[38]
port 911 nsew
flabel metal2 s 258114 -424 258170 56 0 FreeSans 400 90 0 0 analog_noesd_io[39]
port 910 nsew
flabel metal2 s 312914 -424 312970 56 0 FreeSans 400 90 0 0 analog_noesd_io[40]
port 909 nsew
flabel metal2 s 367714 -424 367770 56 0 FreeSans 400 90 0 0 analog_noesd_io[41]
port 908 nsew
flabel metal2 s 422514 -424 422570 56 0 FreeSans 400 90 0 0 analog_noesd_io[42]
port 907 nsew
flabel metal2 s 477314 -424 477370 56 0 FreeSans 400 90 0 0 analog_noesd_io[43]
port 906 nsew
flabel metal3 s -424 141592 56 141663 0 FreeSans 400 0 0 0 gpio_vtrip_sel[37]
port 296 nsew
flabel metal3 633270 422812 633770 427463 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 633270 427763 633770 432563 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 633270 417723 633770 422512 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633270 870611 633770 875273 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633270 875563 633770 880363 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633270 865523 633770 870312 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633270 786384 633770 791164 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 776405 633770 781185 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 471784 633770 476564 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 461805 633770 466585 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 383584 633770 388364 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 633270 373605 633770 378385 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 543541 953270 548321 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 533562 953270 538342 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 301341 953270 306121 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 291362 953270 296142 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -444 875053 56 879715 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 880014 56 884803 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 869963 56 874763 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 837741 56 842521 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 827762 56 832542 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 795541 56 800321 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -444 785562 56 790342 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -444 450941 56 455721 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 440962 56 445742 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 403863 56 408514 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 408814 56 413603 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 398763 56 403563 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 78141 56 82921 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 68162 56 72942 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 36014 56 40803 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 -444 25963 56 30763 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 46784 -443 51564 57 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 36805 -444 41585 56 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 209163 -444 213963 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 199283 -444 203912 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 536984 -444 541764 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 527005 -444 531785 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 580805 -444 585585 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 590784 -444 595564 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel comment s 107715 141850 108715 141850 0 FreeSans 1120000 60 0 0 example
flabel metal3 s 633270 736859 633750 736929 0 FreeSans 400 0 0 0 gpio_analog_en[12]
port 453 nsew
flabel metal3 s 633270 738147 633750 738217 0 FreeSans 400 0 0 0 gpio_analog_pol[12]
port 541 nsew
flabel metal3 s 633270 741183 633750 741253 0 FreeSans 400 0 0 0 gpio_analog_sel[12]
port 497 nsew
flabel metal3 s 633270 737503 633750 737573 0 FreeSans 400 0 0 0 gpio_dm0[12]
port 585 nsew
flabel metal3 s 633270 735663 633750 735733 0 FreeSans 400 0 0 0 gpio_dm1[12]
port 629 nsew
flabel metal3 s 633270 741827 633750 741897 0 FreeSans 400 0 0 0 gpio_dm2[12]
port 673 nsew
flabel metal3 s 633270 742471 633750 742541 0 FreeSans 400 0 0 0 gpio_holdover[12]
port 409 nsew
flabel metal3 s 633270 745507 633750 745577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[12]
port 277 nsew
flabel metal3 s 633270 738699 633750 738769 0 FreeSans 400 0 0 0 gpio_inp_dis[12]
port 233 nsew
flabel metal3 s 633270 746151 633750 746221 0 FreeSans 400 0 0 0 gpio_oeb[12]
port 189 nsew
flabel metal3 s 633270 743023 633750 743093 0 FreeSans 400 0 0 0 gpio_out[12]
port 145 nsew
flabel metal3 s 633270 733823 633750 733893 0 FreeSans 400 0 0 0 gpio_slow_sel[12]
port 365 nsew
flabel metal3 s 633270 744863 633750 744933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[12]
port 321 nsew
flabel metal3 s 633270 731983 633750 732053 0 FreeSans 400 0 0 0 gpio_in[12]
port 717 nsew
flabel metal3 s 633270 826059 633750 826129 0 FreeSans 400 0 0 0 gpio_analog_en[13]
port 452 nsew
flabel metal3 s 633270 827347 633750 827417 0 FreeSans 400 0 0 0 gpio_analog_pol[13]
port 540 nsew
flabel metal3 s 633270 830383 633750 830453 0 FreeSans 400 0 0 0 gpio_analog_sel[13]
port 496 nsew
flabel metal3 s 633270 826703 633750 826773 0 FreeSans 400 0 0 0 gpio_dm0[13]
port 584 nsew
flabel metal3 s 633270 824863 633750 824933 0 FreeSans 400 0 0 0 gpio_dm1[13]
port 628 nsew
flabel metal3 s 633270 831027 633750 831097 0 FreeSans 400 0 0 0 gpio_dm2[13]
port 672 nsew
flabel metal3 s 633270 831671 633750 831741 0 FreeSans 400 0 0 0 gpio_holdover[13]
port 408 nsew
flabel metal3 s 633270 834707 633750 834777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[13]
port 276 nsew
flabel metal3 s 633270 827899 633750 827969 0 FreeSans 400 0 0 0 gpio_inp_dis[13]
port 232 nsew
flabel metal3 s 633270 835351 633750 835421 0 FreeSans 400 0 0 0 gpio_oeb[13]
port 188 nsew
flabel metal3 s 633270 832223 633750 832293 0 FreeSans 400 0 0 0 gpio_out[13]
port 144 nsew
flabel metal3 s 633270 823023 633750 823093 0 FreeSans 400 0 0 0 gpio_slow_sel[13]
port 364 nsew
flabel metal3 s 633270 834063 633750 834133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[13]
port 320 nsew
flabel metal3 s 633270 821183 633750 821253 0 FreeSans 400 0 0 0 gpio_in[13]
port 716 nsew
flabel metal3 s 633270 915259 633750 915329 0 FreeSans 400 0 0 0 gpio_analog_en[14]
port 451 nsew
flabel metal3 s 633270 916547 633750 916617 0 FreeSans 400 0 0 0 gpio_analog_pol[14]
port 539 nsew
flabel metal3 s 633270 919583 633750 919653 0 FreeSans 400 0 0 0 gpio_analog_sel[14]
port 495 nsew
flabel metal3 s 633270 915903 633750 915973 0 FreeSans 400 0 0 0 gpio_dm0[14]
port 583 nsew
flabel metal3 s 633270 914063 633750 914133 0 FreeSans 400 0 0 0 gpio_dm1[14]
port 627 nsew
flabel metal3 s 633270 920227 633750 920297 0 FreeSans 400 0 0 0 gpio_dm2[14]
port 671 nsew
flabel metal3 s 633270 920871 633750 920941 0 FreeSans 400 0 0 0 gpio_holdover[14]
port 407 nsew
flabel metal3 s 633270 923907 633750 923977 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[14]
port 275 nsew
flabel metal3 s 633270 917099 633750 917169 0 FreeSans 400 0 0 0 gpio_inp_dis[14]
port 231 nsew
flabel metal3 s 633270 924551 633750 924621 0 FreeSans 400 0 0 0 gpio_oeb[14]
port 187 nsew
flabel metal3 s 633270 921423 633750 921493 0 FreeSans 400 0 0 0 gpio_out[14]
port 143 nsew
flabel metal3 s 633270 912223 633750 912293 0 FreeSans 400 0 0 0 gpio_slow_sel[14]
port 363 nsew
flabel metal3 s 633270 923263 633750 923333 0 FreeSans 400 0 0 0 gpio_vtrip_sel[14]
port 319 nsew
flabel metal3 s 633270 910383 633750 910453 0 FreeSans 400 0 0 0 gpio_in[14]
port 715 nsew
flabel metal3 s 633270 697471 633750 697541 0 FreeSans 400 0 0 0 gpio_holdover[11]
port 410 nsew
flabel metal3 s 633270 700507 633750 700577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[11]
port 278 nsew
flabel metal3 s 633270 693699 633750 693769 0 FreeSans 400 0 0 0 gpio_inp_dis[11]
port 234 nsew
flabel metal3 s 633270 701151 633750 701221 0 FreeSans 400 0 0 0 gpio_oeb[11]
port 190 nsew
flabel metal3 s 633270 698023 633750 698093 0 FreeSans 400 0 0 0 gpio_out[11]
port 146 nsew
flabel metal3 s 633270 688823 633750 688893 0 FreeSans 400 0 0 0 gpio_slow_sel[11]
port 366 nsew
flabel metal3 s 633270 699863 633750 699933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[11]
port 322 nsew
flabel metal3 s 633270 686983 633750 687053 0 FreeSans 400 0 0 0 gpio_in[11]
port 718 nsew
flabel metal3 s 633270 646859 633750 646929 0 FreeSans 400 0 0 0 gpio_analog_en[10]
port 455 nsew
flabel metal3 s 633270 648147 633750 648217 0 FreeSans 400 0 0 0 gpio_analog_pol[10]
port 543 nsew
flabel metal3 s 633270 651183 633750 651253 0 FreeSans 400 0 0 0 gpio_analog_sel[10]
port 499 nsew
flabel metal3 s 633270 647503 633750 647573 0 FreeSans 400 0 0 0 gpio_dm0[10]
port 587 nsew
flabel metal3 s 633270 645663 633750 645733 0 FreeSans 400 0 0 0 gpio_dm1[10]
port 631 nsew
flabel metal3 s 633270 651827 633750 651897 0 FreeSans 400 0 0 0 gpio_dm2[10]
port 675 nsew
flabel metal3 s 633270 652471 633750 652541 0 FreeSans 400 0 0 0 gpio_holdover[10]
port 411 nsew
flabel metal3 s 633270 655507 633750 655577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[10]
port 279 nsew
flabel metal3 s 633270 648699 633750 648769 0 FreeSans 400 0 0 0 gpio_inp_dis[10]
port 235 nsew
flabel metal3 s 633270 656151 633750 656221 0 FreeSans 400 0 0 0 gpio_oeb[10]
port 191 nsew
flabel metal3 s 633270 653023 633750 653093 0 FreeSans 400 0 0 0 gpio_out[10]
port 147 nsew
flabel metal3 s 633270 643823 633750 643893 0 FreeSans 400 0 0 0 gpio_slow_sel[10]
port 367 nsew
flabel metal3 s 633270 654863 633750 654933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[10]
port 323 nsew
flabel metal3 s 633270 641983 633750 642053 0 FreeSans 400 0 0 0 gpio_in[10]
port 719 nsew
flabel metal3 s 633270 511459 633750 511529 0 FreeSans 400 0 0 0 gpio_analog_en[7]
port 458 nsew
flabel metal3 s 633270 512747 633750 512817 0 FreeSans 400 0 0 0 gpio_analog_pol[7]
port 546 nsew
flabel metal3 s 633270 515783 633750 515853 0 FreeSans 400 0 0 0 gpio_analog_sel[7]
port 502 nsew
flabel metal3 s 633270 512103 633750 512173 0 FreeSans 400 0 0 0 gpio_dm0[7]
port 590 nsew
flabel metal3 s 633270 510263 633750 510333 0 FreeSans 400 0 0 0 gpio_dm1[7]
port 634 nsew
flabel metal3 s 633270 516427 633750 516497 0 FreeSans 400 0 0 0 gpio_dm2[7]
port 678 nsew
flabel metal3 s 633270 517071 633750 517141 0 FreeSans 400 0 0 0 gpio_holdover[7]
port 414 nsew
flabel metal3 s 633270 520107 633750 520177 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[7]
port 282 nsew
flabel metal3 s 633270 513299 633750 513369 0 FreeSans 400 0 0 0 gpio_inp_dis[7]
port 238 nsew
flabel metal3 s 633270 520751 633750 520821 0 FreeSans 400 0 0 0 gpio_oeb[7]
port 194 nsew
flabel metal3 s 633270 517623 633750 517693 0 FreeSans 400 0 0 0 gpio_out[7]
port 150 nsew
flabel metal3 s 633270 508423 633750 508493 0 FreeSans 400 0 0 0 gpio_slow_sel[7]
port 370 nsew
flabel metal3 s 633270 519463 633750 519533 0 FreeSans 400 0 0 0 gpio_vtrip_sel[7]
port 326 nsew
flabel metal3 s 633270 506583 633750 506653 0 FreeSans 400 0 0 0 gpio_in[7]
port 722 nsew
flabel metal3 s 633270 556659 633750 556729 0 FreeSans 400 0 0 0 gpio_analog_en[8]
port 457 nsew
flabel metal3 s 633270 557947 633750 558017 0 FreeSans 400 0 0 0 gpio_analog_pol[8]
port 545 nsew
flabel metal3 s 633270 560983 633750 561053 0 FreeSans 400 0 0 0 gpio_analog_sel[8]
port 501 nsew
flabel metal3 s 633270 557303 633750 557373 0 FreeSans 400 0 0 0 gpio_dm0[8]
port 589 nsew
flabel metal3 s 633270 555463 633750 555533 0 FreeSans 400 0 0 0 gpio_dm1[8]
port 633 nsew
flabel metal3 s 633270 561627 633750 561697 0 FreeSans 400 0 0 0 gpio_dm2[8]
port 677 nsew
flabel metal3 s 633270 562271 633750 562341 0 FreeSans 400 0 0 0 gpio_holdover[8]
port 413 nsew
flabel metal3 s 633270 565307 633750 565377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[8]
port 281 nsew
flabel metal3 s 633270 558499 633750 558569 0 FreeSans 400 0 0 0 gpio_inp_dis[8]
port 237 nsew
flabel metal3 s 633270 565951 633750 566021 0 FreeSans 400 0 0 0 gpio_oeb[8]
port 193 nsew
flabel metal3 s 633270 562823 633750 562893 0 FreeSans 400 0 0 0 gpio_out[8]
port 149 nsew
flabel metal3 s 633270 553623 633750 553693 0 FreeSans 400 0 0 0 gpio_slow_sel[8]
port 369 nsew
flabel metal3 s 633270 564663 633750 564733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[8]
port 325 nsew
flabel metal3 s 633270 551783 633750 551853 0 FreeSans 400 0 0 0 gpio_in[8]
port 721 nsew
flabel metal3 s 633270 601659 633750 601729 0 FreeSans 400 0 0 0 gpio_analog_en[9]
port 456 nsew
flabel metal3 s 633270 602947 633750 603017 0 FreeSans 400 0 0 0 gpio_analog_pol[9]
port 544 nsew
flabel metal3 s 633270 605983 633750 606053 0 FreeSans 400 0 0 0 gpio_analog_sel[9]
port 500 nsew
flabel metal3 s 633270 602303 633750 602373 0 FreeSans 400 0 0 0 gpio_dm0[9]
port 588 nsew
flabel metal3 s 633270 600463 633750 600533 0 FreeSans 400 0 0 0 gpio_dm1[9]
port 632 nsew
flabel metal3 s 633270 606627 633750 606697 0 FreeSans 400 0 0 0 gpio_dm2[9]
port 676 nsew
flabel metal3 s 633270 607271 633750 607341 0 FreeSans 400 0 0 0 gpio_holdover[9]
port 412 nsew
flabel metal3 s 633270 610307 633750 610377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[9]
port 280 nsew
flabel metal3 s 633270 603499 633750 603569 0 FreeSans 400 0 0 0 gpio_inp_dis[9]
port 236 nsew
flabel metal3 s 633270 610951 633750 611021 0 FreeSans 400 0 0 0 gpio_oeb[9]
port 192 nsew
flabel metal3 s 633270 607823 633750 607893 0 FreeSans 400 0 0 0 gpio_out[9]
port 148 nsew
flabel metal3 s 633270 598623 633750 598693 0 FreeSans 400 0 0 0 gpio_slow_sel[9]
port 368 nsew
flabel metal3 s 633270 609663 633750 609733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[9]
port 324 nsew
flabel metal3 s 633270 596783 633750 596853 0 FreeSans 400 0 0 0 gpio_in[9]
port 720 nsew
flabel metal3 s 633270 691859 633750 691929 0 FreeSans 400 0 0 0 gpio_analog_en[11]
port 454 nsew
flabel metal3 s 633270 693147 633750 693217 0 FreeSans 400 0 0 0 gpio_analog_pol[11]
port 542 nsew
flabel metal3 s 633270 696183 633750 696253 0 FreeSans 400 0 0 0 gpio_analog_sel[11]
port 498 nsew
flabel metal3 s 633270 692503 633750 692573 0 FreeSans 400 0 0 0 gpio_dm0[11]
port 586 nsew
flabel metal3 s 633270 690663 633750 690733 0 FreeSans 400 0 0 0 gpio_dm1[11]
port 630 nsew
flabel metal3 s 633270 696827 633750 696897 0 FreeSans 400 0 0 0 gpio_dm2[11]
port 674 nsew
flabel metal3 s 633270 244059 633750 244129 0 FreeSans 400 0 0 0 gpio_analog_en[4]
port 461 nsew
flabel metal3 s 633270 245347 633750 245417 0 FreeSans 400 0 0 0 gpio_analog_pol[4]
port 549 nsew
flabel metal3 s 633270 248383 633750 248453 0 FreeSans 400 0 0 0 gpio_analog_sel[4]
port 505 nsew
flabel metal3 s 633270 244703 633750 244773 0 FreeSans 400 0 0 0 gpio_dm0[4]
port 593 nsew
flabel metal3 s 633270 242863 633750 242933 0 FreeSans 400 0 0 0 gpio_dm1[4]
port 637 nsew
flabel metal3 s 633270 249027 633750 249097 0 FreeSans 400 0 0 0 gpio_dm2[4]
port 681 nsew
flabel metal3 s 633270 249671 633750 249741 0 FreeSans 400 0 0 0 gpio_holdover[4]
port 417 nsew
flabel metal3 s 633270 252707 633750 252777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[4]
port 285 nsew
flabel metal3 s 633270 245899 633750 245969 0 FreeSans 400 0 0 0 gpio_inp_dis[4]
port 241 nsew
flabel metal3 s 633270 253351 633750 253421 0 FreeSans 400 0 0 0 gpio_oeb[4]
port 197 nsew
flabel metal3 s 633270 250223 633750 250293 0 FreeSans 400 0 0 0 gpio_out[4]
port 153 nsew
flabel metal3 s 633270 241023 633750 241093 0 FreeSans 400 0 0 0 gpio_slow_sel[4]
port 373 nsew
flabel metal3 s 633270 252063 633750 252133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[4]
port 329 nsew
flabel metal3 s 633270 239183 633750 239253 0 FreeSans 400 0 0 0 gpio_in[4]
port 725 nsew
flabel metal3 s 633270 289059 633750 289129 0 FreeSans 400 0 0 0 gpio_analog_en[5]
port 460 nsew
flabel metal3 s 633270 290347 633750 290417 0 FreeSans 400 0 0 0 gpio_analog_pol[5]
port 548 nsew
flabel metal3 s 633270 293383 633750 293453 0 FreeSans 400 0 0 0 gpio_analog_sel[5]
port 504 nsew
flabel metal3 s 633270 289703 633750 289773 0 FreeSans 400 0 0 0 gpio_dm0[5]
port 592 nsew
flabel metal3 s 633270 287863 633750 287933 0 FreeSans 400 0 0 0 gpio_dm1[5]
port 636 nsew
flabel metal3 s 633270 294027 633750 294097 0 FreeSans 400 0 0 0 gpio_dm2[5]
port 680 nsew
flabel metal3 s 633270 294671 633750 294741 0 FreeSans 400 0 0 0 gpio_holdover[5]
port 416 nsew
flabel metal3 s 633270 297707 633750 297777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[5]
port 284 nsew
flabel metal3 s 633270 290899 633750 290969 0 FreeSans 400 0 0 0 gpio_inp_dis[5]
port 240 nsew
flabel metal3 s 633270 298351 633750 298421 0 FreeSans 400 0 0 0 gpio_oeb[5]
port 196 nsew
flabel metal3 s 633270 295223 633750 295293 0 FreeSans 400 0 0 0 gpio_out[5]
port 152 nsew
flabel metal3 s 633270 286023 633750 286093 0 FreeSans 400 0 0 0 gpio_slow_sel[5]
port 372 nsew
flabel metal3 s 633270 297063 633750 297133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[5]
port 328 nsew
flabel metal3 s 633270 284183 633750 284253 0 FreeSans 400 0 0 0 gpio_in[5]
port 724 nsew
flabel metal3 s 633270 334259 633750 334329 0 FreeSans 400 0 0 0 gpio_analog_en[6]
port 459 nsew
flabel metal3 s 633270 335547 633750 335617 0 FreeSans 400 0 0 0 gpio_analog_pol[6]
port 547 nsew
flabel metal3 s 633270 338583 633750 338653 0 FreeSans 400 0 0 0 gpio_analog_sel[6]
port 503 nsew
flabel metal3 s 633270 334903 633750 334973 0 FreeSans 400 0 0 0 gpio_dm0[6]
port 591 nsew
flabel metal3 s 633270 333063 633750 333133 0 FreeSans 400 0 0 0 gpio_dm1[6]
port 635 nsew
flabel metal3 s 633270 339227 633750 339297 0 FreeSans 400 0 0 0 gpio_dm2[6]
port 679 nsew
flabel metal3 s 633270 339871 633750 339941 0 FreeSans 400 0 0 0 gpio_holdover[6]
port 415 nsew
flabel metal3 s 633270 342907 633750 342977 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[6]
port 283 nsew
flabel metal3 s 633270 336099 633750 336169 0 FreeSans 400 0 0 0 gpio_inp_dis[6]
port 239 nsew
flabel metal3 s 633270 343551 633750 343621 0 FreeSans 400 0 0 0 gpio_oeb[6]
port 195 nsew
flabel metal3 s 633270 340423 633750 340493 0 FreeSans 400 0 0 0 gpio_out[6]
port 151 nsew
flabel metal3 s 633270 331223 633750 331293 0 FreeSans 400 0 0 0 gpio_slow_sel[6]
port 371 nsew
flabel metal3 s 633270 342263 633750 342333 0 FreeSans 400 0 0 0 gpio_vtrip_sel[6]
port 327 nsew
flabel metal3 s 633270 329383 633750 329453 0 FreeSans 400 0 0 0 gpio_in[6]
port 723 nsew
flabel metal3 s 633270 108859 633750 108929 0 FreeSans 400 0 0 0 gpio_analog_en[1]
port 464 nsew
flabel metal3 s 633270 110147 633750 110217 0 FreeSans 400 0 0 0 gpio_analog_pol[1]
port 552 nsew
flabel metal3 s 633270 113183 633750 113253 0 FreeSans 400 0 0 0 gpio_analog_sel[1]
port 508 nsew
flabel metal3 s 633270 109503 633750 109573 0 FreeSans 400 0 0 0 gpio_dm0[1]
port 596 nsew
flabel metal3 s 633270 107663 633750 107733 0 FreeSans 400 0 0 0 gpio_dm1[1]
port 640 nsew
flabel metal3 s 633270 113827 633750 113897 0 FreeSans 400 0 0 0 gpio_dm2[1]
port 684 nsew
flabel metal3 s 633270 114471 633750 114541 0 FreeSans 400 0 0 0 gpio_holdover[1]
port 420 nsew
flabel metal3 s 633270 117507 633750 117577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[1]
port 288 nsew
flabel metal3 s 633270 110699 633750 110769 0 FreeSans 400 0 0 0 gpio_inp_dis[1]
port 244 nsew
flabel metal3 s 633270 118151 633750 118221 0 FreeSans 400 0 0 0 gpio_oeb[1]
port 200 nsew
flabel metal3 s 633270 115023 633750 115093 0 FreeSans 400 0 0 0 gpio_out[1]
port 156 nsew
flabel metal3 s 633270 105823 633750 105893 0 FreeSans 400 0 0 0 gpio_slow_sel[1]
port 376 nsew
flabel metal3 s 633270 116863 633750 116933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[1]
port 332 nsew
flabel metal3 s 633270 103983 633750 104053 0 FreeSans 400 0 0 0 gpio_in[1]
port 728 nsew
flabel metal3 s 633270 153859 633750 153929 0 FreeSans 400 0 0 0 gpio_analog_en[2]
port 463 nsew
flabel metal3 s 633270 155147 633750 155217 0 FreeSans 400 0 0 0 gpio_analog_pol[2]
port 551 nsew
flabel metal3 s 633270 158183 633750 158253 0 FreeSans 400 0 0 0 gpio_analog_sel[2]
port 507 nsew
flabel metal3 s 633270 154503 633750 154573 0 FreeSans 400 0 0 0 gpio_dm0[2]
port 595 nsew
flabel metal3 s 633270 152663 633750 152733 0 FreeSans 400 0 0 0 gpio_dm1[2]
port 639 nsew
flabel metal3 s 633270 158827 633750 158897 0 FreeSans 400 0 0 0 gpio_dm2[2]
port 683 nsew
flabel metal3 s 633270 159471 633750 159541 0 FreeSans 400 0 0 0 gpio_holdover[2]
port 419 nsew
flabel metal3 s 633270 162507 633750 162577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[2]
port 287 nsew
flabel metal3 s 633270 155699 633750 155769 0 FreeSans 400 0 0 0 gpio_inp_dis[2]
port 243 nsew
flabel metal3 s 633270 163151 633750 163221 0 FreeSans 400 0 0 0 gpio_oeb[2]
port 199 nsew
flabel metal3 s 633270 160023 633750 160093 0 FreeSans 400 0 0 0 gpio_out[2]
port 155 nsew
flabel metal3 s 633270 150823 633750 150893 0 FreeSans 400 0 0 0 gpio_slow_sel[2]
port 375 nsew
flabel metal3 s 633270 161863 633750 161933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[2]
port 331 nsew
flabel metal3 s 633270 148983 633750 149053 0 FreeSans 400 0 0 0 gpio_in[2]
port 727 nsew
flabel metal3 s 633270 199059 633750 199129 0 FreeSans 400 0 0 0 gpio_analog_en[3]
port 462 nsew
flabel metal3 s 633270 200347 633750 200417 0 FreeSans 400 0 0 0 gpio_analog_pol[3]
port 550 nsew
flabel metal3 s 633270 203383 633750 203453 0 FreeSans 400 0 0 0 gpio_analog_sel[3]
port 506 nsew
flabel metal3 s 633270 197863 633750 197933 0 FreeSans 400 0 0 0 gpio_dm1[3]
port 638 nsew
flabel metal3 s 633270 204027 633750 204097 0 FreeSans 400 0 0 0 gpio_dm2[3]
port 682 nsew
flabel metal3 s 633270 199703 633750 199773 0 FreeSans 400 0 0 0 gpio_dm0[3]
port 594 nsew
flabel metal3 s 633270 204671 633750 204741 0 FreeSans 400 0 0 0 gpio_holdover[3]
port 418 nsew
flabel metal3 s 633270 207707 633750 207777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[3]
port 286 nsew
flabel metal3 s 633270 200899 633750 200969 0 FreeSans 400 0 0 0 gpio_inp_dis[3]
port 242 nsew
flabel metal3 s 633270 208351 633750 208421 0 FreeSans 400 0 0 0 gpio_oeb[3]
port 198 nsew
flabel metal3 s 633270 205223 633750 205293 0 FreeSans 400 0 0 0 gpio_out[3]
port 154 nsew
flabel metal3 s 633270 196023 633750 196093 0 FreeSans 400 0 0 0 gpio_slow_sel[3]
port 374 nsew
flabel metal3 s 633270 207063 633750 207133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[3]
port 330 nsew
flabel metal3 s 633270 63659 633750 63729 0 FreeSans 400 0 0 0 gpio_analog_en[0]
port 465 nsew
flabel metal3 s 633270 64947 633750 65017 0 FreeSans 400 0 0 0 gpio_analog_pol[0]
port 553 nsew
flabel metal3 s 633270 67983 633750 68053 0 FreeSans 400 0 0 0 gpio_analog_sel[0]
port 509 nsew
flabel metal3 s 633270 64303 633750 64373 0 FreeSans 400 0 0 0 gpio_dm0[0]
port 597 nsew
flabel metal3 s 633270 62463 633750 62533 0 FreeSans 400 0 0 0 gpio_dm1[0]
port 641 nsew
flabel metal3 s 633270 68627 633750 68697 0 FreeSans 400 0 0 0 gpio_dm2[0]
port 685 nsew
flabel metal3 s 633270 69271 633750 69341 0 FreeSans 400 0 0 0 gpio_holdover[0]
port 421 nsew
flabel metal3 s 633270 72307 633750 72377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[0]
port 289 nsew
flabel metal3 s 633270 65499 633750 65569 0 FreeSans 400 0 0 0 gpio_inp_dis[0]
port 245 nsew
flabel metal3 s 633270 72951 633750 73021 0 FreeSans 400 0 0 0 gpio_oeb[0]
port 201 nsew
flabel metal3 s 633270 69823 633750 69893 0 FreeSans 400 0 0 0 gpio_out[0]
port 157 nsew
flabel metal3 s 633270 60623 633750 60693 0 FreeSans 400 0 0 0 gpio_slow_sel[0]
port 377 nsew
flabel metal3 s 633270 71663 633750 71733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[0]
port 333 nsew
flabel metal3 s 633270 58783 633750 58853 0 FreeSans 400 0 0 0 gpio_in[0]
port 729 nsew
flabel metal3 s 633270 194183 633750 194253 0 FreeSans 400 0 0 0 gpio_in[3]
port 726 nsew
flabel metal3 633270 61267 633750 61337 0 FreeSans 400 0 0 0 analog_io[0]
port 905 nsew
flabel metal3 633270 63107 633750 63177 0 FreeSans 400 0 0 0 analog_noesd_io[0]
port 949 nsew
flabel metal3 633270 108307 633750 108377 0 FreeSans 400 0 0 0 analog_noesd_io[1]
port 948 nsew
flabel metal3 633270 106467 633750 106537 0 FreeSans 400 0 0 0 analog_io[1]
port 904 nsew
flabel metal3 633270 73503 633750 73573 0 FreeSans 400 0 0 0 gpio_in_h[0]
port 773 nsew
flabel metal3 633270 118703 633750 118773 0 FreeSans 400 0 0 0 gpio_in_h[1]
port 772 nsew
flabel metal3 633270 151467 633750 151537 0 FreeSans 400 0 0 0 analog_io[2]
port 903 nsew
flabel metal3 633270 153307 633750 153377 0 FreeSans 400 0 0 0 analog_noesd_io[2]
port 947 nsew
flabel metal3 633270 163703 633750 163773 0 FreeSans 400 0 0 0 gpio_in_h[2]
port 771 nsew
flabel metal3 633270 196667 633750 196737 0 FreeSans 400 0 0 0 analog_io[3]
port 902 nsew
flabel metal3 633270 198507 633750 198577 0 FreeSans 400 0 0 0 analog_noesd_io[3]
port 946 nsew
flabel metal3 633270 208903 633750 208973 0 FreeSans 400 0 0 0 gpio_in_h[3]
port 770 nsew
flabel metal3 633270 241667 633750 241737 0 FreeSans 400 0 0 0 analog_io[4]
port 901 nsew
flabel metal3 633270 243507 633750 243577 0 FreeSans 400 0 0 0 analog_noesd_io[4]
port 945 nsew
flabel metal3 633270 253903 633750 253973 0 FreeSans 400 0 0 0 gpio_in_h[4]
port 769 nsew
flabel metal3 633270 286667 633750 286737 0 FreeSans 400 0 0 0 analog_io[5]
port 900 nsew
flabel metal3 633270 288507 633750 288577 0 FreeSans 400 0 0 0 analog_noesd_io[5]
port 944 nsew
flabel metal3 633270 298903 633750 298973 0 FreeSans 400 0 0 0 gpio_in_h[5]
port 768 nsew
flabel metal3 633270 331867 633750 331937 0 FreeSans 400 0 0 0 analog_io[6]
port 899 nsew
flabel metal3 633270 333707 633750 333777 0 FreeSans 400 0 0 0 analog_noesd_io[6]
port 943 nsew
flabel metal3 633270 344103 633750 344173 0 FreeSans 400 0 0 0 gpio_in_h[6]
port 767 nsew
flabel metal3 s 633270 509067 633750 509137 0 FreeSans 400 0 0 0 analog_io[7]
port 898 nsew
flabel metal3 s 633270 510907 633750 510977 0 FreeSans 400 0 0 0 analog_noesd_io[7]
port 942 nsew
flabel metal3 s 633270 521303 633750 521373 0 FreeSans 400 0 0 0 gpio_in_h[7]
port 766 nsew
flabel metal3 s 633270 554267 633750 554337 0 FreeSans 400 0 0 0 analog_io[8]
port 897 nsew
flabel metal3 s 633270 556107 633750 556177 0 FreeSans 400 0 0 0 analog_noesd_io[8]
port 941 nsew
flabel metal3 s 633270 566503 633750 566573 0 FreeSans 400 0 0 0 gpio_in_h[8]
port 765 nsew
flabel metal3 s 633270 599267 633750 599337 0 FreeSans 400 0 0 0 analog_io[9]
port 896 nsew
flabel metal3 s 633270 601107 633750 601177 0 FreeSans 400 0 0 0 analog_noesd_io[9]
port 940 nsew
flabel metal3 s 633270 611503 633750 611573 0 FreeSans 400 0 0 0 gpio_in_h[9]
port 764 nsew
flabel metal3 s 633270 644467 633750 644537 0 FreeSans 400 0 0 0 analog_io[10]
port 895 nsew
flabel metal3 s 633270 646307 633750 646377 0 FreeSans 400 0 0 0 analog_noesd_io[10]
port 939 nsew
flabel metal3 s 633270 656703 633750 656773 0 FreeSans 400 0 0 0 gpio_in_h[10]
port 763 nsew
flabel metal3 s 633270 689467 633750 689537 0 FreeSans 400 0 0 0 analog_io[11]
port 894 nsew
flabel metal3 s 633270 691307 633750 691377 0 FreeSans 400 0 0 0 analog_noesd_io[11]
port 938 nsew
flabel metal3 s 633270 701703 633750 701773 0 FreeSans 400 0 0 0 gpio_in_h[11]
port 762 nsew
flabel metal3 s 633270 746703 633750 746773 0 FreeSans 400 0 0 0 gpio_in_h[12]
port 761 nsew
flabel metal3 s 633270 835903 633750 835973 0 FreeSans 400 0 0 0 gpio_in_h[13]
port 760 nsew
flabel metal3 s 633270 925103 633750 925173 0 FreeSans 400 0 0 0 gpio_in_h[14]
port 759 nsew
flabel metal3 s 633270 734467 633750 734537 0 FreeSans 400 0 0 0 analog_io[12]
port 893 nsew
flabel metal3 s 633270 823667 633750 823737 0 FreeSans 400 0 0 0 analog_io[13]
port 892 nsew
flabel metal3 s 633270 912867 633750 912937 0 FreeSans 400 0 0 0 analog_io[14]
port 891 nsew
flabel metal3 s 633270 736307 633750 736377 0 FreeSans 400 0 0 0 analog_noesd_io[12]
port 937 nsew
flabel metal3 s 633270 825507 633750 825577 0 FreeSans 400 0 0 0 analog_noesd_io[13]
port 936 nsew
flabel metal3 s 633270 914707 633750 914777 0 FreeSans 400 0 0 0 analog_noesd_io[14]
port 935 nsew
flabel metal3 s -424 922197 56 922267 0 FreeSans 400 0 0 0 gpio_analog_en[24]
port 441 nsew
flabel metal3 s -424 920909 56 920979 0 FreeSans 400 0 0 0 gpio_analog_pol[24]
port 529 nsew
flabel metal3 s -424 917873 56 917943 0 FreeSans 400 0 0 0 gpio_analog_sel[24]
port 485 nsew
flabel metal3 s -424 921553 56 921623 0 FreeSans 400 0 0 0 gpio_dm0[24]
port 573 nsew
flabel metal3 s -424 923393 56 923463 0 FreeSans 400 0 0 0 gpio_dm1[24]
port 617 nsew
flabel metal3 s -424 917229 56 917299 0 FreeSans 400 0 0 0 gpio_dm2[24]
port 661 nsew
flabel metal3 s -424 916585 56 916655 0 FreeSans 400 0 0 0 gpio_holdover[24]
port 397 nsew
flabel metal3 s -424 913549 56 913619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[24]
port 265 nsew
flabel metal3 s -424 920357 56 920427 0 FreeSans 400 0 0 0 gpio_inp_dis[24]
port 221 nsew
flabel metal3 s -424 912905 56 912975 0 FreeSans 400 0 0 0 gpio_oeb[24]
port 177 nsew
flabel metal3 s -424 916033 56 916103 0 FreeSans 400 0 0 0 gpio_out[24]
port 133 nsew
flabel metal3 s -424 925233 56 925303 0 FreeSans 400 0 0 0 gpio_slow_sel[24]
port 353 nsew
flabel metal3 s -424 914193 56 914263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[24]
port 309 nsew
flabel metal3 s -424 927073 56 927143 0 FreeSans 400 0 0 0 gpio_in[24]
port 705 nsew
flabel metal3 s -424 912353 56 912423 0 FreeSans 400 0 0 0 gpio_in_h[24]
port 749 nsew
flabel metal3 s -424 924589 56 924659 0 FreeSans 400 0 0 0 analog_io[24]
port 881 nsew
flabel metal3 s -424 922749 56 922819 0 FreeSans 400 0 0 0 analog_noesd_io[24]
port 925 nsew
flabel metal3 s -424 752397 56 752467 0 FreeSans 400 0 0 0 gpio_analog_en[25]
port 440 nsew
flabel metal3 s -424 751109 56 751179 0 FreeSans 400 0 0 0 gpio_analog_pol[25]
port 528 nsew
flabel metal3 s -424 748073 56 748143 0 FreeSans 400 0 0 0 gpio_analog_sel[25]
port 484 nsew
flabel metal3 s -424 751753 56 751823 0 FreeSans 400 0 0 0 gpio_dm0[25]
port 572 nsew
flabel metal3 s -424 753593 56 753663 0 FreeSans 400 0 0 0 gpio_dm1[25]
port 616 nsew
flabel metal3 s -424 747429 56 747499 0 FreeSans 400 0 0 0 gpio_dm2[25]
port 660 nsew
flabel metal3 s -424 746785 56 746855 0 FreeSans 400 0 0 0 gpio_holdover[25]
port 396 nsew
flabel metal3 s -424 743749 56 743819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[25]
port 264 nsew
flabel metal3 s -424 750557 56 750627 0 FreeSans 400 0 0 0 gpio_inp_dis[25]
port 220 nsew
flabel metal3 s -424 743105 56 743175 0 FreeSans 400 0 0 0 gpio_oeb[25]
port 176 nsew
flabel metal3 s -424 746233 56 746303 0 FreeSans 400 0 0 0 gpio_out[25]
port 132 nsew
flabel metal3 s -424 755433 56 755503 0 FreeSans 400 0 0 0 gpio_slow_sel[25]
port 352 nsew
flabel metal3 s -424 757273 56 757343 0 FreeSans 400 0 0 0 gpio_in[25]
port 704 nsew
flabel metal3 s -424 535753 56 535823 0 FreeSans 400 0 0 0 gpio_dm0[30]
port 567 nsew
flabel metal3 s -424 537593 56 537663 0 FreeSans 400 0 0 0 gpio_dm1[30]
port 611 nsew
flabel metal3 s -424 531429 56 531499 0 FreeSans 400 0 0 0 gpio_dm2[30]
port 655 nsew
flabel metal3 s -424 530785 56 530855 0 FreeSans 400 0 0 0 gpio_holdover[30]
port 391 nsew
flabel metal3 s -424 527749 56 527819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[30]
port 259 nsew
flabel metal3 s -424 534557 56 534627 0 FreeSans 400 0 0 0 gpio_inp_dis[30]
port 215 nsew
flabel metal3 s -424 527105 56 527175 0 FreeSans 400 0 0 0 gpio_oeb[30]
port 171 nsew
flabel metal3 s -424 530233 56 530303 0 FreeSans 400 0 0 0 gpio_out[30]
port 127 nsew
flabel metal3 s -424 539433 56 539503 0 FreeSans 400 0 0 0 gpio_slow_sel[30]
port 347 nsew
flabel metal3 s -424 528393 56 528463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[30]
port 303 nsew
flabel metal3 s -424 541273 56 541343 0 FreeSans 400 0 0 0 gpio_in[30]
port 699 nsew
flabel metal3 s -424 493197 56 493267 0 FreeSans 400 0 0 0 gpio_analog_en[31]
port 434 nsew
flabel metal3 s -424 491909 56 491979 0 FreeSans 400 0 0 0 gpio_analog_pol[31]
port 522 nsew
flabel metal3 s -424 488873 56 488943 0 FreeSans 400 0 0 0 gpio_analog_sel[31]
port 478 nsew
flabel metal3 s -424 492553 56 492623 0 FreeSans 400 0 0 0 gpio_dm0[31]
port 566 nsew
flabel metal3 s -424 494393 56 494463 0 FreeSans 400 0 0 0 gpio_dm1[31]
port 610 nsew
flabel metal3 s -424 488229 56 488299 0 FreeSans 400 0 0 0 gpio_dm2[31]
port 654 nsew
flabel metal3 s -424 487585 56 487655 0 FreeSans 400 0 0 0 gpio_holdover[31]
port 390 nsew
flabel metal3 s -424 484549 56 484619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[31]
port 258 nsew
flabel metal3 s -424 491357 56 491427 0 FreeSans 400 0 0 0 gpio_inp_dis[31]
port 214 nsew
flabel metal3 s -424 483905 56 483975 0 FreeSans 400 0 0 0 gpio_oeb[31]
port 170 nsew
flabel metal3 s -424 487033 56 487103 0 FreeSans 400 0 0 0 gpio_out[31]
port 126 nsew
flabel metal3 s -424 496233 56 496303 0 FreeSans 400 0 0 0 gpio_slow_sel[31]
port 346 nsew
flabel metal3 s -424 485193 56 485263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[31]
port 302 nsew
flabel metal3 s -424 498073 56 498143 0 FreeSans 400 0 0 0 gpio_in[31]
port 698 nsew
flabel metal3 s -424 709197 56 709267 0 FreeSans 400 0 0 0 gpio_analog_en[26]
port 439 nsew
flabel metal3 s -424 707909 56 707979 0 FreeSans 400 0 0 0 gpio_analog_pol[26]
port 527 nsew
flabel metal3 s -424 704873 56 704943 0 FreeSans 400 0 0 0 gpio_analog_sel[26]
port 483 nsew
flabel metal3 s -424 708553 56 708623 0 FreeSans 400 0 0 0 gpio_dm0[26]
port 571 nsew
flabel metal3 s -424 710393 56 710463 0 FreeSans 400 0 0 0 gpio_dm1[26]
port 615 nsew
flabel metal3 s -424 704229 56 704299 0 FreeSans 400 0 0 0 gpio_dm2[26]
port 659 nsew
flabel metal3 s -424 703585 56 703655 0 FreeSans 400 0 0 0 gpio_holdover[26]
port 395 nsew
flabel metal3 s -424 700549 56 700619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[26]
port 263 nsew
flabel metal3 s -424 707357 56 707427 0 FreeSans 400 0 0 0 gpio_inp_dis[26]
port 219 nsew
flabel metal3 s -424 699905 56 699975 0 FreeSans 400 0 0 0 gpio_oeb[26]
port 175 nsew
flabel metal3 s -424 703033 56 703103 0 FreeSans 400 0 0 0 gpio_out[26]
port 131 nsew
flabel metal3 s -424 712233 56 712303 0 FreeSans 400 0 0 0 gpio_slow_sel[26]
port 351 nsew
flabel metal3 s -424 701193 56 701263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[26]
port 307 nsew
flabel metal3 s -424 714073 56 714143 0 FreeSans 400 0 0 0 gpio_in[26]
port 703 nsew
flabel metal3 s -424 665997 56 666067 0 FreeSans 400 0 0 0 gpio_analog_en[27]
port 438 nsew
flabel metal3 s -424 664709 56 664779 0 FreeSans 400 0 0 0 gpio_analog_pol[27]
port 526 nsew
flabel metal3 s -424 661673 56 661743 0 FreeSans 400 0 0 0 gpio_analog_sel[27]
port 482 nsew
flabel metal3 s -424 665353 56 665423 0 FreeSans 400 0 0 0 gpio_dm0[27]
port 570 nsew
flabel metal3 s -424 667193 56 667263 0 FreeSans 400 0 0 0 gpio_dm1[27]
port 614 nsew
flabel metal3 s -424 661029 56 661099 0 FreeSans 400 0 0 0 gpio_dm2[27]
port 658 nsew
flabel metal3 s -424 660385 56 660455 0 FreeSans 400 0 0 0 gpio_holdover[27]
port 394 nsew
flabel metal3 s -424 657349 56 657419 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[27]
port 262 nsew
flabel metal3 s -424 664157 56 664227 0 FreeSans 400 0 0 0 gpio_inp_dis[27]
port 218 nsew
flabel metal3 s -424 656705 56 656775 0 FreeSans 400 0 0 0 gpio_oeb[27]
port 174 nsew
flabel metal3 s -424 659833 56 659903 0 FreeSans 400 0 0 0 gpio_out[27]
port 130 nsew
flabel metal3 s -424 669033 56 669103 0 FreeSans 400 0 0 0 gpio_slow_sel[27]
port 350 nsew
flabel metal3 s -424 657993 56 658063 0 FreeSans 400 0 0 0 gpio_vtrip_sel[27]
port 306 nsew
flabel metal3 s -424 670873 56 670943 0 FreeSans 400 0 0 0 gpio_in[27]
port 702 nsew
flabel metal3 s -424 622797 56 622867 0 FreeSans 400 0 0 0 gpio_analog_en[28]
port 437 nsew
flabel metal3 s -424 621509 56 621579 0 FreeSans 400 0 0 0 gpio_analog_pol[28]
port 525 nsew
flabel metal3 s -424 618473 56 618543 0 FreeSans 400 0 0 0 gpio_analog_sel[28]
port 481 nsew
flabel metal3 s -424 622153 56 622223 0 FreeSans 400 0 0 0 gpio_dm0[28]
port 569 nsew
flabel metal3 s -424 623993 56 624063 0 FreeSans 400 0 0 0 gpio_dm1[28]
port 613 nsew
flabel metal3 s -424 617829 56 617899 0 FreeSans 400 0 0 0 gpio_dm2[28]
port 657 nsew
flabel metal3 s -424 617185 56 617255 0 FreeSans 400 0 0 0 gpio_holdover[28]
port 393 nsew
flabel metal3 s -424 614149 56 614219 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[28]
port 261 nsew
flabel metal3 s -424 620957 56 621027 0 FreeSans 400 0 0 0 gpio_inp_dis[28]
port 217 nsew
flabel metal3 s -424 613505 56 613575 0 FreeSans 400 0 0 0 gpio_oeb[28]
port 173 nsew
flabel metal3 s -424 616633 56 616703 0 FreeSans 400 0 0 0 gpio_out[28]
port 129 nsew
flabel metal3 s -424 625833 56 625903 0 FreeSans 400 0 0 0 gpio_slow_sel[28]
port 349 nsew
flabel metal3 s -424 614793 56 614863 0 FreeSans 400 0 0 0 gpio_vtrip_sel[28]
port 305 nsew
flabel metal3 s -424 627673 56 627743 0 FreeSans 400 0 0 0 gpio_in[28]
port 701 nsew
flabel metal3 s -424 579597 56 579667 0 FreeSans 400 0 0 0 gpio_analog_en[29]
port 436 nsew
flabel metal3 s -424 578309 56 578379 0 FreeSans 400 0 0 0 gpio_analog_pol[29]
port 524 nsew
flabel metal3 s -424 575273 56 575343 0 FreeSans 400 0 0 0 gpio_analog_sel[29]
port 480 nsew
flabel metal3 s -424 578953 56 579023 0 FreeSans 400 0 0 0 gpio_dm0[29]
port 568 nsew
flabel metal3 s -424 580793 56 580863 0 FreeSans 400 0 0 0 gpio_dm1[29]
port 612 nsew
flabel metal3 s -424 574629 56 574699 0 FreeSans 400 0 0 0 gpio_dm2[29]
port 656 nsew
flabel metal3 s -424 573985 56 574055 0 FreeSans 400 0 0 0 gpio_holdover[29]
port 392 nsew
flabel metal3 s -424 570949 56 571019 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[29]
port 260 nsew
flabel metal3 s -424 577757 56 577827 0 FreeSans 400 0 0 0 gpio_inp_dis[29]
port 216 nsew
flabel metal3 s -424 570305 56 570375 0 FreeSans 400 0 0 0 gpio_oeb[29]
port 172 nsew
flabel metal3 s -424 573433 56 573503 0 FreeSans 400 0 0 0 gpio_out[29]
port 128 nsew
flabel metal3 s -424 582633 56 582703 0 FreeSans 400 0 0 0 gpio_slow_sel[29]
port 348 nsew
flabel metal3 s -424 571593 56 571663 0 FreeSans 400 0 0 0 gpio_vtrip_sel[29]
port 304 nsew
flabel metal3 s -424 584473 56 584543 0 FreeSans 400 0 0 0 gpio_in[29]
port 700 nsew
flabel metal3 s -424 536397 56 536467 0 FreeSans 400 0 0 0 gpio_analog_en[30]
port 435 nsew
flabel metal3 s -424 535109 56 535179 0 FreeSans 400 0 0 0 gpio_analog_pol[30]
port 523 nsew
flabel metal3 s -424 532073 56 532143 0 FreeSans 400 0 0 0 gpio_analog_sel[30]
port 479 nsew
flabel metal3 s -424 193993 56 194064 0 FreeSans 400 0 0 0 gpio_dm1[36]
port 605 nsew
flabel metal3 s -424 187829 56 187900 0 FreeSans 400 0 0 0 gpio_dm2[36]
port 649 nsew
flabel metal3 s -424 187185 56 187256 0 FreeSans 400 0 0 0 gpio_holdover[36]
port 385 nsew
flabel metal3 s -424 184149 56 184220 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[36]
port 253 nsew
flabel metal3 s -424 190957 56 191028 0 FreeSans 400 0 0 0 gpio_inp_dis[36]
port 209 nsew
flabel metal3 s -424 183505 56 183576 0 FreeSans 400 0 0 0 gpio_oeb[36]
port 165 nsew
flabel metal3 s -424 186633 56 186704 0 FreeSans 400 0 0 0 gpio_out[36]
port 121 nsew
flabel metal3 s -424 195833 56 195904 0 FreeSans 400 0 0 0 gpio_slow_sel[36]
port 341 nsew
flabel metal3 s -424 184793 56 184864 0 FreeSans 400 0 0 0 gpio_vtrip_sel[36]
port 297 nsew
flabel metal3 s -424 197673 56 197744 0 FreeSans 400 0 0 0 gpio_in[36]
port 693 nsew
flabel metal3 s -424 149597 56 149668 0 FreeSans 400 0 0 0 gpio_analog_en[37]
port 428 nsew
flabel metal3 s -424 148309 56 148380 0 FreeSans 400 0 0 0 gpio_analog_pol[37]
port 516 nsew
flabel metal3 s -424 145273 56 145344 0 FreeSans 400 0 0 0 gpio_analog_sel[37]
port 472 nsew
flabel metal3 s -424 148953 56 149024 0 FreeSans 400 0 0 0 gpio_dm0[37]
port 560 nsew
flabel metal3 s -424 150793 56 150864 0 FreeSans 400 0 0 0 gpio_dm1[37]
port 604 nsew
flabel metal3 s -424 144629 56 144700 0 FreeSans 400 0 0 0 gpio_dm2[37]
port 648 nsew
flabel metal3 s -424 143985 56 144056 0 FreeSans 400 0 0 0 gpio_holdover[37]
port 384 nsew
flabel metal3 s -424 140949 56 141020 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[37]
port 252 nsew
flabel metal3 s -424 140305 56 140376 0 FreeSans 400 0 0 0 gpio_oeb[37]
port 164 nsew
flabel metal3 s -424 143433 56 143504 0 FreeSans 400 0 0 0 gpio_out[37]
port 120 nsew
flabel metal3 s -424 152633 56 152704 0 FreeSans 400 0 0 0 gpio_slow_sel[37]
port 340 nsew
flabel metal3 s -424 154473 56 154544 0 FreeSans 400 0 0 0 gpio_in[37]
port 692 nsew
flabel metal3 s -424 365597 56 365667 0 FreeSans 400 0 0 0 gpio_analog_en[32]
port 433 nsew
flabel metal3 s -424 364309 56 364379 0 FreeSans 400 0 0 0 gpio_analog_pol[32]
port 521 nsew
flabel metal3 s -424 361273 56 361343 0 FreeSans 400 0 0 0 gpio_analog_sel[32]
port 477 nsew
flabel metal3 s -424 364953 56 365023 0 FreeSans 400 0 0 0 gpio_dm0[32]
port 565 nsew
flabel metal3 s -424 366793 56 366863 0 FreeSans 400 0 0 0 gpio_dm1[32]
port 609 nsew
flabel metal3 s -424 360629 56 360699 0 FreeSans 400 0 0 0 gpio_dm2[32]
port 653 nsew
flabel metal3 s -424 359985 56 360055 0 FreeSans 400 0 0 0 gpio_holdover[32]
port 389 nsew
flabel metal3 s -424 356949 56 357019 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[32]
port 257 nsew
flabel metal3 s -424 363757 56 363827 0 FreeSans 400 0 0 0 gpio_inp_dis[32]
port 213 nsew
flabel metal3 s -424 356305 56 356375 0 FreeSans 400 0 0 0 gpio_oeb[32]
port 169 nsew
flabel metal3 s -424 359433 56 359503 0 FreeSans 400 0 0 0 gpio_out[32]
port 125 nsew
flabel metal3 s -424 368633 56 368703 0 FreeSans 400 0 0 0 gpio_slow_sel[32]
port 345 nsew
flabel metal3 s -424 357593 56 357663 0 FreeSans 400 0 0 0 gpio_vtrip_sel[32]
port 301 nsew
flabel metal3 s -424 370473 56 370543 0 FreeSans 400 0 0 0 gpio_in[32]
port 697 nsew
flabel metal3 s -424 322397 56 322467 0 FreeSans 400 0 0 0 gpio_analog_en[33]
port 432 nsew
flabel metal3 s -424 318073 56 318143 0 FreeSans 400 0 0 0 gpio_analog_sel[33]
port 476 nsew
flabel metal3 s -424 323593 56 323663 0 FreeSans 400 0 0 0 gpio_dm1[33]
port 608 nsew
flabel metal3 s -424 317429 56 317499 0 FreeSans 400 0 0 0 gpio_dm2[33]
port 652 nsew
flabel metal3 s -424 321753 56 321823 0 FreeSans 400 0 0 0 gpio_dm0[33]
port 564 nsew
flabel metal3 s -424 316785 56 316855 0 FreeSans 400 0 0 0 gpio_holdover[33]
port 388 nsew
flabel metal3 s -424 313749 56 313819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[33]
port 256 nsew
flabel metal3 s -424 320557 56 320627 0 FreeSans 400 0 0 0 gpio_inp_dis[33]
port 212 nsew
flabel metal3 s -424 313105 56 313175 0 FreeSans 400 0 0 0 gpio_oeb[33]
port 168 nsew
flabel metal3 s -424 316233 56 316303 0 FreeSans 400 0 0 0 gpio_out[33]
port 124 nsew
flabel metal3 s -424 325433 56 325503 0 FreeSans 400 0 0 0 gpio_slow_sel[33]
port 344 nsew
flabel metal3 s -424 314393 56 314463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[33]
port 300 nsew
flabel metal3 s -424 327273 56 327343 0 FreeSans 400 0 0 0 gpio_in[33]
port 696 nsew
flabel metal3 s -424 279197 56 279267 0 FreeSans 400 0 0 0 gpio_analog_en[34]
port 431 nsew
flabel metal3 s -424 277909 56 277979 0 FreeSans 400 0 0 0 gpio_analog_pol[34]
port 519 nsew
flabel metal3 s -424 274873 56 274943 0 FreeSans 400 0 0 0 gpio_analog_sel[34]
port 475 nsew
flabel metal3 s -424 278553 56 278623 0 FreeSans 400 0 0 0 gpio_dm0[34]
port 563 nsew
flabel metal3 s -424 280393 56 280463 0 FreeSans 400 0 0 0 gpio_dm1[34]
port 607 nsew
flabel metal3 s -424 274229 56 274299 0 FreeSans 400 0 0 0 gpio_dm2[34]
port 651 nsew
flabel metal3 s -424 273585 56 273655 0 FreeSans 400 0 0 0 gpio_holdover[34]
port 387 nsew
flabel metal3 s -424 270549 56 270619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[34]
port 255 nsew
flabel metal3 s -424 277357 56 277427 0 FreeSans 400 0 0 0 gpio_inp_dis[34]
port 211 nsew
flabel metal3 s -424 269905 56 269975 0 FreeSans 400 0 0 0 gpio_oeb[34]
port 167 nsew
flabel metal3 s -424 273033 56 273103 0 FreeSans 400 0 0 0 gpio_out[34]
port 123 nsew
flabel metal3 s -424 282233 56 282303 0 FreeSans 400 0 0 0 gpio_slow_sel[34]
port 343 nsew
flabel metal3 s -424 271193 56 271263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[34]
port 299 nsew
flabel metal3 s -424 284073 56 284143 0 FreeSans 400 0 0 0 gpio_in[34]
port 695 nsew
flabel metal3 s -424 235997 56 236067 0 FreeSans 400 0 0 0 gpio_analog_en[35]
port 430 nsew
flabel metal3 s -424 234709 56 234779 0 FreeSans 400 0 0 0 gpio_analog_pol[35]
port 518 nsew
flabel metal3 s -424 231673 56 231743 0 FreeSans 400 0 0 0 gpio_analog_sel[35]
port 474 nsew
flabel metal3 s -424 235353 56 235423 0 FreeSans 400 0 0 0 gpio_dm0[35]
port 562 nsew
flabel metal3 s -424 237193 56 237263 0 FreeSans 400 0 0 0 gpio_dm1[35]
port 606 nsew
flabel metal3 s -424 231029 56 231099 0 FreeSans 400 0 0 0 gpio_dm2[35]
port 650 nsew
flabel metal3 s -424 230385 56 230455 0 FreeSans 400 0 0 0 gpio_holdover[35]
port 386 nsew
flabel metal3 s -424 227349 56 227419 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[35]
port 254 nsew
flabel metal3 s -424 234157 56 234227 0 FreeSans 400 0 0 0 gpio_inp_dis[35]
port 210 nsew
flabel metal3 s -424 226705 56 226775 0 FreeSans 400 0 0 0 gpio_oeb[35]
port 166 nsew
flabel metal3 s -424 229833 56 229903 0 FreeSans 400 0 0 0 gpio_out[35]
port 122 nsew
flabel metal3 s -424 239033 56 239103 0 FreeSans 400 0 0 0 gpio_slow_sel[35]
port 342 nsew
flabel metal3 s -424 227993 56 228063 0 FreeSans 400 0 0 0 gpio_vtrip_sel[35]
port 298 nsew
flabel metal3 s -424 240873 56 240943 0 FreeSans 400 0 0 0 gpio_in[35]
port 694 nsew
flabel metal3 s -424 192797 56 192868 0 FreeSans 400 0 0 0 gpio_analog_en[36]
port 429 nsew
flabel metal3 s -424 191509 56 191580 0 FreeSans 400 0 0 0 gpio_analog_pol[36]
port 517 nsew
flabel metal3 s -424 188473 56 188544 0 FreeSans 400 0 0 0 gpio_analog_sel[36]
port 473 nsew
flabel metal3 s -424 192153 56 192224 0 FreeSans 400 0 0 0 gpio_dm0[36]
port 561 nsew
flabel metal3 s -424 147757 56 147828 0 FreeSans 400 0 0 0 gpio_inp_dis[37]
port 208 nsew
flabel metal3 s -424 742553 56 742623 0 FreeSans 400 0 0 0 gpio_in_h[25]
port 748 nsew
flabel metal3 s -424 699353 56 699423 0 FreeSans 400 0 0 0 gpio_in_h[26]
port 747 nsew
flabel metal3 s -424 656153 56 656223 0 FreeSans 400 0 0 0 gpio_in_h[27]
port 746 nsew
flabel metal3 s -424 612953 56 613023 0 FreeSans 400 0 0 0 gpio_in_h[28]
port 745 nsew
flabel metal3 s -424 569753 56 569823 0 FreeSans 400 0 0 0 gpio_in_h[29]
port 744 nsew
flabel metal3 s -424 526553 56 526623 0 FreeSans 400 0 0 0 gpio_in_h[30]
port 743 nsew
flabel metal3 s -424 483353 56 483423 0 FreeSans 400 0 0 0 gpio_in_h[31]
port 742 nsew
flabel metal3 s -424 355753 56 355823 0 FreeSans 400 0 0 0 gpio_in_h[32]
port 741 nsew
flabel metal3 s -424 312553 56 312623 0 FreeSans 400 0 0 0 gpio_in_h[33]
port 740 nsew
flabel metal3 s -424 269353 56 269423 0 FreeSans 400 0 0 0 gpio_in_h[34]
port 739 nsew
flabel metal3 s -424 226153 56 226223 0 FreeSans 400 0 0 0 gpio_in_h[35]
port 738 nsew
flabel metal3 s -424 182953 56 183024 0 FreeSans 400 0 0 0 gpio_in_h[36]
port 737 nsew
flabel metal3 s -424 139753 56 139824 0 FreeSans 400 0 0 0 gpio_in_h[37]
port 736 nsew
flabel metal3 s -424 754789 56 754859 0 FreeSans 400 0 0 0 analog_io[25]
port 880 nsew
flabel metal3 s -424 711589 56 711659 0 FreeSans 400 0 0 0 analog_io[26]
port 879 nsew
flabel metal3 s -424 668389 56 668459 0 FreeSans 400 0 0 0 analog_io[27]
port 878 nsew
flabel metal3 s -424 625189 56 625259 0 FreeSans 400 0 0 0 analog_io[28]
port 877 nsew
flabel metal3 s -424 581989 56 582059 0 FreeSans 400 0 0 0 analog_io[29]
port 876 nsew
flabel metal3 s -424 538789 56 538859 0 FreeSans 400 0 0 0 analog_io[30]
port 875 nsew
flabel metal3 s -424 495589 56 495659 0 FreeSans 400 0 0 0 analog_io[31]
port 874 nsew
flabel metal3 s -424 367989 56 368059 0 FreeSans 400 0 0 0 analog_io[32]
port 873 nsew
flabel metal3 s -424 324789 56 324859 0 FreeSans 400 0 0 0 analog_io[33]
port 872 nsew
flabel metal3 s -424 281589 56 281659 0 FreeSans 400 0 0 0 analog_io[34]
port 871 nsew
flabel metal3 s -424 238389 56 238459 0 FreeSans 400 0 0 0 analog_io[35]
port 870 nsew
flabel metal3 s -424 195189 56 195260 0 FreeSans 400 0 0 0 analog_io[36]
port 869 nsew
flabel metal3 s -424 151989 56 152060 0 FreeSans 400 0 0 0 analog_io[37]
port 868 nsew
flabel metal3 s -424 752949 56 753019 0 FreeSans 400 0 0 0 analog_noesd_io[25]
port 924 nsew
flabel metal3 s -424 709749 56 709819 0 FreeSans 400 0 0 0 analog_noesd_io[26]
port 923 nsew
flabel metal3 s -424 666549 56 666619 0 FreeSans 400 0 0 0 analog_noesd_io[27]
port 922 nsew
flabel metal3 s -424 623349 56 623419 0 FreeSans 400 0 0 0 analog_noesd_io[28]
port 921 nsew
flabel metal3 s -424 580149 56 580219 0 FreeSans 400 0 0 0 analog_noesd_io[29]
port 920 nsew
flabel metal3 s -424 536949 56 537019 0 FreeSans 400 0 0 0 analog_noesd_io[30]
port 919 nsew
flabel metal3 s -424 493749 56 493819 0 FreeSans 400 0 0 0 analog_noesd_io[31]
port 918 nsew
flabel metal3 s -424 366149 56 366219 0 FreeSans 400 0 0 0 analog_noesd_io[32]
port 917 nsew
flabel metal3 s -424 322949 56 323019 0 FreeSans 400 0 0 0 analog_noesd_io[33]
port 916 nsew
flabel metal3 s -424 279749 56 279819 0 FreeSans 400 0 0 0 analog_noesd_io[34]
port 915 nsew
flabel metal3 s -424 236549 56 236619 0 FreeSans 400 0 0 0 analog_noesd_io[35]
port 914 nsew
flabel metal3 s -424 193349 56 193420 0 FreeSans 400 0 0 0 analog_noesd_io[36]
port 913 nsew
flabel metal3 s -424 150149 56 150220 0 FreeSans 400 0 0 0 analog_noesd_io[37]
port 912 nsew
flabel metal3 s -424 744393 56 744463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[25]
port 308 nsew
flabel metal3 s -424 321109 56 321179 0 FreeSans 400 0 0 0 gpio_analog_pol[33]
port 520 nsew
flabel metal3 -264 906644 56 906704 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal3 -264 736644 56 736704 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel metal3 -264 693644 56 693704 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 -264 650644 56 650704 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 -264 607644 56 607704 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 -264 564644 56 564704 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 -264 521644 56 521704 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 -264 478644 56 478704 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 -264 349644 56 349704 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 -264 306644 56 306704 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 -264 263644 56 263704 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 -264 220644 56 220704 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 -264 177644 56 177704 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 -264 134644 56 134704 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal2 s 488380 -260 488432 56 0 FreeSans 400 90 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 s 492635 -260 492687 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[43]
port 774 nsew
flabel metal2 s 433580 -260 433632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 s 437778 -260 437830 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[42]
port 775 nsew
flabel metal2 s 378780 -260 378832 56 0 FreeSans 400 90 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 s 382978 -260 383030 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[41]
port 776 nsew
flabel metal2 s 323980 -260 324032 56 0 FreeSans 400 90 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 s 328165 -282 328217 34 0 FreeSans 400 90 0 0 gpio_loopback_zero[40]
port 777 nsew
flabel metal2 s 269180 -260 269232 56 0 FreeSans 400 90 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 s 273360 -260 273412 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[39]
port 778 nsew
flabel metal2 s 160580 -260 160632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 s 163791 -259 163843 57 0 FreeSans 400 90 0 0 gpio_loopback_zero[38]
port 779 nsew
flabel metal2 s 110164 -116 110220 56 0 FreeSans 400 90 0 0 resetb_l
port 37 nsew
flabel metal2 s 99571 -90 99637 56 0 FreeSans 400 90 0 0 resetb_h
port 36 nsew
flabel metal3 -283 53372 56 53442 0 FreeSans 400 0 0 0 por_l
port 35 nsew
flabel metal3 -283 53595 56 53665 0 FreeSans 400 0 0 0 porb_l
port 34 nsew
flabel metal2 s 605082 -260 605134 56 0 FreeSans 400 90 0 0 mask_rev[0]
port 69 nsew
flabel metal3 -283 53147 56 53217 0 FreeSans 400 0 0 0 porb_h
port 33 nsew
flabel metal2 578298 953270 578359 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[15]
port 846 nsew
flabel metal2 478898 953270 478959 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[16]
port 845 nsew
flabel metal2 427698 953270 427759 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[17]
port 844 nsew
flabel metal2 338698 953270 338759 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[18]
port 843 nsew
flabel metal2 234298 953270 234359 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[19]
port 842 nsew
flabel metal2 183098 953270 183159 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[20]
port 841 nsew
flabel metal2 131898 953270 131959 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[21]
port 840 nsew
flabel metal2 80698 953270 80759 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[22]
port 839 nsew
flabel metal2 29498 953270 29559 953590 0 FreeSans 400 90 0 0 gpio_loopback_one[23]
port 838 nsew
flabel metal3 633270 927005 633590 927067 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 633270 837005 633590 837067 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 633270 748005 633590 748067 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 633270 703005 633590 703067 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 633270 658005 633590 658067 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 633270 613005 633590 613067 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 633270 568005 633590 568067 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 633270 523005 633590 523067 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 633270 346005 633590 346067 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 633270 301005 633590 301067 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 633270 256005 633590 256067 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 633270 211005 633590 211067 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 633270 166005 633590 166067 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 633270 121005 633590 121067 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 633270 76005 633590 76067 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal2 s 605978 -260 606030 56 0 FreeSans 400 90 0 0 mask_rev[4]
port 65 nsew
flabel metal2 s 606202 -260 606254 56 0 FreeSans 400 90 0 0 mask_rev[5]
port 64 nsew
flabel metal2 s 606426 -260 606478 56 0 FreeSans 400 90 0 0 mask_rev[6]
port 63 nsew
flabel metal2 s 606650 -260 606702 56 0 FreeSans 400 90 0 0 mask_rev[7]
port 62 nsew
flabel metal2 s 606874 -260 606926 56 0 FreeSans 400 90 0 0 mask_rev[8]
port 61 nsew
flabel metal2 s 607098 -260 607150 56 0 FreeSans 400 90 0 0 mask_rev[9]
port 60 nsew
flabel metal2 s 607322 -260 607374 56 0 FreeSans 400 90 0 0 mask_rev[10]
port 59 nsew
flabel metal2 s 607546 -260 607598 56 0 FreeSans 400 90 0 0 mask_rev[11]
port 58 nsew
flabel metal2 s 607770 -260 607822 56 0 FreeSans 400 90 0 0 mask_rev[12]
port 57 nsew
flabel metal2 s 607994 -260 608046 56 0 FreeSans 400 90 0 0 mask_rev[13]
port 56 nsew
flabel metal2 s 608218 -260 608270 56 0 FreeSans 400 90 0 0 mask_rev[14]
port 55 nsew
flabel metal2 s 608442 -260 608494 56 0 FreeSans 400 90 0 0 mask_rev[15]
port 54 nsew
flabel metal2 s 608666 -260 608718 56 0 FreeSans 400 90 0 0 mask_rev[16]
port 53 nsew
flabel metal2 s 608890 -260 608942 56 0 FreeSans 400 90 0 0 mask_rev[17]
port 52 nsew
flabel metal2 s 609114 -260 609166 56 0 FreeSans 400 90 0 0 mask_rev[18]
port 51 nsew
flabel metal2 s 609338 -260 609390 56 0 FreeSans 400 90 0 0 mask_rev[19]
port 50 nsew
flabel metal2 s 609562 -260 609614 56 0 FreeSans 400 90 0 0 mask_rev[20]
port 49 nsew
flabel metal2 s 609786 -260 609838 56 0 FreeSans 400 90 0 0 mask_rev[21]
port 48 nsew
flabel metal2 s 610010 -260 610062 56 0 FreeSans 400 90 0 0 mask_rev[22]
port 47 nsew
flabel metal2 s 610234 -260 610286 56 0 FreeSans 400 90 0 0 mask_rev[23]
port 46 nsew
flabel metal2 s 610458 -260 610510 56 0 FreeSans 400 90 0 0 mask_rev[24]
port 45 nsew
flabel metal2 s 610682 -260 610734 56 0 FreeSans 400 90 0 0 mask_rev[25]
port 44 nsew
flabel metal2 s 610906 -260 610958 56 0 FreeSans 400 90 0 0 mask_rev[26]
port 43 nsew
flabel metal2 s 611130 -260 611182 56 0 FreeSans 400 90 0 0 mask_rev[27]
port 42 nsew
flabel metal2 s 611354 -260 611406 56 0 FreeSans 400 90 0 0 mask_rev[28]
port 41 nsew
flabel metal2 s 611578 -260 611630 56 0 FreeSans 400 90 0 0 mask_rev[29]
port 40 nsew
flabel metal2 s 611802 -260 611854 56 0 FreeSans 400 90 0 0 mask_rev[30]
port 39 nsew
flabel metal2 s 612026 -260 612078 56 0 FreeSans 400 90 0 0 mask_rev[31]
port 38 nsew
flabel metal2 s 605754 -260 605806 56 0 FreeSans 400 90 0 0 mask_rev[3]
port 66 nsew
flabel metal2 s 605530 -260 605582 56 0 FreeSans 400 90 0 0 mask_rev[2]
port 67 nsew
flabel metal2 s 605306 -260 605358 56 0 FreeSans 400 90 0 0 mask_rev[1]
port 68 nsew
flabel metal3 633270 78007 633590 78069 0 FreeSans 400 0 0 0 gpio_loopback_zero[0]
port 817 nsew
flabel metal3 633270 123007 633590 123069 0 FreeSans 400 0 0 0 gpio_loopback_zero[1]
port 816 nsew
flabel metal3 633270 168007 633590 168069 0 FreeSans 400 0 0 0 gpio_loopback_zero[2]
port 815 nsew
flabel metal3 633270 213007 633590 213069 0 FreeSans 400 0 0 0 gpio_loopback_zero[3]
port 814 nsew
flabel metal3 633270 258007 633590 258069 0 FreeSans 400 0 0 0 gpio_loopback_zero[4]
port 813 nsew
flabel metal3 633270 303007 633590 303069 0 FreeSans 400 0 0 0 gpio_loopback_zero[5]
port 812 nsew
flabel metal3 633270 348007 633590 348069 0 FreeSans 400 0 0 0 gpio_loopback_zero[6]
port 811 nsew
flabel metal3 633270 525007 633590 525069 0 FreeSans 400 0 0 0 gpio_loopback_zero[7]
port 810 nsew
flabel metal3 633270 570007 633590 570069 0 FreeSans 400 0 0 0 gpio_loopback_zero[8]
port 809 nsew
flabel metal3 633270 615007 633590 615069 0 FreeSans 400 0 0 0 gpio_loopback_zero[9]
port 808 nsew
flabel metal3 633270 660007 633590 660069 0 FreeSans 400 0 0 0 gpio_loopback_zero[10]
port 807 nsew
flabel metal3 633270 705007 633590 705069 0 FreeSans 400 0 0 0 gpio_loopback_zero[11]
port 806 nsew
flabel metal3 633270 750007 633590 750069 0 FreeSans 400 0 0 0 gpio_loopback_zero[12]
port 805 nsew
flabel metal3 633270 839007 633590 839069 0 FreeSans 400 0 0 0 gpio_loopback_zero[13]
port 804 nsew
flabel metal3 633270 929007 633590 929069 0 FreeSans 400 0 0 0 gpio_loopback_zero[14]
port 803 nsew
flabel metal3 -264 734644 56 734704 0 FreeSans 400 0 0 0 gpio_loopback_zero[25]
port 792 nsew
flabel metal3 -264 648644 56 648704 0 FreeSans 400 0 0 0 gpio_loopback_zero[27]
port 790 nsew
flabel metal3 -264 562644 56 562704 0 FreeSans 400 0 0 0 gpio_loopback_zero[29]
port 788 nsew
flabel metal3 -264 476644 56 476704 0 FreeSans 400 0 0 0 gpio_loopback_zero[31]
port 786 nsew
flabel metal3 -264 304644 56 304704 0 FreeSans 400 0 0 0 gpio_loopback_zero[33]
port 784 nsew
flabel metal3 -264 218644 56 218704 0 FreeSans 400 0 0 0 gpio_loopback_zero[35]
port 782 nsew
flabel metal3 -264 132644 56 132704 0 FreeSans 400 0 0 0 gpio_loopback_zero[37]
port 780 nsew
flabel metal3 -264 904644 56 904704 0 FreeSans 400 0 0 0 gpio_loopback_zero[24]
port 793 nsew
flabel metal3 -264 691644 56 691704 0 FreeSans 400 0 0 0 gpio_loopback_zero[26]
port 791 nsew
flabel metal3 -264 605644 56 605704 0 FreeSans 400 0 0 0 gpio_loopback_zero[28]
port 789 nsew
flabel metal3 -264 519644 56 519704 0 FreeSans 400 0 0 0 gpio_loopback_zero[30]
port 787 nsew
flabel metal3 -264 347644 56 347704 0 FreeSans 400 0 0 0 gpio_loopback_zero[32]
port 785 nsew
flabel metal3 -264 261644 56 261704 0 FreeSans 400 0 0 0 gpio_loopback_zero[34]
port 783 nsew
flabel metal3 -264 175644 56 175704 0 FreeSans 400 0 0 0 gpio_loopback_zero[36]
port 781 nsew
flabel metal2 27497 953270 27558 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[23]
port 794 nsew
flabel metal2 78697 953270 78758 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[22]
port 795 nsew
flabel metal2 129897 953270 129958 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[21]
port 796 nsew
flabel metal2 181097 953270 181158 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[20]
port 797 nsew
flabel metal2 232297 953270 232358 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[19]
port 798 nsew
flabel metal2 336697 953270 336758 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[18]
port 799 nsew
flabel metal2 425697 953270 425758 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[17]
port 800 nsew
flabel metal2 476897 953270 476958 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[16]
port 801 nsew
flabel metal2 576297 953270 576358 953590 0 FreeSans 400 90 0 0 gpio_loopback_zero[15]
port 802 nsew
<< properties >>
string FIXED_BBOX 0 0 633326 953326
<< end >>
